`timescale 1ns / 1ps
module letras (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (k[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= k[vcount- posy][hcount- posx][7:5];
				green <= k[vcount- posy][hcount- posx][4:2];
            blue 	<= k[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 150;
parameter RESOLUCION_Y = 25;
wire [8:0] k[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign k[9][17] = 9'b111111111;
assign k[9][18] = 9'b111111111;
assign k[9][19] = 9'b111111111;
assign k[9][20] = 9'b111111111;
assign k[9][21] = 9'b111111111;
assign k[9][22] = 9'b111111111;
assign k[9][23] = 9'b111111111;
assign k[9][24] = 9'b111111111;
assign k[9][25] = 9'b111111111;
assign k[9][31] = 9'b110110110;
assign k[9][32] = 9'b111111111;
assign k[9][33] = 9'b111111111;
assign k[9][34] = 9'b111111111;
assign k[9][35] = 9'b111111111;
assign k[9][36] = 9'b111111111;
assign k[9][42] = 9'b110110110;
assign k[9][43] = 9'b111111111;
assign k[9][44] = 9'b111111111;
assign k[9][45] = 9'b111111111;
assign k[9][52] = 9'b111111111;
assign k[9][53] = 9'b111111111;
assign k[9][54] = 9'b111111111;
assign k[9][57] = 9'b111111111;
assign k[9][58] = 9'b111111111;
assign k[9][59] = 9'b111111111;
assign k[9][60] = 9'b111111111;
assign k[9][61] = 9'b111111111;
assign k[9][62] = 9'b111111111;
assign k[9][63] = 9'b111111111;
assign k[9][64] = 9'b111111111;
assign k[9][65] = 9'b111111111;
assign k[9][66] = 9'b111111111;
assign k[9][67] = 9'b111111111;
assign k[9][68] = 9'b111111111;
assign k[9][69] = 9'b111111111;
assign k[9][81] = 9'b111111111;
assign k[9][82] = 9'b111111111;
assign k[9][83] = 9'b111111111;
assign k[9][84] = 9'b111111111;
assign k[9][85] = 9'b111111111;
assign k[9][86] = 9'b111111111;
assign k[9][87] = 9'b111111111;
assign k[9][88] = 9'b111111111;
assign k[9][89] = 9'b111111111;
assign k[9][94] = 9'b111111111;
assign k[9][95] = 9'b111111111;
assign k[9][96] = 9'b111111111;
assign k[9][97] = 9'b110110110;
assign k[9][103] = 9'b111111111;
assign k[9][104] = 9'b111111111;
assign k[9][105] = 9'b111111111;
assign k[9][106] = 9'b111111111;
assign k[9][108] = 9'b111111111;
assign k[9][109] = 9'b111111111;
assign k[9][110] = 9'b111111111;
assign k[9][111] = 9'b111111111;
assign k[9][112] = 9'b111111111;
assign k[9][113] = 9'b111111111;
assign k[9][114] = 9'b111111111;
assign k[9][115] = 9'b111111111;
assign k[9][116] = 9'b111111111;
assign k[9][117] = 9'b111111111;
assign k[9][118] = 9'b111111111;
assign k[9][119] = 9'b111111111;
assign k[9][120] = 9'b111111111;
assign k[9][123] = 9'b111111111;
assign k[9][124] = 9'b111111111;
assign k[9][125] = 9'b111111111;
assign k[9][126] = 9'b111111111;
assign k[9][127] = 9'b111111111;
assign k[9][128] = 9'b111111111;
assign k[9][129] = 9'b111111111;
assign k[9][130] = 9'b111111111;
assign k[9][131] = 9'b111111111;
assign k[9][132] = 9'b111111111;
assign k[9][133] = 9'b111111111;
assign k[10][16] = 9'b111111111;
assign k[10][17] = 9'b111111111;
assign k[10][18] = 9'b111111111;
assign k[10][19] = 9'b111111111;
assign k[10][20] = 9'b111111111;
assign k[10][21] = 9'b111111111;
assign k[10][22] = 9'b111111111;
assign k[10][23] = 9'b111111111;
assign k[10][24] = 9'b111111111;
assign k[10][25] = 9'b111111111;
assign k[10][30] = 9'b111111111;
assign k[10][31] = 9'b111111111;
assign k[10][32] = 9'b111111111;
assign k[10][33] = 9'b111111111;
assign k[10][34] = 9'b111111111;
assign k[10][35] = 9'b111111111;
assign k[10][36] = 9'b111111111;
assign k[10][37] = 9'b111111111;
assign k[10][42] = 9'b111111111;
assign k[10][43] = 9'b111111111;
assign k[10][44] = 9'b111111111;
assign k[10][45] = 9'b111111111;
assign k[10][46] = 9'b111111111;
assign k[10][50] = 9'b111111111;
assign k[10][51] = 9'b111111111;
assign k[10][52] = 9'b111111111;
assign k[10][53] = 9'b111111111;
assign k[10][54] = 9'b111111111;
assign k[10][55] = 9'b110110110;
assign k[10][57] = 9'b111111111;
assign k[10][58] = 9'b111111111;
assign k[10][59] = 9'b111111111;
assign k[10][60] = 9'b111111111;
assign k[10][61] = 9'b111111111;
assign k[10][62] = 9'b111111111;
assign k[10][63] = 9'b111111111;
assign k[10][64] = 9'b111111111;
assign k[10][65] = 9'b111111111;
assign k[10][66] = 9'b111111111;
assign k[10][67] = 9'b111111111;
assign k[10][68] = 9'b111111111;
assign k[10][69] = 9'b111111111;
assign k[10][80] = 9'b111111111;
assign k[10][81] = 9'b111111111;
assign k[10][82] = 9'b111111111;
assign k[10][83] = 9'b111111111;
assign k[10][84] = 9'b111111111;
assign k[10][85] = 9'b111111111;
assign k[10][86] = 9'b111111111;
assign k[10][87] = 9'b111111111;
assign k[10][88] = 9'b111111111;
assign k[10][89] = 9'b111111111;
assign k[10][90] = 9'b111111111;
assign k[10][94] = 9'b111111111;
assign k[10][95] = 9'b111111111;
assign k[10][96] = 9'b111111111;
assign k[10][97] = 9'b111111111;
assign k[10][103] = 9'b111111111;
assign k[10][104] = 9'b111111111;
assign k[10][105] = 9'b111111111;
assign k[10][106] = 9'b111111111;
assign k[10][108] = 9'b111111111;
assign k[10][109] = 9'b111111111;
assign k[10][110] = 9'b111111111;
assign k[10][111] = 9'b111111111;
assign k[10][112] = 9'b111111111;
assign k[10][113] = 9'b111111111;
assign k[10][114] = 9'b111111111;
assign k[10][115] = 9'b111111111;
assign k[10][116] = 9'b111111111;
assign k[10][117] = 9'b111111111;
assign k[10][118] = 9'b111111111;
assign k[10][119] = 9'b111111111;
assign k[10][120] = 9'b111111111;
assign k[10][123] = 9'b111111111;
assign k[10][124] = 9'b111111111;
assign k[10][125] = 9'b111111111;
assign k[10][126] = 9'b111111111;
assign k[10][127] = 9'b111111111;
assign k[10][128] = 9'b111111111;
assign k[10][129] = 9'b111111111;
assign k[10][130] = 9'b111111111;
assign k[10][131] = 9'b111111111;
assign k[10][132] = 9'b111111111;
assign k[10][133] = 9'b111111111;
assign k[10][134] = 9'b111111111;
assign k[11][15] = 9'b111111111;
assign k[11][16] = 9'b111111111;
assign k[11][17] = 9'b111111111;
assign k[11][18] = 9'b111111111;
assign k[11][29] = 9'b110010010;
assign k[11][30] = 9'b111111111;
assign k[11][31] = 9'b111111111;
assign k[11][32] = 9'b111111111;
assign k[11][33] = 9'b110110110;
assign k[11][35] = 9'b111111111;
assign k[11][36] = 9'b111111111;
assign k[11][37] = 9'b111111111;
assign k[11][38] = 9'b111111111;
assign k[11][42] = 9'b111111111;
assign k[11][43] = 9'b111111111;
assign k[11][44] = 9'b111111111;
assign k[11][45] = 9'b111111111;
assign k[11][46] = 9'b111111111;
assign k[11][47] = 9'b111111111;
assign k[11][50] = 9'b111111111;
assign k[11][51] = 9'b111111111;
assign k[11][52] = 9'b111111111;
assign k[11][53] = 9'b111111111;
assign k[11][54] = 9'b111111111;
assign k[11][55] = 9'b110110110;
assign k[11][57] = 9'b111111111;
assign k[11][58] = 9'b111111111;
assign k[11][59] = 9'b111111111;
assign k[11][60] = 9'b111111111;
assign k[11][79] = 9'b111111111;
assign k[11][80] = 9'b111111111;
assign k[11][81] = 9'b111111111;
assign k[11][82] = 9'b111111111;
assign k[11][88] = 9'b111111111;
assign k[11][89] = 9'b111111111;
assign k[11][90] = 9'b111111111;
assign k[11][91] = 9'b111111111;
assign k[11][94] = 9'b111111111;
assign k[11][95] = 9'b111111111;
assign k[11][96] = 9'b111111111;
assign k[11][97] = 9'b111111111;
assign k[11][103] = 9'b111111111;
assign k[11][104] = 9'b111111111;
assign k[11][105] = 9'b111111111;
assign k[11][106] = 9'b111111111;
assign k[11][108] = 9'b111111111;
assign k[11][109] = 9'b111111111;
assign k[11][110] = 9'b111111111;
assign k[11][111] = 9'b111111111;
assign k[11][123] = 9'b111111111;
assign k[11][124] = 9'b111111111;
assign k[11][125] = 9'b111111111;
assign k[11][126] = 9'b111111111;
assign k[11][132] = 9'b111111111;
assign k[11][133] = 9'b111111111;
assign k[11][134] = 9'b111111111;
assign k[11][135] = 9'b111111111;
assign k[12][13] = 9'b111111111;
assign k[12][14] = 9'b111111111;
assign k[12][15] = 9'b111111111;
assign k[12][16] = 9'b111111111;
assign k[12][28] = 9'b111111111;
assign k[12][29] = 9'b111111111;
assign k[12][30] = 9'b111111111;
assign k[12][31] = 9'b111111111;
assign k[12][37] = 9'b111111111;
assign k[12][38] = 9'b111111111;
assign k[12][39] = 9'b111111111;
assign k[12][40] = 9'b111111111;
assign k[12][42] = 9'b111111111;
assign k[12][43] = 9'b111111111;
assign k[12][44] = 9'b111111111;
assign k[12][45] = 9'b111111111;
assign k[12][46] = 9'b111111111;
assign k[12][47] = 9'b111111111;
assign k[12][48] = 9'b111111111;
assign k[12][49] = 9'b111111111;
assign k[12][50] = 9'b111111111;
assign k[12][51] = 9'b111111111;
assign k[12][52] = 9'b111111111;
assign k[12][53] = 9'b111111111;
assign k[12][54] = 9'b111111111;
assign k[12][55] = 9'b110110110;
assign k[12][57] = 9'b111111111;
assign k[12][58] = 9'b111111111;
assign k[12][59] = 9'b111111111;
assign k[12][60] = 9'b111111111;
assign k[12][79] = 9'b111111111;
assign k[12][80] = 9'b111111111;
assign k[12][81] = 9'b111111111;
assign k[12][82] = 9'b111111111;
assign k[12][88] = 9'b111111111;
assign k[12][89] = 9'b111111111;
assign k[12][90] = 9'b111111111;
assign k[12][91] = 9'b111111111;
assign k[12][94] = 9'b111111111;
assign k[12][95] = 9'b111111111;
assign k[12][96] = 9'b111111111;
assign k[12][97] = 9'b110110110;
assign k[12][103] = 9'b111111111;
assign k[12][104] = 9'b111111111;
assign k[12][105] = 9'b111111111;
assign k[12][106] = 9'b111111111;
assign k[12][108] = 9'b111111111;
assign k[12][109] = 9'b111111111;
assign k[12][110] = 9'b111111111;
assign k[12][111] = 9'b111111111;
assign k[12][123] = 9'b111111111;
assign k[12][124] = 9'b111111111;
assign k[12][125] = 9'b111111111;
assign k[12][126] = 9'b111111111;
assign k[12][132] = 9'b111111111;
assign k[12][133] = 9'b111111111;
assign k[12][134] = 9'b111111111;
assign k[12][135] = 9'b111111111;
assign k[13][13] = 9'b111111111;
assign k[13][14] = 9'b111111111;
assign k[13][15] = 9'b111111111;
assign k[13][16] = 9'b111111111;
assign k[13][21] = 9'b111111111;
assign k[13][22] = 9'b111111111;
assign k[13][23] = 9'b111111111;
assign k[13][24] = 9'b111111111;
assign k[13][25] = 9'b111111111;
assign k[13][28] = 9'b111111111;
assign k[13][29] = 9'b111111111;
assign k[13][30] = 9'b111111111;
assign k[13][31] = 9'b111111111;
assign k[13][37] = 9'b111111111;
assign k[13][38] = 9'b111111111;
assign k[13][39] = 9'b111111111;
assign k[13][40] = 9'b111111111;
assign k[13][42] = 9'b111111111;
assign k[13][43] = 9'b111111111;
assign k[13][44] = 9'b111111111;
assign k[13][45] = 9'b111111111;
assign k[13][46] = 9'b111111111;
assign k[13][47] = 9'b111111111;
assign k[13][48] = 9'b111111111;
assign k[13][49] = 9'b111111111;
assign k[13][50] = 9'b111111111;
assign k[13][51] = 9'b111111111;
assign k[13][52] = 9'b111111111;
assign k[13][53] = 9'b111111111;
assign k[13][54] = 9'b111111111;
assign k[13][55] = 9'b110110110;
assign k[13][57] = 9'b111111111;
assign k[13][58] = 9'b111111111;
assign k[13][59] = 9'b111111111;
assign k[13][60] = 9'b111111111;
assign k[13][61] = 9'b111111111;
assign k[13][62] = 9'b111111111;
assign k[13][63] = 9'b111111111;
assign k[13][64] = 9'b111111111;
assign k[13][65] = 9'b111111111;
assign k[13][66] = 9'b111111111;
assign k[13][67] = 9'b111111111;
assign k[13][79] = 9'b111111111;
assign k[13][80] = 9'b111111111;
assign k[13][81] = 9'b111111111;
assign k[13][82] = 9'b111111111;
assign k[13][88] = 9'b111111111;
assign k[13][89] = 9'b111111111;
assign k[13][90] = 9'b111111111;
assign k[13][91] = 9'b111111111;
assign k[13][94] = 9'b111111111;
assign k[13][95] = 9'b111111111;
assign k[13][96] = 9'b111111111;
assign k[13][97] = 9'b111111111;
assign k[13][98] = 9'b111111111;
assign k[13][101] = 9'b111111111;
assign k[13][102] = 9'b111111111;
assign k[13][103] = 9'b111111111;
assign k[13][104] = 9'b111111111;
assign k[13][105] = 9'b111111111;
assign k[13][106] = 9'b111111111;
assign k[13][108] = 9'b111111111;
assign k[13][109] = 9'b111111111;
assign k[13][110] = 9'b111111111;
assign k[13][111] = 9'b111111111;
assign k[13][112] = 9'b111111111;
assign k[13][113] = 9'b111111111;
assign k[13][114] = 9'b111111111;
assign k[13][115] = 9'b111111111;
assign k[13][116] = 9'b111111111;
assign k[13][117] = 9'b111111111;
assign k[13][118] = 9'b111111111;
assign k[13][123] = 9'b111111111;
assign k[13][124] = 9'b111111111;
assign k[13][125] = 9'b111111111;
assign k[13][126] = 9'b111111111;
assign k[13][131] = 9'b111111111;
assign k[13][132] = 9'b111111111;
assign k[13][133] = 9'b111111111;
assign k[13][134] = 9'b111111111;
assign k[13][135] = 9'b111111111;
assign k[14][13] = 9'b111111111;
assign k[14][14] = 9'b111111111;
assign k[14][15] = 9'b111111111;
assign k[14][16] = 9'b111111111;
assign k[14][20] = 9'b111111111;
assign k[14][21] = 9'b111111111;
assign k[14][22] = 9'b111111111;
assign k[14][23] = 9'b111111111;
assign k[14][24] = 9'b111111111;
assign k[14][25] = 9'b111111111;
assign k[14][28] = 9'b111111111;
assign k[14][29] = 9'b111111111;
assign k[14][30] = 9'b111111111;
assign k[14][31] = 9'b111111111;
assign k[14][37] = 9'b111111111;
assign k[14][38] = 9'b111111111;
assign k[14][39] = 9'b111111111;
assign k[14][40] = 9'b111111111;
assign k[14][42] = 9'b111111111;
assign k[14][43] = 9'b111111111;
assign k[14][44] = 9'b111111111;
assign k[14][45] = 9'b111111111;
assign k[14][46] = 9'b111111111;
assign k[14][47] = 9'b111111111;
assign k[14][48] = 9'b111111111;
assign k[14][49] = 9'b111111111;
assign k[14][50] = 9'b111111111;
assign k[14][51] = 9'b111111111;
assign k[14][52] = 9'b111111111;
assign k[14][53] = 9'b111111111;
assign k[14][54] = 9'b111111111;
assign k[14][55] = 9'b110110110;
assign k[14][57] = 9'b111111111;
assign k[14][58] = 9'b111111111;
assign k[14][59] = 9'b111111111;
assign k[14][60] = 9'b111111111;
assign k[14][61] = 9'b111111111;
assign k[14][62] = 9'b111111111;
assign k[14][63] = 9'b111111111;
assign k[14][64] = 9'b111111111;
assign k[14][65] = 9'b111111111;
assign k[14][66] = 9'b111111111;
assign k[14][67] = 9'b111111111;
assign k[14][79] = 9'b111111111;
assign k[14][80] = 9'b111111111;
assign k[14][81] = 9'b111111111;
assign k[14][82] = 9'b111111111;
assign k[14][88] = 9'b111111111;
assign k[14][89] = 9'b111111111;
assign k[14][90] = 9'b111111111;
assign k[14][91] = 9'b111111111;
assign k[14][94] = 9'b111111111;
assign k[14][95] = 9'b111111111;
assign k[14][96] = 9'b111111111;
assign k[14][97] = 9'b111111111;
assign k[14][98] = 9'b111111111;
assign k[14][101] = 9'b111111111;
assign k[14][102] = 9'b111111111;
assign k[14][103] = 9'b111111111;
assign k[14][104] = 9'b111111111;
assign k[14][105] = 9'b111111111;
assign k[14][106] = 9'b111111111;
assign k[14][108] = 9'b111111111;
assign k[14][109] = 9'b111111111;
assign k[14][110] = 9'b111111111;
assign k[14][111] = 9'b111111111;
assign k[14][112] = 9'b111111111;
assign k[14][113] = 9'b111111111;
assign k[14][114] = 9'b111111111;
assign k[14][115] = 9'b111111111;
assign k[14][116] = 9'b111111111;
assign k[14][117] = 9'b111111111;
assign k[14][118] = 9'b111111111;
assign k[14][119] = 9'b110110110;
assign k[14][123] = 9'b111111111;
assign k[14][124] = 9'b111111111;
assign k[14][125] = 9'b111111111;
assign k[14][126] = 9'b111111111;
assign k[14][130] = 9'b111111111;
assign k[14][131] = 9'b111111111;
assign k[14][132] = 9'b111111111;
assign k[14][133] = 9'b111111111;
assign k[14][134] = 9'b111111111;
assign k[14][135] = 9'b111111111;
assign k[15][13] = 9'b111111111;
assign k[15][14] = 9'b111111111;
assign k[15][15] = 9'b111111111;
assign k[15][16] = 9'b111111111;
assign k[15][22] = 9'b111111111;
assign k[15][23] = 9'b111111111;
assign k[15][24] = 9'b111111111;
assign k[15][25] = 9'b111111111;
assign k[15][28] = 9'b111111111;
assign k[15][29] = 9'b111111111;
assign k[15][30] = 9'b111111111;
assign k[15][31] = 9'b111111111;
assign k[15][32] = 9'b111111111;
assign k[15][33] = 9'b111111111;
assign k[15][34] = 9'b111111111;
assign k[15][35] = 9'b111111111;
assign k[15][36] = 9'b111111111;
assign k[15][37] = 9'b111111111;
assign k[15][38] = 9'b111111111;
assign k[15][39] = 9'b111111111;
assign k[15][40] = 9'b111111111;
assign k[15][42] = 9'b111111111;
assign k[15][43] = 9'b111111111;
assign k[15][44] = 9'b111111111;
assign k[15][45] = 9'b111111111;
assign k[15][46] = 9'b111111111;
assign k[15][48] = 9'b111111111;
assign k[15][49] = 9'b111111111;
assign k[15][51] = 9'b111111111;
assign k[15][52] = 9'b111111111;
assign k[15][53] = 9'b111111111;
assign k[15][54] = 9'b111111111;
assign k[15][55] = 9'b110110110;
assign k[15][57] = 9'b111111111;
assign k[15][58] = 9'b111111111;
assign k[15][59] = 9'b111111111;
assign k[15][60] = 9'b111111111;
assign k[15][79] = 9'b111111111;
assign k[15][80] = 9'b111111111;
assign k[15][81] = 9'b111111111;
assign k[15][82] = 9'b111111111;
assign k[15][88] = 9'b111111111;
assign k[15][89] = 9'b111111111;
assign k[15][90] = 9'b111111111;
assign k[15][91] = 9'b111111111;
assign k[15][95] = 9'b111111111;
assign k[15][96] = 9'b111111111;
assign k[15][97] = 9'b111111111;
assign k[15][98] = 9'b111111111;
assign k[15][99] = 9'b111111111;
assign k[15][100] = 9'b111111111;
assign k[15][101] = 9'b111111111;
assign k[15][102] = 9'b111111111;
assign k[15][103] = 9'b111111111;
assign k[15][104] = 9'b111111111;
assign k[15][108] = 9'b111111111;
assign k[15][109] = 9'b111111111;
assign k[15][110] = 9'b111111111;
assign k[15][111] = 9'b111111111;
assign k[15][123] = 9'b111111111;
assign k[15][124] = 9'b111111111;
assign k[15][125] = 9'b111111111;
assign k[15][126] = 9'b111111111;
assign k[15][127] = 9'b111111111;
assign k[15][128] = 9'b111111111;
assign k[15][129] = 9'b111111111;
assign k[15][130] = 9'b111111111;
assign k[15][131] = 9'b111111111;
assign k[16][13] = 9'b111111111;
assign k[16][14] = 9'b111111111;
assign k[16][15] = 9'b111111111;
assign k[16][16] = 9'b111111111;
assign k[16][17] = 9'b111111111;
assign k[16][22] = 9'b111111111;
assign k[16][23] = 9'b111111111;
assign k[16][24] = 9'b111111111;
assign k[16][25] = 9'b111111111;
assign k[16][28] = 9'b111111111;
assign k[16][29] = 9'b111111111;
assign k[16][30] = 9'b111111111;
assign k[16][31] = 9'b111111111;
assign k[16][32] = 9'b111111111;
assign k[16][33] = 9'b111111111;
assign k[16][34] = 9'b111111111;
assign k[16][35] = 9'b111111111;
assign k[16][36] = 9'b111111111;
assign k[16][37] = 9'b111111111;
assign k[16][38] = 9'b111111111;
assign k[16][39] = 9'b111111111;
assign k[16][40] = 9'b111111111;
assign k[16][42] = 9'b111111111;
assign k[16][43] = 9'b111111111;
assign k[16][44] = 9'b111111111;
assign k[16][45] = 9'b111111111;
assign k[16][48] = 9'b111111111;
assign k[16][49] = 9'b111111111;
assign k[16][52] = 9'b111111111;
assign k[16][53] = 9'b111111111;
assign k[16][54] = 9'b111111111;
assign k[16][55] = 9'b110110110;
assign k[16][57] = 9'b111111111;
assign k[16][58] = 9'b111111111;
assign k[16][59] = 9'b111111111;
assign k[16][60] = 9'b111111111;
assign k[16][79] = 9'b111111111;
assign k[16][80] = 9'b111111111;
assign k[16][81] = 9'b111111111;
assign k[16][82] = 9'b111111111;
assign k[16][88] = 9'b111111111;
assign k[16][89] = 9'b111111111;
assign k[16][90] = 9'b111111111;
assign k[16][91] = 9'b111111111;
assign k[16][96] = 9'b111111111;
assign k[16][97] = 9'b111111111;
assign k[16][98] = 9'b111111111;
assign k[16][99] = 9'b111111111;
assign k[16][100] = 9'b111111111;
assign k[16][101] = 9'b111111111;
assign k[16][102] = 9'b111111111;
assign k[16][103] = 9'b111111111;
assign k[16][104] = 9'b111111111;
assign k[16][108] = 9'b111111111;
assign k[16][109] = 9'b111111111;
assign k[16][110] = 9'b111111111;
assign k[16][111] = 9'b111111111;
assign k[16][123] = 9'b111111111;
assign k[16][124] = 9'b111111111;
assign k[16][125] = 9'b111111111;
assign k[16][126] = 9'b111111111;
assign k[16][127] = 9'b111111111;
assign k[16][128] = 9'b111111111;
assign k[16][129] = 9'b111111111;
assign k[16][130] = 9'b111111111;
assign k[16][131] = 9'b111111111;
assign k[16][132] = 9'b111111111;
assign k[16][133] = 9'b111111111;
assign k[17][15] = 9'b111111111;
assign k[17][16] = 9'b111111111;
assign k[17][17] = 9'b111111111;
assign k[17][18] = 9'b111111111;
assign k[17][22] = 9'b111111111;
assign k[17][23] = 9'b111111111;
assign k[17][24] = 9'b111111111;
assign k[17][25] = 9'b111111111;
assign k[17][28] = 9'b111111111;
assign k[17][29] = 9'b111111111;
assign k[17][30] = 9'b111111111;
assign k[17][31] = 9'b111111111;
assign k[17][37] = 9'b111111111;
assign k[17][38] = 9'b111111111;
assign k[17][39] = 9'b111111111;
assign k[17][40] = 9'b111111111;
assign k[17][42] = 9'b111111111;
assign k[17][43] = 9'b111111111;
assign k[17][44] = 9'b111111111;
assign k[17][45] = 9'b111111111;
assign k[17][51] = 9'b111111111;
assign k[17][52] = 9'b111111111;
assign k[17][53] = 9'b111111111;
assign k[17][54] = 9'b111111111;
assign k[17][55] = 9'b110110110;
assign k[17][57] = 9'b111111111;
assign k[17][58] = 9'b111111111;
assign k[17][59] = 9'b111111111;
assign k[17][60] = 9'b111111111;
assign k[17][79] = 9'b111111111;
assign k[17][80] = 9'b111111111;
assign k[17][81] = 9'b111111111;
assign k[17][82] = 9'b111111111;
assign k[17][88] = 9'b111111111;
assign k[17][89] = 9'b111111111;
assign k[17][90] = 9'b111111111;
assign k[17][91] = 9'b111111111;
assign k[17][97] = 9'b111111111;
assign k[17][98] = 9'b111111111;
assign k[17][99] = 9'b111111111;
assign k[17][100] = 9'b111111111;
assign k[17][101] = 9'b111111111;
assign k[17][102] = 9'b111111111;
assign k[17][108] = 9'b111111111;
assign k[17][109] = 9'b111111111;
assign k[17][110] = 9'b111111111;
assign k[17][111] = 9'b111111111;
assign k[17][123] = 9'b111111111;
assign k[17][124] = 9'b111111111;
assign k[17][125] = 9'b111111111;
assign k[17][126] = 9'b111111111;
assign k[17][128] = 9'b111111111;
assign k[17][129] = 9'b111111111;
assign k[17][130] = 9'b111111111;
assign k[17][131] = 9'b111111111;
assign k[17][132] = 9'b111111111;
assign k[17][133] = 9'b111111111;
assign k[18][17] = 9'b111111111;
assign k[18][18] = 9'b111111111;
assign k[18][19] = 9'b111111111;
assign k[18][20] = 9'b111111111;
assign k[18][21] = 9'b111111111;
assign k[18][22] = 9'b111111111;
assign k[18][23] = 9'b111111111;
assign k[18][24] = 9'b111111111;
assign k[18][25] = 9'b111111111;
assign k[18][28] = 9'b111111111;
assign k[18][29] = 9'b111111111;
assign k[18][30] = 9'b111111111;
assign k[18][31] = 9'b111111111;
assign k[18][37] = 9'b111111111;
assign k[18][38] = 9'b111111111;
assign k[18][39] = 9'b111111111;
assign k[18][40] = 9'b111111111;
assign k[18][42] = 9'b111111111;
assign k[18][43] = 9'b111111111;
assign k[18][44] = 9'b111111111;
assign k[18][45] = 9'b111111111;
assign k[18][51] = 9'b111111111;
assign k[18][52] = 9'b111111111;
assign k[18][53] = 9'b111111111;
assign k[18][54] = 9'b111111111;
assign k[18][55] = 9'b110110110;
assign k[18][57] = 9'b111111111;
assign k[18][58] = 9'b111111111;
assign k[18][59] = 9'b111111111;
assign k[18][60] = 9'b111111111;
assign k[18][61] = 9'b111111111;
assign k[18][62] = 9'b111111111;
assign k[18][63] = 9'b111111111;
assign k[18][64] = 9'b111111111;
assign k[18][65] = 9'b111111111;
assign k[18][66] = 9'b111111111;
assign k[18][67] = 9'b111111111;
assign k[18][68] = 9'b111111111;
assign k[18][69] = 9'b111111111;
assign k[18][81] = 9'b111111111;
assign k[18][82] = 9'b111111111;
assign k[18][83] = 9'b111111111;
assign k[18][84] = 9'b111111111;
assign k[18][85] = 9'b111111111;
assign k[18][86] = 9'b111111111;
assign k[18][87] = 9'b111111111;
assign k[18][88] = 9'b111111111;
assign k[18][89] = 9'b111111111;
assign k[18][99] = 9'b111111111;
assign k[18][100] = 9'b111111111;
assign k[18][108] = 9'b111111111;
assign k[18][109] = 9'b111111111;
assign k[18][110] = 9'b111111111;
assign k[18][111] = 9'b111111111;
assign k[18][112] = 9'b111111111;
assign k[18][113] = 9'b111111111;
assign k[18][114] = 9'b111111111;
assign k[18][115] = 9'b111111111;
assign k[18][116] = 9'b111111111;
assign k[18][117] = 9'b111111111;
assign k[18][118] = 9'b111111111;
assign k[18][119] = 9'b111111111;
assign k[18][120] = 9'b111111111;
assign k[18][123] = 9'b111111111;
assign k[18][124] = 9'b111111111;
assign k[18][125] = 9'b111111111;
assign k[18][126] = 9'b111111111;
assign k[18][130] = 9'b111111111;
assign k[18][131] = 9'b111111111;
assign k[18][132] = 9'b111111111;
assign k[18][133] = 9'b111111111;
assign k[18][134] = 9'b111111111;
assign k[18][135] = 9'b111111111;
assign k[19][17] = 9'b111111111;
assign k[19][18] = 9'b111111111;
assign k[19][19] = 9'b111111111;
assign k[19][20] = 9'b111111111;
assign k[19][21] = 9'b111111111;
assign k[19][22] = 9'b111111111;
assign k[19][23] = 9'b111111111;
assign k[19][24] = 9'b111111111;
assign k[19][25] = 9'b111111111;
assign k[19][28] = 9'b111111111;
assign k[19][29] = 9'b111111111;
assign k[19][30] = 9'b111111111;
assign k[19][31] = 9'b111111111;
assign k[19][37] = 9'b111111111;
assign k[19][38] = 9'b111111111;
assign k[19][39] = 9'b111111111;
assign k[19][40] = 9'b111111111;
assign k[19][43] = 9'b111111111;
assign k[19][44] = 9'b111111111;
assign k[19][45] = 9'b111111111;
assign k[19][52] = 9'b111111111;
assign k[19][53] = 9'b111111111;
assign k[19][54] = 9'b111111111;
assign k[19][57] = 9'b111111111;
assign k[19][58] = 9'b111111111;
assign k[19][59] = 9'b111111111;
assign k[19][60] = 9'b111111111;
assign k[19][61] = 9'b111111111;
assign k[19][62] = 9'b111111111;
assign k[19][63] = 9'b111111111;
assign k[19][64] = 9'b111111111;
assign k[19][65] = 9'b111111111;
assign k[19][66] = 9'b111111111;
assign k[19][67] = 9'b111111111;
assign k[19][68] = 9'b111111111;
assign k[19][69] = 9'b111111111;
assign k[19][81] = 9'b111111111;
assign k[19][82] = 9'b111111111;
assign k[19][83] = 9'b111111111;
assign k[19][84] = 9'b111111111;
assign k[19][85] = 9'b111111111;
assign k[19][86] = 9'b111111111;
assign k[19][87] = 9'b111111111;
assign k[19][88] = 9'b111111111;
assign k[19][89] = 9'b111111111;
assign k[19][99] = 9'b111111111;
assign k[19][100] = 9'b111111111;
assign k[19][108] = 9'b110110110;
assign k[19][109] = 9'b111111111;
assign k[19][110] = 9'b111111111;
assign k[19][111] = 9'b111111111;
assign k[19][112] = 9'b111111111;
assign k[19][113] = 9'b111111111;
assign k[19][114] = 9'b111111111;
assign k[19][115] = 9'b111111111;
assign k[19][116] = 9'b111111111;
assign k[19][117] = 9'b111111111;
assign k[19][118] = 9'b111111111;
assign k[19][119] = 9'b111111111;
assign k[19][120] = 9'b111111111;
assign k[19][123] = 9'b111111111;
assign k[19][124] = 9'b111111111;
assign k[19][125] = 9'b111111111;
assign k[19][126] = 9'b111111111;
assign k[19][130] = 9'b110110110;
assign k[19][131] = 9'b111111111;
assign k[19][132] = 9'b111111111;
assign k[19][133] = 9'b111111111;
assign k[19][134] = 9'b111111111;
assign k[19][135] = 9'b111111111;
//Total de Lineas = 778
endmodule

