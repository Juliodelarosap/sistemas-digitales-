/*`timescale 1ns / 1ps
module prueba_5 (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (micromatrizz[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= micromatrizz[vcount- posy][hcount- posx][7:5];
				green <= micromatrizz[vcount- posy][hcount- posx][4:2];
            blue 	<= micromatrizz[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 640;
parameter RESOLUCION_Y = 100;
wire [8:0] micromatrizz[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign micromatrizz[0][0] = 9'b111111111;
assign micromatrizz[0][1] = 9'b111111111;
assign micromatrizz[0][2] = 9'b111111111;
assign micromatrizz[0][3] = 9'b111111111;
assign micromatrizz[0][4] = 9'b111111111;
assign micromatrizz[0][5] = 9'b111111111;
assign micromatrizz[0][6] = 9'b111111111;
assign micromatrizz[0][7] = 9'b111111111;
assign micromatrizz[0][8] = 9'b111111111;
assign micromatrizz[0][9] = 9'b111111111;
assign micromatrizz[0][10] = 9'b111111111;
assign micromatrizz[0][11] = 9'b111111111;
assign micromatrizz[0][12] = 9'b111111111;
assign micromatrizz[0][13] = 9'b111111111;
assign micromatrizz[0][14] = 9'b111111111;
assign micromatrizz[0][15] = 9'b111111111;
assign micromatrizz[0][16] = 9'b111111111;
assign micromatrizz[0][17] = 9'b111111111;
assign micromatrizz[0][18] = 9'b111111111;
assign micromatrizz[0][19] = 9'b111111111;
assign micromatrizz[0][20] = 9'b111111111;
assign micromatrizz[0][21] = 9'b111111111;
assign micromatrizz[0][22] = 9'b111111111;
assign micromatrizz[0][23] = 9'b111111111;
assign micromatrizz[0][24] = 9'b111111111;
assign micromatrizz[0][25] = 9'b111111111;
assign micromatrizz[0][26] = 9'b111111111;
assign micromatrizz[0][27] = 9'b111111111;
assign micromatrizz[0][28] = 9'b111111111;
assign micromatrizz[0][29] = 9'b111111111;
assign micromatrizz[0][30] = 9'b111111111;
assign micromatrizz[0][31] = 9'b111111111;
assign micromatrizz[0][32] = 9'b111111111;
assign micromatrizz[0][33] = 9'b111111111;
assign micromatrizz[0][34] = 9'b111111111;
assign micromatrizz[0][35] = 9'b111111111;
assign micromatrizz[0][36] = 9'b111111111;
assign micromatrizz[0][37] = 9'b111111111;
assign micromatrizz[0][38] = 9'b111111111;
assign micromatrizz[0][39] = 9'b111111111;
assign micromatrizz[0][40] = 9'b111111111;
assign micromatrizz[0][41] = 9'b111111111;
assign micromatrizz[0][42] = 9'b111111111;
assign micromatrizz[0][43] = 9'b111111111;
assign micromatrizz[0][44] = 9'b111111111;
assign micromatrizz[0][45] = 9'b111111111;
assign micromatrizz[0][46] = 9'b111111111;
assign micromatrizz[0][47] = 9'b111111111;
assign micromatrizz[0][48] = 9'b111111111;
assign micromatrizz[0][49] = 9'b111111111;
assign micromatrizz[0][50] = 9'b111111111;
assign micromatrizz[0][51] = 9'b111111111;
assign micromatrizz[0][52] = 9'b111111111;
assign micromatrizz[0][53] = 9'b111111111;
assign micromatrizz[0][54] = 9'b111111111;
assign micromatrizz[0][55] = 9'b111111111;
assign micromatrizz[0][56] = 9'b111111111;
assign micromatrizz[0][57] = 9'b111111111;
assign micromatrizz[0][58] = 9'b111111111;
assign micromatrizz[0][59] = 9'b111111111;
assign micromatrizz[0][60] = 9'b111111111;
assign micromatrizz[0][61] = 9'b111111111;
assign micromatrizz[0][62] = 9'b111111111;
assign micromatrizz[0][63] = 9'b111111111;
assign micromatrizz[0][64] = 9'b111111111;
assign micromatrizz[0][65] = 9'b111111111;
assign micromatrizz[0][66] = 9'b111111111;
assign micromatrizz[0][67] = 9'b111111111;
assign micromatrizz[0][68] = 9'b111111111;
assign micromatrizz[0][69] = 9'b111111111;
assign micromatrizz[0][70] = 9'b111111111;
assign micromatrizz[0][71] = 9'b111111111;
assign micromatrizz[0][72] = 9'b111111111;
assign micromatrizz[0][73] = 9'b111111111;
assign micromatrizz[0][74] = 9'b111111111;
assign micromatrizz[0][75] = 9'b111111111;
assign micromatrizz[0][76] = 9'b111111111;
assign micromatrizz[0][77] = 9'b111111111;
assign micromatrizz[0][78] = 9'b111111111;
assign micromatrizz[0][79] = 9'b111111111;
assign micromatrizz[0][80] = 9'b111111111;
assign micromatrizz[0][81] = 9'b111111111;
assign micromatrizz[0][82] = 9'b111111111;
assign micromatrizz[0][83] = 9'b111111111;
assign micromatrizz[0][84] = 9'b111111111;
assign micromatrizz[0][85] = 9'b111111111;
assign micromatrizz[0][86] = 9'b111111111;
assign micromatrizz[0][87] = 9'b111111111;
assign micromatrizz[0][88] = 9'b111111111;
assign micromatrizz[0][89] = 9'b111111111;
assign micromatrizz[0][90] = 9'b111111111;
assign micromatrizz[0][91] = 9'b111111111;
assign micromatrizz[0][92] = 9'b111111111;
assign micromatrizz[0][93] = 9'b111111111;
assign micromatrizz[0][94] = 9'b111111111;
assign micromatrizz[0][95] = 9'b111111111;
assign micromatrizz[0][96] = 9'b111111111;
assign micromatrizz[0][97] = 9'b111111111;
assign micromatrizz[0][98] = 9'b111111111;
assign micromatrizz[0][99] = 9'b111111111;
assign micromatrizz[0][100] = 9'b111111111;
assign micromatrizz[0][101] = 9'b111111111;
assign micromatrizz[0][102] = 9'b111111111;
assign micromatrizz[0][103] = 9'b111111111;
assign micromatrizz[0][104] = 9'b111111111;
assign micromatrizz[0][105] = 9'b111111111;
assign micromatrizz[0][106] = 9'b111111111;
assign micromatrizz[0][107] = 9'b111111111;
assign micromatrizz[0][108] = 9'b111111111;
assign micromatrizz[0][109] = 9'b111111111;
assign micromatrizz[0][110] = 9'b111111111;
assign micromatrizz[0][111] = 9'b111111111;
assign micromatrizz[0][112] = 9'b111111111;
assign micromatrizz[0][113] = 9'b111111111;
assign micromatrizz[0][114] = 9'b111111111;
assign micromatrizz[0][115] = 9'b111111111;
assign micromatrizz[0][116] = 9'b111111111;
assign micromatrizz[0][117] = 9'b111111111;
assign micromatrizz[0][118] = 9'b111111111;
assign micromatrizz[0][119] = 9'b111111111;
assign micromatrizz[0][120] = 9'b111111111;
assign micromatrizz[0][121] = 9'b111111111;
assign micromatrizz[0][122] = 9'b111111111;
assign micromatrizz[0][123] = 9'b111111111;
assign micromatrizz[0][124] = 9'b111111111;
assign micromatrizz[0][125] = 9'b111111111;
assign micromatrizz[0][126] = 9'b111111111;
assign micromatrizz[0][127] = 9'b111111111;
assign micromatrizz[0][128] = 9'b111111111;
assign micromatrizz[0][129] = 9'b111111111;
assign micromatrizz[0][130] = 9'b111111111;
assign micromatrizz[0][131] = 9'b111111111;
assign micromatrizz[0][132] = 9'b111111111;
assign micromatrizz[0][133] = 9'b111111111;
assign micromatrizz[0][134] = 9'b111111111;
assign micromatrizz[0][135] = 9'b111111111;
assign micromatrizz[0][136] = 9'b111111111;
assign micromatrizz[0][137] = 9'b111111111;
assign micromatrizz[0][138] = 9'b111111111;
assign micromatrizz[0][139] = 9'b111111111;
assign micromatrizz[0][140] = 9'b111111111;
assign micromatrizz[0][141] = 9'b111111111;
assign micromatrizz[0][142] = 9'b111111111;
assign micromatrizz[0][143] = 9'b111111111;
assign micromatrizz[0][144] = 9'b111111111;
assign micromatrizz[0][145] = 9'b111111111;
assign micromatrizz[0][146] = 9'b111111111;
assign micromatrizz[0][147] = 9'b111111111;
assign micromatrizz[0][148] = 9'b111111111;
assign micromatrizz[0][149] = 9'b111111111;
assign micromatrizz[0][150] = 9'b111111111;
assign micromatrizz[0][151] = 9'b111111111;
assign micromatrizz[0][152] = 9'b111111111;
assign micromatrizz[0][153] = 9'b111111111;
assign micromatrizz[0][154] = 9'b111111111;
assign micromatrizz[0][155] = 9'b111111111;
assign micromatrizz[0][156] = 9'b111111111;
assign micromatrizz[0][157] = 9'b111111111;
assign micromatrizz[0][158] = 9'b111111111;
assign micromatrizz[0][159] = 9'b111111111;
assign micromatrizz[0][160] = 9'b111111111;
assign micromatrizz[0][161] = 9'b111111111;
assign micromatrizz[0][162] = 9'b111111111;
assign micromatrizz[0][163] = 9'b111111111;
assign micromatrizz[0][164] = 9'b111111111;
assign micromatrizz[0][165] = 9'b111111111;
assign micromatrizz[0][166] = 9'b111111111;
assign micromatrizz[0][167] = 9'b111111111;
assign micromatrizz[0][168] = 9'b111111111;
assign micromatrizz[0][169] = 9'b111111111;
assign micromatrizz[0][170] = 9'b111111111;
assign micromatrizz[0][171] = 9'b111111111;
assign micromatrizz[0][172] = 9'b111111111;
assign micromatrizz[0][173] = 9'b111111111;
assign micromatrizz[0][174] = 9'b111111111;
assign micromatrizz[0][175] = 9'b111111111;
assign micromatrizz[0][176] = 9'b111111111;
assign micromatrizz[0][177] = 9'b111111111;
assign micromatrizz[0][178] = 9'b111111111;
assign micromatrizz[0][179] = 9'b111111111;
assign micromatrizz[0][180] = 9'b111111111;
assign micromatrizz[0][181] = 9'b111111111;
assign micromatrizz[0][182] = 9'b111111111;
assign micromatrizz[0][183] = 9'b111111111;
assign micromatrizz[0][184] = 9'b111111111;
assign micromatrizz[0][185] = 9'b111111111;
assign micromatrizz[0][186] = 9'b111111111;
assign micromatrizz[0][187] = 9'b111111111;
assign micromatrizz[0][188] = 9'b111111111;
assign micromatrizz[0][189] = 9'b111111111;
assign micromatrizz[0][190] = 9'b111111111;
assign micromatrizz[0][191] = 9'b111111111;
assign micromatrizz[0][192] = 9'b111111111;
assign micromatrizz[0][193] = 9'b111111111;
assign micromatrizz[0][194] = 9'b111111111;
assign micromatrizz[0][195] = 9'b111111111;
assign micromatrizz[0][196] = 9'b111111111;
assign micromatrizz[0][197] = 9'b111111111;
assign micromatrizz[0][198] = 9'b111111111;
assign micromatrizz[0][199] = 9'b111111111;
assign micromatrizz[0][200] = 9'b111111111;
assign micromatrizz[0][201] = 9'b111111111;
assign micromatrizz[0][202] = 9'b111111111;
assign micromatrizz[0][203] = 9'b111111111;
assign micromatrizz[0][204] = 9'b111111111;
assign micromatrizz[0][205] = 9'b111111111;
assign micromatrizz[0][206] = 9'b111111111;
assign micromatrizz[0][207] = 9'b111111111;
assign micromatrizz[0][208] = 9'b111111111;
assign micromatrizz[0][209] = 9'b111111111;
assign micromatrizz[0][210] = 9'b111111111;
assign micromatrizz[0][211] = 9'b111111111;
assign micromatrizz[0][212] = 9'b111111111;
assign micromatrizz[0][213] = 9'b111111111;
assign micromatrizz[0][214] = 9'b111111111;
assign micromatrizz[0][215] = 9'b111111111;
assign micromatrizz[0][216] = 9'b111111111;
assign micromatrizz[0][217] = 9'b111111111;
assign micromatrizz[0][218] = 9'b111111111;
assign micromatrizz[0][219] = 9'b111111111;
assign micromatrizz[0][220] = 9'b111111111;
assign micromatrizz[0][221] = 9'b111111111;
assign micromatrizz[0][222] = 9'b111111111;
assign micromatrizz[0][223] = 9'b111111111;
assign micromatrizz[0][224] = 9'b111111111;
assign micromatrizz[0][225] = 9'b111111111;
assign micromatrizz[0][226] = 9'b111111111;
assign micromatrizz[0][227] = 9'b111111111;
assign micromatrizz[0][228] = 9'b111111111;
assign micromatrizz[0][229] = 9'b111111111;
assign micromatrizz[0][230] = 9'b111111111;
assign micromatrizz[0][231] = 9'b111111111;
assign micromatrizz[0][232] = 9'b111111111;
assign micromatrizz[0][233] = 9'b111111111;
assign micromatrizz[0][234] = 9'b111111111;
assign micromatrizz[0][235] = 9'b111111111;
assign micromatrizz[0][236] = 9'b111111111;
assign micromatrizz[0][237] = 9'b111111111;
assign micromatrizz[0][238] = 9'b111111111;
assign micromatrizz[0][239] = 9'b111111111;
assign micromatrizz[0][240] = 9'b111111111;
assign micromatrizz[0][241] = 9'b111111111;
assign micromatrizz[0][242] = 9'b111111111;
assign micromatrizz[0][243] = 9'b111111111;
assign micromatrizz[0][244] = 9'b111111111;
assign micromatrizz[0][245] = 9'b111111111;
assign micromatrizz[0][246] = 9'b111111111;
assign micromatrizz[0][247] = 9'b111111111;
assign micromatrizz[0][248] = 9'b111111111;
assign micromatrizz[0][249] = 9'b111111111;
assign micromatrizz[0][250] = 9'b111111111;
assign micromatrizz[0][251] = 9'b111111111;
assign micromatrizz[0][252] = 9'b111111111;
assign micromatrizz[0][253] = 9'b111111111;
assign micromatrizz[0][254] = 9'b111111111;
assign micromatrizz[0][255] = 9'b111111111;
assign micromatrizz[0][256] = 9'b111111111;
assign micromatrizz[0][257] = 9'b111111111;
assign micromatrizz[0][258] = 9'b111111111;
assign micromatrizz[0][259] = 9'b111111111;
assign micromatrizz[0][260] = 9'b111111111;
assign micromatrizz[0][261] = 9'b111111111;
assign micromatrizz[0][262] = 9'b111111111;
assign micromatrizz[0][263] = 9'b111111111;
assign micromatrizz[0][264] = 9'b111111111;
assign micromatrizz[0][265] = 9'b111111111;
assign micromatrizz[0][266] = 9'b111111111;
assign micromatrizz[0][267] = 9'b111111111;
assign micromatrizz[0][268] = 9'b111111111;
assign micromatrizz[0][269] = 9'b111111111;
assign micromatrizz[0][270] = 9'b111111111;
assign micromatrizz[0][271] = 9'b111111111;
assign micromatrizz[0][272] = 9'b111111111;
assign micromatrizz[0][273] = 9'b111111111;
assign micromatrizz[0][274] = 9'b111111111;
assign micromatrizz[0][275] = 9'b111111111;
assign micromatrizz[0][276] = 9'b111111111;
assign micromatrizz[0][277] = 9'b111111111;
assign micromatrizz[0][278] = 9'b111111111;
assign micromatrizz[0][279] = 9'b111111111;
assign micromatrizz[0][280] = 9'b111111111;
assign micromatrizz[0][281] = 9'b111111111;
assign micromatrizz[0][282] = 9'b111111111;
assign micromatrizz[0][283] = 9'b111111111;
assign micromatrizz[0][284] = 9'b111111111;
assign micromatrizz[0][285] = 9'b111111111;
assign micromatrizz[0][286] = 9'b111111111;
assign micromatrizz[0][287] = 9'b111111111;
assign micromatrizz[0][288] = 9'b111111111;
assign micromatrizz[0][289] = 9'b111111111;
assign micromatrizz[0][290] = 9'b111111111;
assign micromatrizz[0][291] = 9'b111111111;
assign micromatrizz[0][292] = 9'b111111111;
assign micromatrizz[0][293] = 9'b111111111;
assign micromatrizz[0][294] = 9'b111111111;
assign micromatrizz[0][295] = 9'b111111111;
assign micromatrizz[0][296] = 9'b111111111;
assign micromatrizz[0][297] = 9'b111111111;
assign micromatrizz[0][298] = 9'b111111111;
assign micromatrizz[0][299] = 9'b111111111;
assign micromatrizz[0][300] = 9'b111111111;
assign micromatrizz[0][301] = 9'b111111111;
assign micromatrizz[0][302] = 9'b111111111;
assign micromatrizz[0][303] = 9'b111111111;
assign micromatrizz[0][304] = 9'b111111111;
assign micromatrizz[0][305] = 9'b111111111;
assign micromatrizz[0][306] = 9'b111111111;
assign micromatrizz[0][307] = 9'b111111111;
assign micromatrizz[0][308] = 9'b111111111;
assign micromatrizz[0][309] = 9'b111111111;
assign micromatrizz[0][310] = 9'b111111111;
assign micromatrizz[0][311] = 9'b111111111;
assign micromatrizz[0][312] = 9'b111111111;
assign micromatrizz[0][313] = 9'b111111111;
assign micromatrizz[0][314] = 9'b111111111;
assign micromatrizz[0][315] = 9'b111111111;
assign micromatrizz[0][316] = 9'b111111111;
assign micromatrizz[0][317] = 9'b111111111;
assign micromatrizz[0][318] = 9'b111111111;
assign micromatrizz[0][319] = 9'b111111111;
assign micromatrizz[0][320] = 9'b111111111;
assign micromatrizz[0][321] = 9'b111111111;
assign micromatrizz[0][322] = 9'b111111111;
assign micromatrizz[0][323] = 9'b111111111;
assign micromatrizz[0][324] = 9'b111111111;
assign micromatrizz[0][325] = 9'b111111111;
assign micromatrizz[0][326] = 9'b111111111;
assign micromatrizz[0][327] = 9'b111111111;
assign micromatrizz[0][328] = 9'b111111111;
assign micromatrizz[0][329] = 9'b111111111;
assign micromatrizz[0][330] = 9'b111111111;
assign micromatrizz[0][331] = 9'b111111111;
assign micromatrizz[0][332] = 9'b111111111;
assign micromatrizz[0][333] = 9'b111111111;
assign micromatrizz[0][334] = 9'b111111111;
assign micromatrizz[0][335] = 9'b111111111;
assign micromatrizz[0][336] = 9'b111111111;
assign micromatrizz[0][337] = 9'b111111111;
assign micromatrizz[0][338] = 9'b111111111;
assign micromatrizz[0][339] = 9'b111111111;
assign micromatrizz[0][340] = 9'b111111111;
assign micromatrizz[0][341] = 9'b111111111;
assign micromatrizz[0][342] = 9'b111111111;
assign micromatrizz[0][343] = 9'b111111111;
assign micromatrizz[0][344] = 9'b111111111;
assign micromatrizz[0][345] = 9'b111111111;
assign micromatrizz[0][346] = 9'b111111111;
assign micromatrizz[0][347] = 9'b111111111;
assign micromatrizz[0][348] = 9'b111111111;
assign micromatrizz[0][349] = 9'b111111111;
assign micromatrizz[0][350] = 9'b111111111;
assign micromatrizz[0][351] = 9'b111111111;
assign micromatrizz[0][352] = 9'b111111111;
assign micromatrizz[0][353] = 9'b111111111;
assign micromatrizz[0][354] = 9'b111111111;
assign micromatrizz[0][355] = 9'b111111111;
assign micromatrizz[0][356] = 9'b111111111;
assign micromatrizz[0][357] = 9'b111111111;
assign micromatrizz[0][358] = 9'b111111111;
assign micromatrizz[0][359] = 9'b111111111;
assign micromatrizz[0][360] = 9'b111111111;
assign micromatrizz[0][361] = 9'b111111111;
assign micromatrizz[0][362] = 9'b111111111;
assign micromatrizz[0][363] = 9'b111111111;
assign micromatrizz[0][364] = 9'b111111111;
assign micromatrizz[0][365] = 9'b111111111;
assign micromatrizz[0][366] = 9'b111111111;
assign micromatrizz[0][367] = 9'b111111111;
assign micromatrizz[0][368] = 9'b111111111;
assign micromatrizz[0][369] = 9'b111111111;
assign micromatrizz[0][370] = 9'b111111111;
assign micromatrizz[0][371] = 9'b111111111;
assign micromatrizz[0][372] = 9'b111111111;
assign micromatrizz[0][373] = 9'b111111111;
assign micromatrizz[0][374] = 9'b111111111;
assign micromatrizz[0][375] = 9'b111111111;
assign micromatrizz[0][376] = 9'b111111111;
assign micromatrizz[0][377] = 9'b111111111;
assign micromatrizz[0][378] = 9'b111111111;
assign micromatrizz[0][379] = 9'b111111111;
assign micromatrizz[0][380] = 9'b111111111;
assign micromatrizz[0][381] = 9'b111111111;
assign micromatrizz[0][382] = 9'b111111111;
assign micromatrizz[0][383] = 9'b111111111;
assign micromatrizz[0][384] = 9'b111111111;
assign micromatrizz[0][385] = 9'b111111111;
assign micromatrizz[0][386] = 9'b111111111;
assign micromatrizz[0][387] = 9'b111111111;
assign micromatrizz[0][388] = 9'b111111111;
assign micromatrizz[0][389] = 9'b111111111;
assign micromatrizz[0][390] = 9'b111111111;
assign micromatrizz[0][391] = 9'b111111111;
assign micromatrizz[0][392] = 9'b111111111;
assign micromatrizz[0][393] = 9'b111111111;
assign micromatrizz[0][394] = 9'b111111111;
assign micromatrizz[0][395] = 9'b111111111;
assign micromatrizz[0][396] = 9'b111111111;
assign micromatrizz[0][397] = 9'b111111111;
assign micromatrizz[0][398] = 9'b111111111;
assign micromatrizz[0][399] = 9'b111111111;
assign micromatrizz[0][400] = 9'b111111111;
assign micromatrizz[0][401] = 9'b111111111;
assign micromatrizz[0][402] = 9'b111111111;
assign micromatrizz[0][403] = 9'b111111111;
assign micromatrizz[0][404] = 9'b111111111;
assign micromatrizz[0][405] = 9'b111111111;
assign micromatrizz[0][406] = 9'b111111111;
assign micromatrizz[0][407] = 9'b111111111;
assign micromatrizz[0][408] = 9'b111111111;
assign micromatrizz[0][409] = 9'b111111111;
assign micromatrizz[0][410] = 9'b111111111;
assign micromatrizz[0][411] = 9'b111111111;
assign micromatrizz[0][412] = 9'b111111111;
assign micromatrizz[0][413] = 9'b111111111;
assign micromatrizz[0][414] = 9'b111111111;
assign micromatrizz[0][415] = 9'b111111111;
assign micromatrizz[0][416] = 9'b111111111;
assign micromatrizz[0][417] = 9'b111111111;
assign micromatrizz[0][418] = 9'b111111111;
assign micromatrizz[0][419] = 9'b111111111;
assign micromatrizz[0][420] = 9'b111111111;
assign micromatrizz[0][421] = 9'b111111111;
assign micromatrizz[0][422] = 9'b111111111;
assign micromatrizz[0][423] = 9'b111111111;
assign micromatrizz[0][424] = 9'b111111111;
assign micromatrizz[0][425] = 9'b111111111;
assign micromatrizz[0][426] = 9'b111111111;
assign micromatrizz[0][427] = 9'b111111111;
assign micromatrizz[0][428] = 9'b111111111;
assign micromatrizz[0][429] = 9'b111111111;
assign micromatrizz[0][430] = 9'b111111111;
assign micromatrizz[0][431] = 9'b111111111;
assign micromatrizz[0][432] = 9'b111111111;
assign micromatrizz[0][433] = 9'b111111111;
assign micromatrizz[0][434] = 9'b111111111;
assign micromatrizz[0][435] = 9'b111111111;
assign micromatrizz[0][436] = 9'b111111111;
assign micromatrizz[0][437] = 9'b111111111;
assign micromatrizz[0][438] = 9'b111111111;
assign micromatrizz[0][439] = 9'b111111111;
assign micromatrizz[0][440] = 9'b111111111;
assign micromatrizz[0][441] = 9'b111111111;
assign micromatrizz[0][442] = 9'b111111111;
assign micromatrizz[0][443] = 9'b111111111;
assign micromatrizz[0][444] = 9'b111111111;
assign micromatrizz[0][445] = 9'b111111111;
assign micromatrizz[0][446] = 9'b111111111;
assign micromatrizz[0][447] = 9'b111111111;
assign micromatrizz[0][448] = 9'b111111111;
assign micromatrizz[0][449] = 9'b111111111;
assign micromatrizz[0][450] = 9'b111111111;
assign micromatrizz[0][451] = 9'b111111111;
assign micromatrizz[0][452] = 9'b111111111;
assign micromatrizz[0][453] = 9'b111111111;
assign micromatrizz[0][454] = 9'b111111111;
assign micromatrizz[0][455] = 9'b111111111;
assign micromatrizz[0][456] = 9'b111111111;
assign micromatrizz[0][457] = 9'b111111111;
assign micromatrizz[0][458] = 9'b111111111;
assign micromatrizz[0][459] = 9'b111111111;
assign micromatrizz[0][460] = 9'b111111111;
assign micromatrizz[0][461] = 9'b111111111;
assign micromatrizz[0][462] = 9'b111111111;
assign micromatrizz[0][463] = 9'b111111111;
assign micromatrizz[0][464] = 9'b111111111;
assign micromatrizz[0][465] = 9'b111111111;
assign micromatrizz[0][466] = 9'b111111111;
assign micromatrizz[0][467] = 9'b111111111;
assign micromatrizz[0][468] = 9'b111111111;
assign micromatrizz[0][469] = 9'b111111111;
assign micromatrizz[0][470] = 9'b111111111;
assign micromatrizz[0][471] = 9'b111111111;
assign micromatrizz[0][472] = 9'b111111111;
assign micromatrizz[0][473] = 9'b111111111;
assign micromatrizz[0][474] = 9'b111111111;
assign micromatrizz[0][475] = 9'b111111111;
assign micromatrizz[0][476] = 9'b111111111;
assign micromatrizz[0][477] = 9'b111111111;
assign micromatrizz[0][478] = 9'b111111111;
assign micromatrizz[0][479] = 9'b111111111;
assign micromatrizz[0][480] = 9'b111111111;
assign micromatrizz[0][481] = 9'b111111111;
assign micromatrizz[0][482] = 9'b111111111;
assign micromatrizz[0][483] = 9'b111111111;
assign micromatrizz[0][484] = 9'b111111111;
assign micromatrizz[0][485] = 9'b111111111;
assign micromatrizz[0][486] = 9'b111111111;
assign micromatrizz[0][487] = 9'b111111111;
assign micromatrizz[0][488] = 9'b111111111;
assign micromatrizz[0][489] = 9'b111111111;
assign micromatrizz[0][490] = 9'b111111111;
assign micromatrizz[0][491] = 9'b111111111;
assign micromatrizz[0][492] = 9'b111111111;
assign micromatrizz[0][493] = 9'b111111111;
assign micromatrizz[0][494] = 9'b111111111;
assign micromatrizz[0][495] = 9'b111111111;
assign micromatrizz[0][496] = 9'b111111111;
assign micromatrizz[0][497] = 9'b111111111;
assign micromatrizz[0][498] = 9'b111111111;
assign micromatrizz[0][499] = 9'b111111111;
assign micromatrizz[0][500] = 9'b111111111;
assign micromatrizz[0][501] = 9'b111111111;
assign micromatrizz[0][502] = 9'b111111111;
assign micromatrizz[0][503] = 9'b111111111;
assign micromatrizz[0][504] = 9'b111111111;
assign micromatrizz[0][505] = 9'b111111111;
assign micromatrizz[0][506] = 9'b111111111;
assign micromatrizz[0][507] = 9'b111111111;
assign micromatrizz[0][508] = 9'b111111111;
assign micromatrizz[0][509] = 9'b111111111;
assign micromatrizz[0][510] = 9'b111111111;
assign micromatrizz[0][511] = 9'b111111111;
assign micromatrizz[0][512] = 9'b111111111;
assign micromatrizz[0][513] = 9'b111111111;
assign micromatrizz[0][514] = 9'b111111111;
assign micromatrizz[0][515] = 9'b111111111;
assign micromatrizz[0][516] = 9'b111111111;
assign micromatrizz[0][517] = 9'b111111111;
assign micromatrizz[0][518] = 9'b111111111;
assign micromatrizz[0][519] = 9'b111111111;
assign micromatrizz[0][520] = 9'b111111111;
assign micromatrizz[0][521] = 9'b111111111;
assign micromatrizz[0][522] = 9'b111111111;
assign micromatrizz[0][523] = 9'b111111111;
assign micromatrizz[0][524] = 9'b111111111;
assign micromatrizz[0][525] = 9'b111111111;
assign micromatrizz[0][526] = 9'b111111111;
assign micromatrizz[0][527] = 9'b111111111;
assign micromatrizz[0][528] = 9'b111111111;
assign micromatrizz[0][529] = 9'b111111111;
assign micromatrizz[0][530] = 9'b111111111;
assign micromatrizz[0][531] = 9'b111111111;
assign micromatrizz[0][532] = 9'b111111111;
assign micromatrizz[0][533] = 9'b111111111;
assign micromatrizz[0][534] = 9'b111111111;
assign micromatrizz[0][535] = 9'b111111111;
assign micromatrizz[0][536] = 9'b111111111;
assign micromatrizz[0][537] = 9'b111111111;
assign micromatrizz[0][538] = 9'b111111111;
assign micromatrizz[0][539] = 9'b111111111;
assign micromatrizz[0][540] = 9'b111111111;
assign micromatrizz[0][541] = 9'b111111111;
assign micromatrizz[0][542] = 9'b111111111;
assign micromatrizz[0][543] = 9'b111111111;
assign micromatrizz[0][544] = 9'b111111111;
assign micromatrizz[0][545] = 9'b111111111;
assign micromatrizz[0][546] = 9'b111111111;
assign micromatrizz[0][547] = 9'b111111111;
assign micromatrizz[0][548] = 9'b111111111;
assign micromatrizz[0][549] = 9'b111111111;
assign micromatrizz[0][550] = 9'b111111111;
assign micromatrizz[0][551] = 9'b111111111;
assign micromatrizz[0][552] = 9'b111111111;
assign micromatrizz[0][553] = 9'b111111111;
assign micromatrizz[0][554] = 9'b111111111;
assign micromatrizz[0][555] = 9'b111111111;
assign micromatrizz[0][556] = 9'b111111111;
assign micromatrizz[0][557] = 9'b111111111;
assign micromatrizz[0][558] = 9'b111111111;
assign micromatrizz[0][559] = 9'b111111111;
assign micromatrizz[0][560] = 9'b111111111;
assign micromatrizz[0][561] = 9'b111111111;
assign micromatrizz[0][562] = 9'b111111111;
assign micromatrizz[0][563] = 9'b111111111;
assign micromatrizz[0][564] = 9'b111111111;
assign micromatrizz[0][565] = 9'b111111111;
assign micromatrizz[0][566] = 9'b111111111;
assign micromatrizz[0][567] = 9'b111111111;
assign micromatrizz[0][568] = 9'b111111111;
assign micromatrizz[0][569] = 9'b111111111;
assign micromatrizz[0][570] = 9'b111111111;
assign micromatrizz[0][571] = 9'b111111111;
assign micromatrizz[0][572] = 9'b111111111;
assign micromatrizz[0][573] = 9'b111111111;
assign micromatrizz[0][574] = 9'b111111111;
assign micromatrizz[0][575] = 9'b111111111;
assign micromatrizz[0][576] = 9'b111111111;
assign micromatrizz[0][577] = 9'b111111111;
assign micromatrizz[0][578] = 9'b111111111;
assign micromatrizz[0][579] = 9'b111111111;
assign micromatrizz[0][580] = 9'b111111111;
assign micromatrizz[0][581] = 9'b111111111;
assign micromatrizz[0][582] = 9'b111111111;
assign micromatrizz[0][583] = 9'b111111111;
assign micromatrizz[0][584] = 9'b111111111;
assign micromatrizz[0][585] = 9'b111111111;
assign micromatrizz[0][586] = 9'b111111111;
assign micromatrizz[0][587] = 9'b111111111;
assign micromatrizz[0][588] = 9'b111111111;
assign micromatrizz[0][589] = 9'b111111111;
assign micromatrizz[0][590] = 9'b111111111;
assign micromatrizz[0][591] = 9'b111111111;
assign micromatrizz[0][592] = 9'b111111111;
assign micromatrizz[0][593] = 9'b111111111;
assign micromatrizz[0][594] = 9'b111111111;
assign micromatrizz[0][595] = 9'b111111111;
assign micromatrizz[0][596] = 9'b111111111;
assign micromatrizz[0][597] = 9'b111111111;
assign micromatrizz[0][598] = 9'b111111111;
assign micromatrizz[0][599] = 9'b111111111;
assign micromatrizz[0][600] = 9'b111111111;
assign micromatrizz[0][601] = 9'b111111111;
assign micromatrizz[0][602] = 9'b111111111;
assign micromatrizz[0][603] = 9'b111111111;
assign micromatrizz[0][604] = 9'b111111111;
assign micromatrizz[0][605] = 9'b111111111;
assign micromatrizz[0][606] = 9'b111111111;
assign micromatrizz[0][607] = 9'b111111111;
assign micromatrizz[0][608] = 9'b111111111;
assign micromatrizz[0][609] = 9'b111111111;
assign micromatrizz[0][610] = 9'b111111111;
assign micromatrizz[0][611] = 9'b111111111;
assign micromatrizz[0][612] = 9'b111111111;
assign micromatrizz[0][613] = 9'b111111111;
assign micromatrizz[0][614] = 9'b111111111;
assign micromatrizz[0][615] = 9'b111111111;
assign micromatrizz[0][616] = 9'b111111111;
assign micromatrizz[0][617] = 9'b111111111;
assign micromatrizz[0][618] = 9'b111111111;
assign micromatrizz[0][619] = 9'b111111111;
assign micromatrizz[0][620] = 9'b111111111;
assign micromatrizz[0][621] = 9'b111111111;
assign micromatrizz[0][622] = 9'b111111111;
assign micromatrizz[0][623] = 9'b111111111;
assign micromatrizz[0][624] = 9'b111111111;
assign micromatrizz[0][625] = 9'b111111111;
assign micromatrizz[0][626] = 9'b111111111;
assign micromatrizz[0][627] = 9'b111111111;
assign micromatrizz[0][628] = 9'b111111111;
assign micromatrizz[0][629] = 9'b111111111;
assign micromatrizz[0][630] = 9'b111111111;
assign micromatrizz[0][631] = 9'b111111111;
assign micromatrizz[0][632] = 9'b111111111;
assign micromatrizz[0][633] = 9'b111111111;
assign micromatrizz[0][634] = 9'b111111111;
assign micromatrizz[0][635] = 9'b111111111;
assign micromatrizz[0][636] = 9'b111111111;
assign micromatrizz[0][637] = 9'b111111111;
assign micromatrizz[0][638] = 9'b111111111;
assign micromatrizz[0][639] = 9'b111111111;
assign micromatrizz[1][0] = 9'b111111111;
assign micromatrizz[1][1] = 9'b111111111;
assign micromatrizz[1][2] = 9'b111111111;
assign micromatrizz[1][3] = 9'b111111111;
assign micromatrizz[1][4] = 9'b111111111;
assign micromatrizz[1][5] = 9'b111111111;
assign micromatrizz[1][6] = 9'b111111111;
assign micromatrizz[1][7] = 9'b111111111;
assign micromatrizz[1][8] = 9'b111111111;
assign micromatrizz[1][9] = 9'b111111111;
assign micromatrizz[1][10] = 9'b111111111;
assign micromatrizz[1][11] = 9'b111111111;
assign micromatrizz[1][12] = 9'b111111111;
assign micromatrizz[1][13] = 9'b111111111;
assign micromatrizz[1][14] = 9'b111111111;
assign micromatrizz[1][15] = 9'b111111111;
assign micromatrizz[1][16] = 9'b111111111;
assign micromatrizz[1][17] = 9'b111111111;
assign micromatrizz[1][18] = 9'b111111111;
assign micromatrizz[1][19] = 9'b111111111;
assign micromatrizz[1][20] = 9'b111111111;
assign micromatrizz[1][21] = 9'b111111111;
assign micromatrizz[1][22] = 9'b111111111;
assign micromatrizz[1][23] = 9'b111111111;
assign micromatrizz[1][24] = 9'b111111111;
assign micromatrizz[1][25] = 9'b111111111;
assign micromatrizz[1][26] = 9'b111111111;
assign micromatrizz[1][27] = 9'b111111111;
assign micromatrizz[1][28] = 9'b111111111;
assign micromatrizz[1][29] = 9'b111111111;
assign micromatrizz[1][30] = 9'b111111111;
assign micromatrizz[1][31] = 9'b111111111;
assign micromatrizz[1][32] = 9'b111111111;
assign micromatrizz[1][33] = 9'b111111111;
assign micromatrizz[1][34] = 9'b111111111;
assign micromatrizz[1][35] = 9'b111111111;
assign micromatrizz[1][36] = 9'b111111111;
assign micromatrizz[1][37] = 9'b111111111;
assign micromatrizz[1][38] = 9'b111111111;
assign micromatrizz[1][39] = 9'b111111111;
assign micromatrizz[1][40] = 9'b111111111;
assign micromatrizz[1][41] = 9'b111111111;
assign micromatrizz[1][42] = 9'b111111111;
assign micromatrizz[1][43] = 9'b111111111;
assign micromatrizz[1][44] = 9'b111111111;
assign micromatrizz[1][45] = 9'b111111111;
assign micromatrizz[1][46] = 9'b111111111;
assign micromatrizz[1][47] = 9'b111111111;
assign micromatrizz[1][48] = 9'b111111111;
assign micromatrizz[1][49] = 9'b111111111;
assign micromatrizz[1][50] = 9'b111111111;
assign micromatrizz[1][51] = 9'b111111111;
assign micromatrizz[1][52] = 9'b111111111;
assign micromatrizz[1][53] = 9'b111111111;
assign micromatrizz[1][54] = 9'b111111111;
assign micromatrizz[1][55] = 9'b111111111;
assign micromatrizz[1][56] = 9'b111111111;
assign micromatrizz[1][57] = 9'b111111111;
assign micromatrizz[1][58] = 9'b111111111;
assign micromatrizz[1][59] = 9'b111111111;
assign micromatrizz[1][60] = 9'b111111111;
assign micromatrizz[1][61] = 9'b111111111;
assign micromatrizz[1][62] = 9'b111111111;
assign micromatrizz[1][63] = 9'b111111111;
assign micromatrizz[1][64] = 9'b111111111;
assign micromatrizz[1][65] = 9'b111111111;
assign micromatrizz[1][66] = 9'b111111111;
assign micromatrizz[1][67] = 9'b111111111;
assign micromatrizz[1][68] = 9'b111111111;
assign micromatrizz[1][69] = 9'b111111111;
assign micromatrizz[1][70] = 9'b111111111;
assign micromatrizz[1][71] = 9'b111111111;
assign micromatrizz[1][72] = 9'b111111111;
assign micromatrizz[1][73] = 9'b111111111;
assign micromatrizz[1][74] = 9'b111111111;
assign micromatrizz[1][75] = 9'b111111111;
assign micromatrizz[1][76] = 9'b111111111;
assign micromatrizz[1][77] = 9'b111111111;
assign micromatrizz[1][78] = 9'b111111111;
assign micromatrizz[1][79] = 9'b111111111;
assign micromatrizz[1][80] = 9'b111111111;
assign micromatrizz[1][81] = 9'b111111111;
assign micromatrizz[1][82] = 9'b111111111;
assign micromatrizz[1][83] = 9'b111111111;
assign micromatrizz[1][84] = 9'b111111111;
assign micromatrizz[1][85] = 9'b111111111;
assign micromatrizz[1][86] = 9'b111111111;
assign micromatrizz[1][87] = 9'b111111111;
assign micromatrizz[1][88] = 9'b111111111;
assign micromatrizz[1][89] = 9'b111111111;
assign micromatrizz[1][90] = 9'b111111111;
assign micromatrizz[1][91] = 9'b111111111;
assign micromatrizz[1][92] = 9'b111111111;
assign micromatrizz[1][93] = 9'b111111111;
assign micromatrizz[1][94] = 9'b111111111;
assign micromatrizz[1][95] = 9'b111111111;
assign micromatrizz[1][96] = 9'b111111111;
assign micromatrizz[1][97] = 9'b111111111;
assign micromatrizz[1][98] = 9'b111111111;
assign micromatrizz[1][99] = 9'b111111111;
assign micromatrizz[1][100] = 9'b111111111;
assign micromatrizz[1][101] = 9'b111111111;
assign micromatrizz[1][102] = 9'b111111111;
assign micromatrizz[1][103] = 9'b111111111;
assign micromatrizz[1][104] = 9'b111111111;
assign micromatrizz[1][105] = 9'b111111111;
assign micromatrizz[1][106] = 9'b111111111;
assign micromatrizz[1][107] = 9'b111111111;
assign micromatrizz[1][108] = 9'b111111111;
assign micromatrizz[1][109] = 9'b111111111;
assign micromatrizz[1][110] = 9'b111111111;
assign micromatrizz[1][111] = 9'b111111111;
assign micromatrizz[1][112] = 9'b111111111;
assign micromatrizz[1][113] = 9'b111111111;
assign micromatrizz[1][114] = 9'b111111111;
assign micromatrizz[1][115] = 9'b111111111;
assign micromatrizz[1][116] = 9'b111111111;
assign micromatrizz[1][117] = 9'b111111111;
assign micromatrizz[1][118] = 9'b111111111;
assign micromatrizz[1][119] = 9'b111111111;
assign micromatrizz[1][120] = 9'b111111111;
assign micromatrizz[1][121] = 9'b111111111;
assign micromatrizz[1][122] = 9'b111111111;
assign micromatrizz[1][123] = 9'b111111111;
assign micromatrizz[1][124] = 9'b111111111;
assign micromatrizz[1][125] = 9'b111111111;
assign micromatrizz[1][126] = 9'b111111111;
assign micromatrizz[1][127] = 9'b111111111;
assign micromatrizz[1][128] = 9'b111111111;
assign micromatrizz[1][129] = 9'b111111111;
assign micromatrizz[1][130] = 9'b111111111;
assign micromatrizz[1][131] = 9'b111111111;
assign micromatrizz[1][132] = 9'b111111111;
assign micromatrizz[1][133] = 9'b111111111;
assign micromatrizz[1][134] = 9'b111111111;
assign micromatrizz[1][135] = 9'b111111111;
assign micromatrizz[1][136] = 9'b111111111;
assign micromatrizz[1][137] = 9'b111111111;
assign micromatrizz[1][138] = 9'b111111111;
assign micromatrizz[1][139] = 9'b111111111;
assign micromatrizz[1][140] = 9'b111111111;
assign micromatrizz[1][141] = 9'b111111111;
assign micromatrizz[1][142] = 9'b111111111;
assign micromatrizz[1][143] = 9'b111111111;
assign micromatrizz[1][144] = 9'b111111111;
assign micromatrizz[1][145] = 9'b111111111;
assign micromatrizz[1][146] = 9'b111111111;
assign micromatrizz[1][147] = 9'b111111111;
assign micromatrizz[1][148] = 9'b111111111;
assign micromatrizz[1][149] = 9'b111111111;
assign micromatrizz[1][150] = 9'b111111111;
assign micromatrizz[1][151] = 9'b111111111;
assign micromatrizz[1][152] = 9'b111111111;
assign micromatrizz[1][153] = 9'b111111111;
assign micromatrizz[1][154] = 9'b111111111;
assign micromatrizz[1][155] = 9'b111111111;
assign micromatrizz[1][156] = 9'b111111111;
assign micromatrizz[1][157] = 9'b111111111;
assign micromatrizz[1][158] = 9'b111111111;
assign micromatrizz[1][159] = 9'b111111111;
assign micromatrizz[1][160] = 9'b111111111;
assign micromatrizz[1][161] = 9'b111111111;
assign micromatrizz[1][162] = 9'b111111111;
assign micromatrizz[1][163] = 9'b111111111;
assign micromatrizz[1][164] = 9'b111111111;
assign micromatrizz[1][165] = 9'b111111111;
assign micromatrizz[1][166] = 9'b111111111;
assign micromatrizz[1][167] = 9'b111111111;
assign micromatrizz[1][168] = 9'b111111111;
assign micromatrizz[1][169] = 9'b111111111;
assign micromatrizz[1][170] = 9'b111111111;
assign micromatrizz[1][171] = 9'b111111111;
assign micromatrizz[1][172] = 9'b111111111;
assign micromatrizz[1][173] = 9'b111111111;
assign micromatrizz[1][174] = 9'b111111111;
assign micromatrizz[1][175] = 9'b111111111;
assign micromatrizz[1][176] = 9'b111111111;
assign micromatrizz[1][177] = 9'b111111111;
assign micromatrizz[1][178] = 9'b111111111;
assign micromatrizz[1][179] = 9'b111111111;
assign micromatrizz[1][180] = 9'b111111111;
assign micromatrizz[1][181] = 9'b111111111;
assign micromatrizz[1][182] = 9'b111111111;
assign micromatrizz[1][183] = 9'b111111111;
assign micromatrizz[1][184] = 9'b111111111;
assign micromatrizz[1][185] = 9'b111111111;
assign micromatrizz[1][186] = 9'b111111111;
assign micromatrizz[1][187] = 9'b111111111;
assign micromatrizz[1][188] = 9'b111111111;
assign micromatrizz[1][189] = 9'b111111111;
assign micromatrizz[1][190] = 9'b111111111;
assign micromatrizz[1][191] = 9'b111111111;
assign micromatrizz[1][192] = 9'b111111111;
assign micromatrizz[1][193] = 9'b111111111;
assign micromatrizz[1][194] = 9'b111111111;
assign micromatrizz[1][195] = 9'b111111111;
assign micromatrizz[1][196] = 9'b111111111;
assign micromatrizz[1][197] = 9'b111111111;
assign micromatrizz[1][198] = 9'b111111111;
assign micromatrizz[1][199] = 9'b111111111;
assign micromatrizz[1][200] = 9'b111111111;
assign micromatrizz[1][201] = 9'b111111111;
assign micromatrizz[1][202] = 9'b111111111;
assign micromatrizz[1][203] = 9'b111111111;
assign micromatrizz[1][204] = 9'b111111111;
assign micromatrizz[1][205] = 9'b111111111;
assign micromatrizz[1][206] = 9'b111111111;
assign micromatrizz[1][207] = 9'b111111111;
assign micromatrizz[1][208] = 9'b111111111;
assign micromatrizz[1][209] = 9'b111111111;
assign micromatrizz[1][210] = 9'b111111111;
assign micromatrizz[1][211] = 9'b111111111;
assign micromatrizz[1][212] = 9'b111111111;
assign micromatrizz[1][213] = 9'b111111111;
assign micromatrizz[1][214] = 9'b111111111;
assign micromatrizz[1][215] = 9'b111111111;
assign micromatrizz[1][216] = 9'b111111111;
assign micromatrizz[1][217] = 9'b111111111;
assign micromatrizz[1][218] = 9'b111111111;
assign micromatrizz[1][219] = 9'b111111111;
assign micromatrizz[1][220] = 9'b111111111;
assign micromatrizz[1][221] = 9'b111111111;
assign micromatrizz[1][222] = 9'b111111111;
assign micromatrizz[1][223] = 9'b111111111;
assign micromatrizz[1][224] = 9'b111111111;
assign micromatrizz[1][225] = 9'b111111111;
assign micromatrizz[1][226] = 9'b111111111;
assign micromatrizz[1][227] = 9'b111111111;
assign micromatrizz[1][228] = 9'b111111111;
assign micromatrizz[1][229] = 9'b111111111;
assign micromatrizz[1][230] = 9'b111111111;
assign micromatrizz[1][231] = 9'b111111111;
assign micromatrizz[1][232] = 9'b111111111;
assign micromatrizz[1][233] = 9'b111111111;
assign micromatrizz[1][234] = 9'b111111111;
assign micromatrizz[1][235] = 9'b111111111;
assign micromatrizz[1][236] = 9'b111111111;
assign micromatrizz[1][237] = 9'b111111111;
assign micromatrizz[1][238] = 9'b111111111;
assign micromatrizz[1][239] = 9'b111111111;
assign micromatrizz[1][240] = 9'b111111111;
assign micromatrizz[1][241] = 9'b111111111;
assign micromatrizz[1][242] = 9'b111111111;
assign micromatrizz[1][243] = 9'b111111111;
assign micromatrizz[1][244] = 9'b111111111;
assign micromatrizz[1][245] = 9'b111111111;
assign micromatrizz[1][246] = 9'b111111111;
assign micromatrizz[1][247] = 9'b111111111;
assign micromatrizz[1][248] = 9'b111111111;
assign micromatrizz[1][249] = 9'b111111111;
assign micromatrizz[1][250] = 9'b111111111;
assign micromatrizz[1][251] = 9'b111111111;
assign micromatrizz[1][252] = 9'b111111111;
assign micromatrizz[1][253] = 9'b111111111;
assign micromatrizz[1][254] = 9'b111111111;
assign micromatrizz[1][255] = 9'b111111111;
assign micromatrizz[1][256] = 9'b111111111;
assign micromatrizz[1][257] = 9'b111111111;
assign micromatrizz[1][258] = 9'b111111111;
assign micromatrizz[1][259] = 9'b111111111;
assign micromatrizz[1][260] = 9'b111111111;
assign micromatrizz[1][261] = 9'b111111111;
assign micromatrizz[1][262] = 9'b111111111;
assign micromatrizz[1][263] = 9'b111111111;
assign micromatrizz[1][264] = 9'b111111111;
assign micromatrizz[1][265] = 9'b111111111;
assign micromatrizz[1][266] = 9'b111111111;
assign micromatrizz[1][267] = 9'b111111111;
assign micromatrizz[1][268] = 9'b111111111;
assign micromatrizz[1][269] = 9'b111111111;
assign micromatrizz[1][270] = 9'b111111111;
assign micromatrizz[1][271] = 9'b111111111;
assign micromatrizz[1][272] = 9'b111111111;
assign micromatrizz[1][273] = 9'b111111111;
assign micromatrizz[1][274] = 9'b111111111;
assign micromatrizz[1][275] = 9'b111111111;
assign micromatrizz[1][276] = 9'b111111111;
assign micromatrizz[1][277] = 9'b111111111;
assign micromatrizz[1][278] = 9'b111111111;
assign micromatrizz[1][279] = 9'b111111111;
assign micromatrizz[1][280] = 9'b111111111;
assign micromatrizz[1][281] = 9'b111111111;
assign micromatrizz[1][282] = 9'b111111111;
assign micromatrizz[1][283] = 9'b111111111;
assign micromatrizz[1][284] = 9'b111111111;
assign micromatrizz[1][285] = 9'b111111111;
assign micromatrizz[1][286] = 9'b111111111;
assign micromatrizz[1][287] = 9'b111111111;
assign micromatrizz[1][288] = 9'b111111111;
assign micromatrizz[1][289] = 9'b111111111;
assign micromatrizz[1][290] = 9'b111111111;
assign micromatrizz[1][291] = 9'b111111111;
assign micromatrizz[1][292] = 9'b111111111;
assign micromatrizz[1][293] = 9'b111111111;
assign micromatrizz[1][294] = 9'b111111111;
assign micromatrizz[1][295] = 9'b111111111;
assign micromatrizz[1][296] = 9'b111111111;
assign micromatrizz[1][297] = 9'b111111111;
assign micromatrizz[1][298] = 9'b111111111;
assign micromatrizz[1][299] = 9'b111111111;
assign micromatrizz[1][300] = 9'b111111111;
assign micromatrizz[1][301] = 9'b111111111;
assign micromatrizz[1][302] = 9'b111111111;
assign micromatrizz[1][303] = 9'b111111111;
assign micromatrizz[1][304] = 9'b111111111;
assign micromatrizz[1][305] = 9'b111111111;
assign micromatrizz[1][306] = 9'b111111111;
assign micromatrizz[1][307] = 9'b111111111;
assign micromatrizz[1][308] = 9'b111111111;
assign micromatrizz[1][309] = 9'b111111111;
assign micromatrizz[1][310] = 9'b111111111;
assign micromatrizz[1][311] = 9'b111111111;
assign micromatrizz[1][312] = 9'b111111111;
assign micromatrizz[1][313] = 9'b111111111;
assign micromatrizz[1][314] = 9'b111111111;
assign micromatrizz[1][315] = 9'b111111111;
assign micromatrizz[1][316] = 9'b111111111;
assign micromatrizz[1][317] = 9'b111111111;
assign micromatrizz[1][318] = 9'b111111111;
assign micromatrizz[1][319] = 9'b111111111;
assign micromatrizz[1][320] = 9'b111111111;
assign micromatrizz[1][321] = 9'b111111111;
assign micromatrizz[1][322] = 9'b111111111;
assign micromatrizz[1][323] = 9'b111111111;
assign micromatrizz[1][324] = 9'b111111111;
assign micromatrizz[1][325] = 9'b111111111;
assign micromatrizz[1][326] = 9'b111111111;
assign micromatrizz[1][327] = 9'b111111111;
assign micromatrizz[1][328] = 9'b111111111;
assign micromatrizz[1][329] = 9'b111111111;
assign micromatrizz[1][330] = 9'b111111111;
assign micromatrizz[1][331] = 9'b111111111;
assign micromatrizz[1][332] = 9'b111111111;
assign micromatrizz[1][333] = 9'b111111111;
assign micromatrizz[1][334] = 9'b111111111;
assign micromatrizz[1][335] = 9'b111111111;
assign micromatrizz[1][336] = 9'b111111111;
assign micromatrizz[1][337] = 9'b111111111;
assign micromatrizz[1][338] = 9'b111111111;
assign micromatrizz[1][339] = 9'b111111111;
assign micromatrizz[1][340] = 9'b111111111;
assign micromatrizz[1][341] = 9'b111111111;
assign micromatrizz[1][342] = 9'b111111111;
assign micromatrizz[1][343] = 9'b111111111;
assign micromatrizz[1][344] = 9'b111111111;
assign micromatrizz[1][345] = 9'b111111111;
assign micromatrizz[1][346] = 9'b111111111;
assign micromatrizz[1][347] = 9'b111111111;
assign micromatrizz[1][348] = 9'b111111111;
assign micromatrizz[1][349] = 9'b111111111;
assign micromatrizz[1][350] = 9'b111111111;
assign micromatrizz[1][351] = 9'b111111111;
assign micromatrizz[1][352] = 9'b111111111;
assign micromatrizz[1][353] = 9'b111111111;
assign micromatrizz[1][354] = 9'b111111111;
assign micromatrizz[1][355] = 9'b111111111;
assign micromatrizz[1][356] = 9'b111111111;
assign micromatrizz[1][357] = 9'b111111111;
assign micromatrizz[1][358] = 9'b111111111;
assign micromatrizz[1][359] = 9'b111111111;
assign micromatrizz[1][360] = 9'b111111111;
assign micromatrizz[1][361] = 9'b111111111;
assign micromatrizz[1][362] = 9'b111111111;
assign micromatrizz[1][363] = 9'b111111111;
assign micromatrizz[1][364] = 9'b111111111;
assign micromatrizz[1][365] = 9'b111111111;
assign micromatrizz[1][366] = 9'b111111111;
assign micromatrizz[1][367] = 9'b111111111;
assign micromatrizz[1][368] = 9'b111111111;
assign micromatrizz[1][369] = 9'b111111111;
assign micromatrizz[1][370] = 9'b111111111;
assign micromatrizz[1][371] = 9'b111111111;
assign micromatrizz[1][372] = 9'b111111111;
assign micromatrizz[1][373] = 9'b111111111;
assign micromatrizz[1][374] = 9'b111111111;
assign micromatrizz[1][375] = 9'b111111111;
assign micromatrizz[1][376] = 9'b111111111;
assign micromatrizz[1][377] = 9'b111111111;
assign micromatrizz[1][378] = 9'b111111111;
assign micromatrizz[1][379] = 9'b111111111;
assign micromatrizz[1][380] = 9'b111111111;
assign micromatrizz[1][381] = 9'b111111111;
assign micromatrizz[1][382] = 9'b111111111;
assign micromatrizz[1][383] = 9'b111111111;
assign micromatrizz[1][384] = 9'b111111111;
assign micromatrizz[1][385] = 9'b111111111;
assign micromatrizz[1][386] = 9'b111111111;
assign micromatrizz[1][387] = 9'b111111111;
assign micromatrizz[1][388] = 9'b111111111;
assign micromatrizz[1][389] = 9'b111111111;
assign micromatrizz[1][390] = 9'b111111111;
assign micromatrizz[1][391] = 9'b111111111;
assign micromatrizz[1][392] = 9'b111111111;
assign micromatrizz[1][393] = 9'b111111111;
assign micromatrizz[1][394] = 9'b111111111;
assign micromatrizz[1][395] = 9'b111111111;
assign micromatrizz[1][396] = 9'b111111111;
assign micromatrizz[1][397] = 9'b111111111;
assign micromatrizz[1][398] = 9'b111111111;
assign micromatrizz[1][399] = 9'b111111111;
assign micromatrizz[1][400] = 9'b111111111;
assign micromatrizz[1][401] = 9'b111111111;
assign micromatrizz[1][402] = 9'b111111111;
assign micromatrizz[1][403] = 9'b111111111;
assign micromatrizz[1][404] = 9'b111111111;
assign micromatrizz[1][405] = 9'b111111111;
assign micromatrizz[1][406] = 9'b111111111;
assign micromatrizz[1][407] = 9'b111111111;
assign micromatrizz[1][408] = 9'b111111111;
assign micromatrizz[1][409] = 9'b111111111;
assign micromatrizz[1][410] = 9'b111111111;
assign micromatrizz[1][411] = 9'b111111111;
assign micromatrizz[1][412] = 9'b111111111;
assign micromatrizz[1][413] = 9'b111111111;
assign micromatrizz[1][414] = 9'b111111111;
assign micromatrizz[1][415] = 9'b111111111;
assign micromatrizz[1][416] = 9'b111111111;
assign micromatrizz[1][417] = 9'b111111111;
assign micromatrizz[1][418] = 9'b111111111;
assign micromatrizz[1][419] = 9'b111111111;
assign micromatrizz[1][420] = 9'b111111111;
assign micromatrizz[1][421] = 9'b111111111;
assign micromatrizz[1][422] = 9'b111111111;
assign micromatrizz[1][423] = 9'b111111111;
assign micromatrizz[1][424] = 9'b111111111;
assign micromatrizz[1][425] = 9'b111111111;
assign micromatrizz[1][426] = 9'b111111111;
assign micromatrizz[1][427] = 9'b111111111;
assign micromatrizz[1][428] = 9'b111111111;
assign micromatrizz[1][429] = 9'b111111111;
assign micromatrizz[1][430] = 9'b111111111;
assign micromatrizz[1][431] = 9'b111111111;
assign micromatrizz[1][432] = 9'b111111111;
assign micromatrizz[1][433] = 9'b111111111;
assign micromatrizz[1][434] = 9'b111111111;
assign micromatrizz[1][435] = 9'b111111111;
assign micromatrizz[1][436] = 9'b111111111;
assign micromatrizz[1][437] = 9'b111111111;
assign micromatrizz[1][438] = 9'b111111111;
assign micromatrizz[1][439] = 9'b111111111;
assign micromatrizz[1][440] = 9'b111111111;
assign micromatrizz[1][441] = 9'b111111111;
assign micromatrizz[1][442] = 9'b111111111;
assign micromatrizz[1][443] = 9'b111111111;
assign micromatrizz[1][444] = 9'b111111111;
assign micromatrizz[1][445] = 9'b111111111;
assign micromatrizz[1][446] = 9'b111111111;
assign micromatrizz[1][447] = 9'b111111111;
assign micromatrizz[1][448] = 9'b111111111;
assign micromatrizz[1][449] = 9'b111111111;
assign micromatrizz[1][450] = 9'b111111111;
assign micromatrizz[1][451] = 9'b111111111;
assign micromatrizz[1][452] = 9'b111111111;
assign micromatrizz[1][453] = 9'b111111111;
assign micromatrizz[1][454] = 9'b111111111;
assign micromatrizz[1][455] = 9'b111111111;
assign micromatrizz[1][456] = 9'b111111111;
assign micromatrizz[1][457] = 9'b111111111;
assign micromatrizz[1][458] = 9'b111111111;
assign micromatrizz[1][459] = 9'b111111111;
assign micromatrizz[1][460] = 9'b111111111;
assign micromatrizz[1][461] = 9'b111111111;
assign micromatrizz[1][462] = 9'b111111111;
assign micromatrizz[1][463] = 9'b111111111;
assign micromatrizz[1][464] = 9'b111111111;
assign micromatrizz[1][465] = 9'b111111111;
assign micromatrizz[1][466] = 9'b111111111;
assign micromatrizz[1][467] = 9'b111111111;
assign micromatrizz[1][468] = 9'b111111111;
assign micromatrizz[1][469] = 9'b111111111;
assign micromatrizz[1][470] = 9'b111111111;
assign micromatrizz[1][471] = 9'b111111111;
assign micromatrizz[1][472] = 9'b111111111;
assign micromatrizz[1][473] = 9'b111111111;
assign micromatrizz[1][474] = 9'b111111111;
assign micromatrizz[1][475] = 9'b111111111;
assign micromatrizz[1][476] = 9'b111111111;
assign micromatrizz[1][477] = 9'b111111111;
assign micromatrizz[1][478] = 9'b111111111;
assign micromatrizz[1][479] = 9'b111111111;
assign micromatrizz[1][480] = 9'b111111111;
assign micromatrizz[1][481] = 9'b111111111;
assign micromatrizz[1][482] = 9'b111111111;
assign micromatrizz[1][483] = 9'b111111111;
assign micromatrizz[1][484] = 9'b111111111;
assign micromatrizz[1][485] = 9'b111111111;
assign micromatrizz[1][486] = 9'b111111111;
assign micromatrizz[1][487] = 9'b111111111;
assign micromatrizz[1][488] = 9'b111111111;
assign micromatrizz[1][489] = 9'b111111111;
assign micromatrizz[1][490] = 9'b111111111;
assign micromatrizz[1][491] = 9'b111111111;
assign micromatrizz[1][492] = 9'b111111111;
assign micromatrizz[1][493] = 9'b111111111;
assign micromatrizz[1][494] = 9'b111111111;
assign micromatrizz[1][495] = 9'b111111111;
assign micromatrizz[1][496] = 9'b111111111;
assign micromatrizz[1][497] = 9'b111111111;
assign micromatrizz[1][498] = 9'b111111111;
assign micromatrizz[1][499] = 9'b111111111;
assign micromatrizz[1][500] = 9'b111111111;
assign micromatrizz[1][501] = 9'b111111111;
assign micromatrizz[1][502] = 9'b111111111;
assign micromatrizz[1][503] = 9'b111111111;
assign micromatrizz[1][504] = 9'b111111111;
assign micromatrizz[1][505] = 9'b111111111;
assign micromatrizz[1][506] = 9'b111111111;
assign micromatrizz[1][507] = 9'b111111111;
assign micromatrizz[1][508] = 9'b111111111;
assign micromatrizz[1][509] = 9'b111111111;
assign micromatrizz[1][510] = 9'b111111111;
assign micromatrizz[1][511] = 9'b111111111;
assign micromatrizz[1][512] = 9'b111111111;
assign micromatrizz[1][513] = 9'b111111111;
assign micromatrizz[1][514] = 9'b111111111;
assign micromatrizz[1][515] = 9'b111111111;
assign micromatrizz[1][516] = 9'b111111111;
assign micromatrizz[1][517] = 9'b111111111;
assign micromatrizz[1][518] = 9'b111111111;
assign micromatrizz[1][519] = 9'b111111111;
assign micromatrizz[1][520] = 9'b111111111;
assign micromatrizz[1][521] = 9'b111111111;
assign micromatrizz[1][522] = 9'b111111111;
assign micromatrizz[1][523] = 9'b111111111;
assign micromatrizz[1][524] = 9'b111111111;
assign micromatrizz[1][525] = 9'b111111111;
assign micromatrizz[1][526] = 9'b111111111;
assign micromatrizz[1][527] = 9'b111111111;
assign micromatrizz[1][528] = 9'b111111111;
assign micromatrizz[1][529] = 9'b111111111;
assign micromatrizz[1][530] = 9'b111111111;
assign micromatrizz[1][531] = 9'b111111111;
assign micromatrizz[1][532] = 9'b111111111;
assign micromatrizz[1][533] = 9'b111111111;
assign micromatrizz[1][534] = 9'b111111111;
assign micromatrizz[1][535] = 9'b111111111;
assign micromatrizz[1][536] = 9'b111111111;
assign micromatrizz[1][537] = 9'b111111111;
assign micromatrizz[1][538] = 9'b111111111;
assign micromatrizz[1][539] = 9'b111111111;
assign micromatrizz[1][540] = 9'b111111111;
assign micromatrizz[1][541] = 9'b111111111;
assign micromatrizz[1][542] = 9'b111111111;
assign micromatrizz[1][543] = 9'b111111111;
assign micromatrizz[1][544] = 9'b111111111;
assign micromatrizz[1][545] = 9'b111111111;
assign micromatrizz[1][546] = 9'b111111111;
assign micromatrizz[1][547] = 9'b111111111;
assign micromatrizz[1][548] = 9'b111111111;
assign micromatrizz[1][549] = 9'b111111111;
assign micromatrizz[1][550] = 9'b111111111;
assign micromatrizz[1][551] = 9'b111111111;
assign micromatrizz[1][552] = 9'b111111111;
assign micromatrizz[1][553] = 9'b111111111;
assign micromatrizz[1][554] = 9'b111111111;
assign micromatrizz[1][555] = 9'b111111111;
assign micromatrizz[1][556] = 9'b111111111;
assign micromatrizz[1][557] = 9'b111111111;
assign micromatrizz[1][558] = 9'b111111111;
assign micromatrizz[1][559] = 9'b111111111;
assign micromatrizz[1][560] = 9'b111111111;
assign micromatrizz[1][561] = 9'b111111111;
assign micromatrizz[1][562] = 9'b111111111;
assign micromatrizz[1][563] = 9'b111111111;
assign micromatrizz[1][564] = 9'b111111111;
assign micromatrizz[1][565] = 9'b111111111;
assign micromatrizz[1][566] = 9'b111111111;
assign micromatrizz[1][567] = 9'b111111111;
assign micromatrizz[1][568] = 9'b111111111;
assign micromatrizz[1][569] = 9'b111111111;
assign micromatrizz[1][570] = 9'b111111111;
assign micromatrizz[1][571] = 9'b111111111;
assign micromatrizz[1][572] = 9'b111111111;
assign micromatrizz[1][573] = 9'b111111111;
assign micromatrizz[1][574] = 9'b111111111;
assign micromatrizz[1][575] = 9'b111111111;
assign micromatrizz[1][576] = 9'b111111111;
assign micromatrizz[1][577] = 9'b111111111;
assign micromatrizz[1][578] = 9'b111111111;
assign micromatrizz[1][579] = 9'b111111111;
assign micromatrizz[1][580] = 9'b111111111;
assign micromatrizz[1][581] = 9'b111111111;
assign micromatrizz[1][582] = 9'b111111111;
assign micromatrizz[1][583] = 9'b111111111;
assign micromatrizz[1][584] = 9'b111111111;
assign micromatrizz[1][585] = 9'b111111111;
assign micromatrizz[1][586] = 9'b111111111;
assign micromatrizz[1][587] = 9'b111111111;
assign micromatrizz[1][588] = 9'b111111111;
assign micromatrizz[1][589] = 9'b111111111;
assign micromatrizz[1][590] = 9'b111111111;
assign micromatrizz[1][591] = 9'b111111111;
assign micromatrizz[1][592] = 9'b111111111;
assign micromatrizz[1][593] = 9'b111111111;
assign micromatrizz[1][594] = 9'b111111111;
assign micromatrizz[1][595] = 9'b111111111;
assign micromatrizz[1][596] = 9'b111111111;
assign micromatrizz[1][597] = 9'b111111111;
assign micromatrizz[1][598] = 9'b111111111;
assign micromatrizz[1][599] = 9'b111111111;
assign micromatrizz[1][600] = 9'b111111111;
assign micromatrizz[1][601] = 9'b111111111;
assign micromatrizz[1][602] = 9'b111111111;
assign micromatrizz[1][603] = 9'b111111111;
assign micromatrizz[1][604] = 9'b111111111;
assign micromatrizz[1][605] = 9'b111111111;
assign micromatrizz[1][606] = 9'b111111111;
assign micromatrizz[1][607] = 9'b111111111;
assign micromatrizz[1][608] = 9'b111111111;
assign micromatrizz[1][609] = 9'b111111111;
assign micromatrizz[1][610] = 9'b111111111;
assign micromatrizz[1][611] = 9'b111111111;
assign micromatrizz[1][612] = 9'b111111111;
assign micromatrizz[1][613] = 9'b111111111;
assign micromatrizz[1][614] = 9'b111111111;
assign micromatrizz[1][615] = 9'b111111111;
assign micromatrizz[1][616] = 9'b111111111;
assign micromatrizz[1][617] = 9'b111111111;
assign micromatrizz[1][618] = 9'b111111111;
assign micromatrizz[1][619] = 9'b111111111;
assign micromatrizz[1][620] = 9'b111111111;
assign micromatrizz[1][621] = 9'b111111111;
assign micromatrizz[1][622] = 9'b111111111;
assign micromatrizz[1][623] = 9'b111111111;
assign micromatrizz[1][624] = 9'b111111111;
assign micromatrizz[1][625] = 9'b111111111;
assign micromatrizz[1][626] = 9'b111111111;
assign micromatrizz[1][627] = 9'b111111111;
assign micromatrizz[1][628] = 9'b111111111;
assign micromatrizz[1][629] = 9'b111111111;
assign micromatrizz[1][630] = 9'b111111111;
assign micromatrizz[1][631] = 9'b111111111;
assign micromatrizz[1][632] = 9'b111111111;
assign micromatrizz[1][633] = 9'b111111111;
assign micromatrizz[1][634] = 9'b111111111;
assign micromatrizz[1][635] = 9'b111111111;
assign micromatrizz[1][636] = 9'b111111111;
assign micromatrizz[1][637] = 9'b111111111;
assign micromatrizz[1][638] = 9'b111111111;
assign micromatrizz[1][639] = 9'b111111111;
assign micromatrizz[2][0] = 9'b111111111;
assign micromatrizz[2][1] = 9'b111111111;
assign micromatrizz[2][2] = 9'b111111111;
assign micromatrizz[2][3] = 9'b111111111;
assign micromatrizz[2][4] = 9'b111111111;
assign micromatrizz[2][5] = 9'b111111111;
assign micromatrizz[2][6] = 9'b111111111;
assign micromatrizz[2][7] = 9'b111111111;
assign micromatrizz[2][8] = 9'b111111111;
assign micromatrizz[2][9] = 9'b111111111;
assign micromatrizz[2][10] = 9'b111111111;
assign micromatrizz[2][11] = 9'b111111111;
assign micromatrizz[2][12] = 9'b111111111;
assign micromatrizz[2][13] = 9'b111111111;
assign micromatrizz[2][14] = 9'b111111111;
assign micromatrizz[2][15] = 9'b111111111;
assign micromatrizz[2][16] = 9'b111111111;
assign micromatrizz[2][17] = 9'b111111111;
assign micromatrizz[2][18] = 9'b111111111;
assign micromatrizz[2][19] = 9'b111111111;
assign micromatrizz[2][20] = 9'b111111111;
assign micromatrizz[2][21] = 9'b111111111;
assign micromatrizz[2][22] = 9'b111111111;
assign micromatrizz[2][23] = 9'b111111111;
assign micromatrizz[2][24] = 9'b111111111;
assign micromatrizz[2][25] = 9'b111111111;
assign micromatrizz[2][26] = 9'b111111111;
assign micromatrizz[2][27] = 9'b111111111;
assign micromatrizz[2][28] = 9'b111111111;
assign micromatrizz[2][29] = 9'b111111111;
assign micromatrizz[2][30] = 9'b111111111;
assign micromatrizz[2][31] = 9'b111111111;
assign micromatrizz[2][32] = 9'b111111111;
assign micromatrizz[2][33] = 9'b111111111;
assign micromatrizz[2][34] = 9'b111111111;
assign micromatrizz[2][35] = 9'b111111111;
assign micromatrizz[2][36] = 9'b111111111;
assign micromatrizz[2][37] = 9'b111111111;
assign micromatrizz[2][38] = 9'b111111111;
assign micromatrizz[2][39] = 9'b111111111;
assign micromatrizz[2][40] = 9'b111111111;
assign micromatrizz[2][41] = 9'b111111111;
assign micromatrizz[2][42] = 9'b111111111;
assign micromatrizz[2][43] = 9'b111111111;
assign micromatrizz[2][44] = 9'b111111111;
assign micromatrizz[2][45] = 9'b111111111;
assign micromatrizz[2][46] = 9'b111111111;
assign micromatrizz[2][47] = 9'b111111111;
assign micromatrizz[2][48] = 9'b111111111;
assign micromatrizz[2][49] = 9'b111111111;
assign micromatrizz[2][50] = 9'b111111111;
assign micromatrizz[2][51] = 9'b111111111;
assign micromatrizz[2][52] = 9'b111111111;
assign micromatrizz[2][53] = 9'b111111111;
assign micromatrizz[2][54] = 9'b111111111;
assign micromatrizz[2][55] = 9'b111111111;
assign micromatrizz[2][56] = 9'b111111111;
assign micromatrizz[2][57] = 9'b111111111;
assign micromatrizz[2][58] = 9'b111111111;
assign micromatrizz[2][59] = 9'b111111111;
assign micromatrizz[2][60] = 9'b111111111;
assign micromatrizz[2][61] = 9'b111111111;
assign micromatrizz[2][62] = 9'b111111111;
assign micromatrizz[2][63] = 9'b111111111;
assign micromatrizz[2][64] = 9'b111111111;
assign micromatrizz[2][65] = 9'b111111111;
assign micromatrizz[2][66] = 9'b111111111;
assign micromatrizz[2][67] = 9'b111111111;
assign micromatrizz[2][68] = 9'b111111111;
assign micromatrizz[2][69] = 9'b111111111;
assign micromatrizz[2][70] = 9'b111111111;
assign micromatrizz[2][71] = 9'b111111111;
assign micromatrizz[2][72] = 9'b111111111;
assign micromatrizz[2][73] = 9'b111111111;
assign micromatrizz[2][74] = 9'b111111111;
assign micromatrizz[2][75] = 9'b111111111;
assign micromatrizz[2][76] = 9'b111111111;
assign micromatrizz[2][77] = 9'b111111111;
assign micromatrizz[2][78] = 9'b111111111;
assign micromatrizz[2][79] = 9'b111111111;
assign micromatrizz[2][80] = 9'b111111111;
assign micromatrizz[2][81] = 9'b111111111;
assign micromatrizz[2][82] = 9'b111111111;
assign micromatrizz[2][83] = 9'b111111111;
assign micromatrizz[2][84] = 9'b111111111;
assign micromatrizz[2][85] = 9'b111111111;
assign micromatrizz[2][86] = 9'b111111111;
assign micromatrizz[2][87] = 9'b111111111;
assign micromatrizz[2][88] = 9'b111111111;
assign micromatrizz[2][89] = 9'b111111111;
assign micromatrizz[2][90] = 9'b111111111;
assign micromatrizz[2][91] = 9'b111111111;
assign micromatrizz[2][92] = 9'b111111111;
assign micromatrizz[2][93] = 9'b111111111;
assign micromatrizz[2][94] = 9'b111111111;
assign micromatrizz[2][95] = 9'b111111111;
assign micromatrizz[2][96] = 9'b111111111;
assign micromatrizz[2][97] = 9'b111111111;
assign micromatrizz[2][98] = 9'b111111111;
assign micromatrizz[2][99] = 9'b111111111;
assign micromatrizz[2][100] = 9'b111111111;
assign micromatrizz[2][101] = 9'b111111111;
assign micromatrizz[2][102] = 9'b111111111;
assign micromatrizz[2][103] = 9'b111111111;
assign micromatrizz[2][104] = 9'b111111111;
assign micromatrizz[2][105] = 9'b111111111;
assign micromatrizz[2][106] = 9'b111111111;
assign micromatrizz[2][107] = 9'b111111111;
assign micromatrizz[2][108] = 9'b111111111;
assign micromatrizz[2][109] = 9'b111111111;
assign micromatrizz[2][110] = 9'b111111111;
assign micromatrizz[2][111] = 9'b111111111;
assign micromatrizz[2][112] = 9'b111111111;
assign micromatrizz[2][113] = 9'b111111111;
assign micromatrizz[2][114] = 9'b111111111;
assign micromatrizz[2][115] = 9'b111111111;
assign micromatrizz[2][116] = 9'b111111111;
assign micromatrizz[2][117] = 9'b111111111;
assign micromatrizz[2][118] = 9'b111111111;
assign micromatrizz[2][119] = 9'b111111111;
assign micromatrizz[2][120] = 9'b111111111;
assign micromatrizz[2][121] = 9'b111111111;
assign micromatrizz[2][122] = 9'b111111111;
assign micromatrizz[2][123] = 9'b111111111;
assign micromatrizz[2][124] = 9'b111111111;
assign micromatrizz[2][125] = 9'b111111111;
assign micromatrizz[2][126] = 9'b111111111;
assign micromatrizz[2][127] = 9'b111111111;
assign micromatrizz[2][128] = 9'b111111111;
assign micromatrizz[2][129] = 9'b111111111;
assign micromatrizz[2][130] = 9'b111111111;
assign micromatrizz[2][131] = 9'b111111111;
assign micromatrizz[2][132] = 9'b111111111;
assign micromatrizz[2][133] = 9'b111111111;
assign micromatrizz[2][134] = 9'b111111111;
assign micromatrizz[2][135] = 9'b111111111;
assign micromatrizz[2][136] = 9'b111111111;
assign micromatrizz[2][137] = 9'b111111111;
assign micromatrizz[2][138] = 9'b111111111;
assign micromatrizz[2][139] = 9'b111111111;
assign micromatrizz[2][140] = 9'b111111111;
assign micromatrizz[2][141] = 9'b111111111;
assign micromatrizz[2][142] = 9'b111111111;
assign micromatrizz[2][143] = 9'b111111111;
assign micromatrizz[2][144] = 9'b111111111;
assign micromatrizz[2][145] = 9'b111111111;
assign micromatrizz[2][146] = 9'b111111111;
assign micromatrizz[2][147] = 9'b111111111;
assign micromatrizz[2][148] = 9'b111111111;
assign micromatrizz[2][149] = 9'b111111111;
assign micromatrizz[2][150] = 9'b111111111;
assign micromatrizz[2][151] = 9'b111111111;
assign micromatrizz[2][152] = 9'b111111111;
assign micromatrizz[2][153] = 9'b111111111;
assign micromatrizz[2][154] = 9'b111111111;
assign micromatrizz[2][155] = 9'b111111111;
assign micromatrizz[2][156] = 9'b111111111;
assign micromatrizz[2][157] = 9'b111111111;
assign micromatrizz[2][158] = 9'b111111111;
assign micromatrizz[2][159] = 9'b111111111;
assign micromatrizz[2][160] = 9'b111111111;
assign micromatrizz[2][161] = 9'b111111111;
assign micromatrizz[2][162] = 9'b111111111;
assign micromatrizz[2][163] = 9'b111111111;
assign micromatrizz[2][164] = 9'b111111111;
assign micromatrizz[2][165] = 9'b111111111;
assign micromatrizz[2][166] = 9'b111111111;
assign micromatrizz[2][167] = 9'b111111111;
assign micromatrizz[2][168] = 9'b111111111;
assign micromatrizz[2][169] = 9'b111111111;
assign micromatrizz[2][170] = 9'b111111111;
assign micromatrizz[2][171] = 9'b111111111;
assign micromatrizz[2][172] = 9'b111111111;
assign micromatrizz[2][173] = 9'b111111111;
assign micromatrizz[2][174] = 9'b111111111;
assign micromatrizz[2][175] = 9'b111111111;
assign micromatrizz[2][176] = 9'b111111111;
assign micromatrizz[2][177] = 9'b111111111;
assign micromatrizz[2][178] = 9'b111111111;
assign micromatrizz[2][179] = 9'b111111111;
assign micromatrizz[2][180] = 9'b111111111;
assign micromatrizz[2][181] = 9'b111111111;
assign micromatrizz[2][182] = 9'b111111111;
assign micromatrizz[2][183] = 9'b111111111;
assign micromatrizz[2][184] = 9'b111111111;
assign micromatrizz[2][185] = 9'b111111111;
assign micromatrizz[2][186] = 9'b111111111;
assign micromatrizz[2][187] = 9'b111111111;
assign micromatrizz[2][188] = 9'b111111111;
assign micromatrizz[2][189] = 9'b111111111;
assign micromatrizz[2][190] = 9'b111111111;
assign micromatrizz[2][191] = 9'b111111111;
assign micromatrizz[2][192] = 9'b111111111;
assign micromatrizz[2][193] = 9'b111111111;
assign micromatrizz[2][194] = 9'b111111111;
assign micromatrizz[2][195] = 9'b111111111;
assign micromatrizz[2][196] = 9'b111111111;
assign micromatrizz[2][197] = 9'b111111111;
assign micromatrizz[2][198] = 9'b111111111;
assign micromatrizz[2][199] = 9'b111111111;
assign micromatrizz[2][200] = 9'b111111111;
assign micromatrizz[2][201] = 9'b111111111;
assign micromatrizz[2][202] = 9'b111111111;
assign micromatrizz[2][203] = 9'b111111111;
assign micromatrizz[2][204] = 9'b111111111;
assign micromatrizz[2][205] = 9'b111111111;
assign micromatrizz[2][206] = 9'b111111111;
assign micromatrizz[2][207] = 9'b111111111;
assign micromatrizz[2][208] = 9'b111111111;
assign micromatrizz[2][209] = 9'b111111111;
assign micromatrizz[2][210] = 9'b111111111;
assign micromatrizz[2][211] = 9'b111111111;
assign micromatrizz[2][212] = 9'b111111111;
assign micromatrizz[2][213] = 9'b111111111;
assign micromatrizz[2][214] = 9'b111111111;
assign micromatrizz[2][215] = 9'b111111111;
assign micromatrizz[2][216] = 9'b111111111;
assign micromatrizz[2][217] = 9'b111111111;
assign micromatrizz[2][218] = 9'b111111111;
assign micromatrizz[2][219] = 9'b111111111;
assign micromatrizz[2][220] = 9'b111111111;
assign micromatrizz[2][221] = 9'b111111111;
assign micromatrizz[2][222] = 9'b111111111;
assign micromatrizz[2][223] = 9'b111111111;
assign micromatrizz[2][224] = 9'b111111111;
assign micromatrizz[2][225] = 9'b111111111;
assign micromatrizz[2][226] = 9'b111111111;
assign micromatrizz[2][227] = 9'b111111111;
assign micromatrizz[2][228] = 9'b111111111;
assign micromatrizz[2][229] = 9'b111111111;
assign micromatrizz[2][230] = 9'b111111111;
assign micromatrizz[2][231] = 9'b111111111;
assign micromatrizz[2][232] = 9'b111111111;
assign micromatrizz[2][233] = 9'b111111111;
assign micromatrizz[2][234] = 9'b111111111;
assign micromatrizz[2][235] = 9'b111111111;
assign micromatrizz[2][236] = 9'b111111111;
assign micromatrizz[2][237] = 9'b111111111;
assign micromatrizz[2][238] = 9'b111111111;
assign micromatrizz[2][239] = 9'b111111111;
assign micromatrizz[2][240] = 9'b111111111;
assign micromatrizz[2][241] = 9'b111111111;
assign micromatrizz[2][242] = 9'b111111111;
assign micromatrizz[2][243] = 9'b111111111;
assign micromatrizz[2][244] = 9'b111111111;
assign micromatrizz[2][245] = 9'b111111111;
assign micromatrizz[2][246] = 9'b111111111;
assign micromatrizz[2][247] = 9'b111111111;
assign micromatrizz[2][248] = 9'b111111111;
assign micromatrizz[2][249] = 9'b111111111;
assign micromatrizz[2][250] = 9'b111111111;
assign micromatrizz[2][251] = 9'b111111111;
assign micromatrizz[2][252] = 9'b111111111;
assign micromatrizz[2][253] = 9'b111111111;
assign micromatrizz[2][254] = 9'b111111111;
assign micromatrizz[2][255] = 9'b111111111;
assign micromatrizz[2][256] = 9'b111111111;
assign micromatrizz[2][257] = 9'b111111111;
assign micromatrizz[2][258] = 9'b111111111;
assign micromatrizz[2][259] = 9'b111111111;
assign micromatrizz[2][260] = 9'b111111111;
assign micromatrizz[2][261] = 9'b111111111;
assign micromatrizz[2][262] = 9'b111111111;
assign micromatrizz[2][263] = 9'b111111111;
assign micromatrizz[2][264] = 9'b111111111;
assign micromatrizz[2][265] = 9'b111111111;
assign micromatrizz[2][266] = 9'b111111111;
assign micromatrizz[2][267] = 9'b111111111;
assign micromatrizz[2][268] = 9'b111111111;
assign micromatrizz[2][269] = 9'b111111111;
assign micromatrizz[2][270] = 9'b111111111;
assign micromatrizz[2][271] = 9'b111111111;
assign micromatrizz[2][272] = 9'b111111111;
assign micromatrizz[2][273] = 9'b111111111;
assign micromatrizz[2][274] = 9'b111111111;
assign micromatrizz[2][275] = 9'b111111111;
assign micromatrizz[2][276] = 9'b111111111;
assign micromatrizz[2][277] = 9'b111111111;
assign micromatrizz[2][278] = 9'b111111111;
assign micromatrizz[2][279] = 9'b111111111;
assign micromatrizz[2][280] = 9'b111111111;
assign micromatrizz[2][281] = 9'b111111111;
assign micromatrizz[2][282] = 9'b111111111;
assign micromatrizz[2][283] = 9'b111111111;
assign micromatrizz[2][284] = 9'b111111111;
assign micromatrizz[2][285] = 9'b111111111;
assign micromatrizz[2][286] = 9'b111111111;
assign micromatrizz[2][287] = 9'b111111111;
assign micromatrizz[2][288] = 9'b111111111;
assign micromatrizz[2][289] = 9'b111111111;
assign micromatrizz[2][290] = 9'b111111111;
assign micromatrizz[2][291] = 9'b111111111;
assign micromatrizz[2][292] = 9'b111111111;
assign micromatrizz[2][293] = 9'b111111111;
assign micromatrizz[2][294] = 9'b111111111;
assign micromatrizz[2][295] = 9'b111111111;
assign micromatrizz[2][296] = 9'b111111111;
assign micromatrizz[2][297] = 9'b111111111;
assign micromatrizz[2][298] = 9'b111111111;
assign micromatrizz[2][299] = 9'b111111111;
assign micromatrizz[2][300] = 9'b111111111;
assign micromatrizz[2][301] = 9'b111111111;
assign micromatrizz[2][302] = 9'b111111111;
assign micromatrizz[2][303] = 9'b111111111;
assign micromatrizz[2][304] = 9'b111111111;
assign micromatrizz[2][305] = 9'b111111111;
assign micromatrizz[2][306] = 9'b111111111;
assign micromatrizz[2][307] = 9'b111111111;
assign micromatrizz[2][308] = 9'b111111111;
assign micromatrizz[2][309] = 9'b111111111;
assign micromatrizz[2][310] = 9'b111111111;
assign micromatrizz[2][311] = 9'b111111111;
assign micromatrizz[2][312] = 9'b111111111;
assign micromatrizz[2][313] = 9'b111111111;
assign micromatrizz[2][314] = 9'b111111111;
assign micromatrizz[2][315] = 9'b111111111;
assign micromatrizz[2][316] = 9'b111111111;
assign micromatrizz[2][317] = 9'b111111111;
assign micromatrizz[2][318] = 9'b111111111;
assign micromatrizz[2][319] = 9'b111111111;
assign micromatrizz[2][320] = 9'b111111111;
assign micromatrizz[2][321] = 9'b111111111;
assign micromatrizz[2][322] = 9'b111111111;
assign micromatrizz[2][323] = 9'b111111111;
assign micromatrizz[2][324] = 9'b111111111;
assign micromatrizz[2][325] = 9'b111111111;
assign micromatrizz[2][326] = 9'b111111111;
assign micromatrizz[2][327] = 9'b111111111;
assign micromatrizz[2][328] = 9'b111111111;
assign micromatrizz[2][329] = 9'b111111111;
assign micromatrizz[2][330] = 9'b111111111;
assign micromatrizz[2][331] = 9'b111111111;
assign micromatrizz[2][332] = 9'b111111111;
assign micromatrizz[2][333] = 9'b111111111;
assign micromatrizz[2][334] = 9'b111111111;
assign micromatrizz[2][335] = 9'b111111111;
assign micromatrizz[2][336] = 9'b111111111;
assign micromatrizz[2][337] = 9'b111111111;
assign micromatrizz[2][338] = 9'b111111111;
assign micromatrizz[2][339] = 9'b111111111;
assign micromatrizz[2][340] = 9'b111111111;
assign micromatrizz[2][341] = 9'b111111111;
assign micromatrizz[2][342] = 9'b111111111;
assign micromatrizz[2][343] = 9'b111111111;
assign micromatrizz[2][344] = 9'b111111111;
assign micromatrizz[2][345] = 9'b111111111;
assign micromatrizz[2][346] = 9'b111111111;
assign micromatrizz[2][347] = 9'b111111111;
assign micromatrizz[2][348] = 9'b111111111;
assign micromatrizz[2][349] = 9'b111111111;
assign micromatrizz[2][350] = 9'b111111111;
assign micromatrizz[2][351] = 9'b111111111;
assign micromatrizz[2][352] = 9'b111111111;
assign micromatrizz[2][353] = 9'b111111111;
assign micromatrizz[2][354] = 9'b111111111;
assign micromatrizz[2][355] = 9'b111111111;
assign micromatrizz[2][356] = 9'b111111111;
assign micromatrizz[2][357] = 9'b111111111;
assign micromatrizz[2][358] = 9'b111111111;
assign micromatrizz[2][359] = 9'b111111111;
assign micromatrizz[2][360] = 9'b111111111;
assign micromatrizz[2][361] = 9'b111111111;
assign micromatrizz[2][362] = 9'b111111111;
assign micromatrizz[2][363] = 9'b111111111;
assign micromatrizz[2][364] = 9'b111111111;
assign micromatrizz[2][365] = 9'b111111111;
assign micromatrizz[2][366] = 9'b111111111;
assign micromatrizz[2][367] = 9'b111111111;
assign micromatrizz[2][368] = 9'b111111111;
assign micromatrizz[2][369] = 9'b111111111;
assign micromatrizz[2][370] = 9'b111111111;
assign micromatrizz[2][371] = 9'b111111111;
assign micromatrizz[2][372] = 9'b111111111;
assign micromatrizz[2][373] = 9'b111111111;
assign micromatrizz[2][374] = 9'b111111111;
assign micromatrizz[2][375] = 9'b111111111;
assign micromatrizz[2][376] = 9'b111111111;
assign micromatrizz[2][377] = 9'b111111111;
assign micromatrizz[2][378] = 9'b111111111;
assign micromatrizz[2][379] = 9'b111111111;
assign micromatrizz[2][380] = 9'b111111111;
assign micromatrizz[2][381] = 9'b111111111;
assign micromatrizz[2][382] = 9'b111111111;
assign micromatrizz[2][383] = 9'b111111111;
assign micromatrizz[2][384] = 9'b111111111;
assign micromatrizz[2][385] = 9'b111111111;
assign micromatrizz[2][386] = 9'b111111111;
assign micromatrizz[2][387] = 9'b111111111;
assign micromatrizz[2][388] = 9'b111111111;
assign micromatrizz[2][389] = 9'b111111111;
assign micromatrizz[2][390] = 9'b111111111;
assign micromatrizz[2][391] = 9'b111111111;
assign micromatrizz[2][392] = 9'b111111111;
assign micromatrizz[2][393] = 9'b111111111;
assign micromatrizz[2][394] = 9'b111111111;
assign micromatrizz[2][395] = 9'b111111111;
assign micromatrizz[2][396] = 9'b111111111;
assign micromatrizz[2][397] = 9'b111111111;
assign micromatrizz[2][398] = 9'b111111111;
assign micromatrizz[2][399] = 9'b111111111;
assign micromatrizz[2][400] = 9'b111111111;
assign micromatrizz[2][401] = 9'b111111111;
assign micromatrizz[2][402] = 9'b111111111;
assign micromatrizz[2][403] = 9'b111111111;
assign micromatrizz[2][404] = 9'b111111111;
assign micromatrizz[2][405] = 9'b111111111;
assign micromatrizz[2][406] = 9'b111111111;
assign micromatrizz[2][407] = 9'b111111111;
assign micromatrizz[2][408] = 9'b111111111;
assign micromatrizz[2][409] = 9'b111111111;
assign micromatrizz[2][410] = 9'b111111111;
assign micromatrizz[2][411] = 9'b111111111;
assign micromatrizz[2][412] = 9'b111111111;
assign micromatrizz[2][413] = 9'b111111111;
assign micromatrizz[2][414] = 9'b111111111;
assign micromatrizz[2][415] = 9'b111111111;
assign micromatrizz[2][416] = 9'b111111111;
assign micromatrizz[2][417] = 9'b111111111;
assign micromatrizz[2][418] = 9'b111111111;
assign micromatrizz[2][419] = 9'b111111111;
assign micromatrizz[2][420] = 9'b111111111;
assign micromatrizz[2][421] = 9'b111111111;
assign micromatrizz[2][422] = 9'b111111111;
assign micromatrizz[2][423] = 9'b111111111;
assign micromatrizz[2][424] = 9'b111111111;
assign micromatrizz[2][425] = 9'b111111111;
assign micromatrizz[2][426] = 9'b111111111;
assign micromatrizz[2][427] = 9'b111111111;
assign micromatrizz[2][428] = 9'b111111111;
assign micromatrizz[2][429] = 9'b111111111;
assign micromatrizz[2][430] = 9'b111111111;
assign micromatrizz[2][431] = 9'b111111111;
assign micromatrizz[2][432] = 9'b111111111;
assign micromatrizz[2][433] = 9'b111111111;
assign micromatrizz[2][434] = 9'b111111111;
assign micromatrizz[2][435] = 9'b111111111;
assign micromatrizz[2][436] = 9'b111111111;
assign micromatrizz[2][437] = 9'b111111111;
assign micromatrizz[2][438] = 9'b111111111;
assign micromatrizz[2][439] = 9'b111111111;
assign micromatrizz[2][440] = 9'b111111111;
assign micromatrizz[2][441] = 9'b111111111;
assign micromatrizz[2][442] = 9'b111111111;
assign micromatrizz[2][443] = 9'b111111111;
assign micromatrizz[2][444] = 9'b111111111;
assign micromatrizz[2][445] = 9'b111111111;
assign micromatrizz[2][446] = 9'b111111111;
assign micromatrizz[2][447] = 9'b111111111;
assign micromatrizz[2][448] = 9'b111111111;
assign micromatrizz[2][449] = 9'b111111111;
assign micromatrizz[2][450] = 9'b111111111;
assign micromatrizz[2][451] = 9'b111111111;
assign micromatrizz[2][452] = 9'b111111111;
assign micromatrizz[2][453] = 9'b111111111;
assign micromatrizz[2][454] = 9'b111111111;
assign micromatrizz[2][455] = 9'b111111111;
assign micromatrizz[2][456] = 9'b111111111;
assign micromatrizz[2][457] = 9'b111111111;
assign micromatrizz[2][458] = 9'b111111111;
assign micromatrizz[2][459] = 9'b111111111;
assign micromatrizz[2][460] = 9'b111111111;
assign micromatrizz[2][461] = 9'b111111111;
assign micromatrizz[2][462] = 9'b111111111;
assign micromatrizz[2][463] = 9'b111111111;
assign micromatrizz[2][464] = 9'b111111111;
assign micromatrizz[2][465] = 9'b111111111;
assign micromatrizz[2][466] = 9'b111111111;
assign micromatrizz[2][467] = 9'b111111111;
assign micromatrizz[2][468] = 9'b111111111;
assign micromatrizz[2][469] = 9'b111111111;
assign micromatrizz[2][470] = 9'b111111111;
assign micromatrizz[2][471] = 9'b111111111;
assign micromatrizz[2][472] = 9'b111111111;
assign micromatrizz[2][473] = 9'b111111111;
assign micromatrizz[2][474] = 9'b111111111;
assign micromatrizz[2][475] = 9'b111111111;
assign micromatrizz[2][476] = 9'b111111111;
assign micromatrizz[2][477] = 9'b111111111;
assign micromatrizz[2][478] = 9'b111111111;
assign micromatrizz[2][479] = 9'b111111111;
assign micromatrizz[2][480] = 9'b111111111;
assign micromatrizz[2][481] = 9'b111111111;
assign micromatrizz[2][482] = 9'b111111111;
assign micromatrizz[2][483] = 9'b111111111;
assign micromatrizz[2][484] = 9'b111111111;
assign micromatrizz[2][485] = 9'b111111111;
assign micromatrizz[2][486] = 9'b111111111;
assign micromatrizz[2][487] = 9'b111111111;
assign micromatrizz[2][488] = 9'b111111111;
assign micromatrizz[2][489] = 9'b111111111;
assign micromatrizz[2][490] = 9'b111111111;
assign micromatrizz[2][491] = 9'b111111111;
assign micromatrizz[2][492] = 9'b111111111;
assign micromatrizz[2][493] = 9'b111111111;
assign micromatrizz[2][494] = 9'b111111111;
assign micromatrizz[2][495] = 9'b111111111;
assign micromatrizz[2][496] = 9'b111111111;
assign micromatrizz[2][497] = 9'b111111111;
assign micromatrizz[2][498] = 9'b111111111;
assign micromatrizz[2][499] = 9'b111111111;
assign micromatrizz[2][500] = 9'b111111111;
assign micromatrizz[2][501] = 9'b111111111;
assign micromatrizz[2][502] = 9'b111111111;
assign micromatrizz[2][503] = 9'b111111111;
assign micromatrizz[2][504] = 9'b111111111;
assign micromatrizz[2][505] = 9'b111111111;
assign micromatrizz[2][506] = 9'b111111111;
assign micromatrizz[2][507] = 9'b111111111;
assign micromatrizz[2][508] = 9'b111111111;
assign micromatrizz[2][509] = 9'b111111111;
assign micromatrizz[2][510] = 9'b111111111;
assign micromatrizz[2][511] = 9'b111111111;
assign micromatrizz[2][512] = 9'b111111111;
assign micromatrizz[2][513] = 9'b111111111;
assign micromatrizz[2][514] = 9'b111111111;
assign micromatrizz[2][515] = 9'b111111111;
assign micromatrizz[2][516] = 9'b111111111;
assign micromatrizz[2][517] = 9'b111111111;
assign micromatrizz[2][518] = 9'b111111111;
assign micromatrizz[2][519] = 9'b111111111;
assign micromatrizz[2][520] = 9'b111111111;
assign micromatrizz[2][521] = 9'b111111111;
assign micromatrizz[2][522] = 9'b111111111;
assign micromatrizz[2][523] = 9'b111111111;
assign micromatrizz[2][524] = 9'b111111111;
assign micromatrizz[2][525] = 9'b111111111;
assign micromatrizz[2][526] = 9'b111111111;
assign micromatrizz[2][527] = 9'b111111111;
assign micromatrizz[2][528] = 9'b111111111;
assign micromatrizz[2][529] = 9'b111111111;
assign micromatrizz[2][530] = 9'b111111111;
assign micromatrizz[2][531] = 9'b111111111;
assign micromatrizz[2][532] = 9'b111111111;
assign micromatrizz[2][533] = 9'b111111111;
assign micromatrizz[2][534] = 9'b111111111;
assign micromatrizz[2][535] = 9'b111111111;
assign micromatrizz[2][536] = 9'b111111111;
assign micromatrizz[2][537] = 9'b111111111;
assign micromatrizz[2][538] = 9'b111111111;
assign micromatrizz[2][539] = 9'b111111111;
assign micromatrizz[2][540] = 9'b111111111;
assign micromatrizz[2][541] = 9'b111111111;
assign micromatrizz[2][542] = 9'b111111111;
assign micromatrizz[2][543] = 9'b111111111;
assign micromatrizz[2][544] = 9'b111111111;
assign micromatrizz[2][545] = 9'b111111111;
assign micromatrizz[2][546] = 9'b111111111;
assign micromatrizz[2][547] = 9'b111111111;
assign micromatrizz[2][548] = 9'b111111111;
assign micromatrizz[2][549] = 9'b111111111;
assign micromatrizz[2][550] = 9'b111111111;
assign micromatrizz[2][551] = 9'b111111111;
assign micromatrizz[2][552] = 9'b111111111;
assign micromatrizz[2][553] = 9'b111111111;
assign micromatrizz[2][554] = 9'b111111111;
assign micromatrizz[2][555] = 9'b111111111;
assign micromatrizz[2][556] = 9'b111111111;
assign micromatrizz[2][557] = 9'b111111111;
assign micromatrizz[2][558] = 9'b111111111;
assign micromatrizz[2][559] = 9'b111111111;
assign micromatrizz[2][560] = 9'b111111111;
assign micromatrizz[2][561] = 9'b111111111;
assign micromatrizz[2][562] = 9'b111111111;
assign micromatrizz[2][563] = 9'b111111111;
assign micromatrizz[2][564] = 9'b111111111;
assign micromatrizz[2][565] = 9'b111111111;
assign micromatrizz[2][566] = 9'b111111111;
assign micromatrizz[2][567] = 9'b111111111;
assign micromatrizz[2][568] = 9'b111111111;
assign micromatrizz[2][569] = 9'b111111111;
assign micromatrizz[2][570] = 9'b111111111;
assign micromatrizz[2][571] = 9'b111111111;
assign micromatrizz[2][572] = 9'b111111111;
assign micromatrizz[2][573] = 9'b111111111;
assign micromatrizz[2][574] = 9'b111111111;
assign micromatrizz[2][575] = 9'b111111111;
assign micromatrizz[2][576] = 9'b111111111;
assign micromatrizz[2][577] = 9'b111111111;
assign micromatrizz[2][578] = 9'b111111111;
assign micromatrizz[2][579] = 9'b111111111;
assign micromatrizz[2][580] = 9'b111111111;
assign micromatrizz[2][581] = 9'b111111111;
assign micromatrizz[2][582] = 9'b111111111;
assign micromatrizz[2][583] = 9'b111111111;
assign micromatrizz[2][584] = 9'b111111111;
assign micromatrizz[2][585] = 9'b111111111;
assign micromatrizz[2][586] = 9'b111111111;
assign micromatrizz[2][587] = 9'b111111111;
assign micromatrizz[2][588] = 9'b111111111;
assign micromatrizz[2][589] = 9'b111111111;
assign micromatrizz[2][590] = 9'b111111111;
assign micromatrizz[2][591] = 9'b111111111;
assign micromatrizz[2][592] = 9'b111111111;
assign micromatrizz[2][593] = 9'b111111111;
assign micromatrizz[2][594] = 9'b111111111;
assign micromatrizz[2][595] = 9'b111111111;
assign micromatrizz[2][596] = 9'b111111111;
assign micromatrizz[2][597] = 9'b111111111;
assign micromatrizz[2][598] = 9'b111111111;
assign micromatrizz[2][599] = 9'b111111111;
assign micromatrizz[2][600] = 9'b111111111;
assign micromatrizz[2][601] = 9'b111111111;
assign micromatrizz[2][602] = 9'b111111111;
assign micromatrizz[2][603] = 9'b111111111;
assign micromatrizz[2][604] = 9'b111111111;
assign micromatrizz[2][605] = 9'b111111111;
assign micromatrizz[2][606] = 9'b111111111;
assign micromatrizz[2][607] = 9'b111111111;
assign micromatrizz[2][608] = 9'b111111111;
assign micromatrizz[2][609] = 9'b111111111;
assign micromatrizz[2][610] = 9'b111111111;
assign micromatrizz[2][611] = 9'b111111111;
assign micromatrizz[2][612] = 9'b111111111;
assign micromatrizz[2][613] = 9'b111111111;
assign micromatrizz[2][614] = 9'b111111111;
assign micromatrizz[2][615] = 9'b111111111;
assign micromatrizz[2][616] = 9'b111111111;
assign micromatrizz[2][617] = 9'b111111111;
assign micromatrizz[2][618] = 9'b111111111;
assign micromatrizz[2][619] = 9'b111111111;
assign micromatrizz[2][620] = 9'b111111111;
assign micromatrizz[2][621] = 9'b111111111;
assign micromatrizz[2][622] = 9'b111111111;
assign micromatrizz[2][623] = 9'b111111111;
assign micromatrizz[2][624] = 9'b111111111;
assign micromatrizz[2][625] = 9'b111111111;
assign micromatrizz[2][626] = 9'b111111111;
assign micromatrizz[2][627] = 9'b111111111;
assign micromatrizz[2][628] = 9'b111111111;
assign micromatrizz[2][629] = 9'b111111111;
assign micromatrizz[2][630] = 9'b111111111;
assign micromatrizz[2][631] = 9'b111111111;
assign micromatrizz[2][632] = 9'b111111111;
assign micromatrizz[2][633] = 9'b111111111;
assign micromatrizz[2][634] = 9'b111111111;
assign micromatrizz[2][635] = 9'b111111111;
assign micromatrizz[2][636] = 9'b111111111;
assign micromatrizz[2][637] = 9'b111111111;
assign micromatrizz[2][638] = 9'b111111111;
assign micromatrizz[2][639] = 9'b111111111;
assign micromatrizz[3][0] = 9'b111111111;
assign micromatrizz[3][1] = 9'b111111111;
assign micromatrizz[3][2] = 9'b111111111;
assign micromatrizz[3][3] = 9'b111111111;
assign micromatrizz[3][4] = 9'b111111111;
assign micromatrizz[3][5] = 9'b111111111;
assign micromatrizz[3][6] = 9'b111111111;
assign micromatrizz[3][7] = 9'b111111111;
assign micromatrizz[3][8] = 9'b111111111;
assign micromatrizz[3][9] = 9'b111111111;
assign micromatrizz[3][10] = 9'b111111111;
assign micromatrizz[3][11] = 9'b111111111;
assign micromatrizz[3][12] = 9'b111111111;
assign micromatrizz[3][13] = 9'b111111111;
assign micromatrizz[3][14] = 9'b111111111;
assign micromatrizz[3][15] = 9'b111111111;
assign micromatrizz[3][16] = 9'b111111111;
assign micromatrizz[3][17] = 9'b111111111;
assign micromatrizz[3][18] = 9'b111111111;
assign micromatrizz[3][19] = 9'b111111111;
assign micromatrizz[3][20] = 9'b111111111;
assign micromatrizz[3][21] = 9'b111111111;
assign micromatrizz[3][22] = 9'b111111111;
assign micromatrizz[3][23] = 9'b111111111;
assign micromatrizz[3][24] = 9'b111111111;
assign micromatrizz[3][25] = 9'b111111111;
assign micromatrizz[3][26] = 9'b111111111;
assign micromatrizz[3][27] = 9'b111111111;
assign micromatrizz[3][28] = 9'b111111111;
assign micromatrizz[3][29] = 9'b111111111;
assign micromatrizz[3][30] = 9'b111111111;
assign micromatrizz[3][31] = 9'b111111111;
assign micromatrizz[3][32] = 9'b111111111;
assign micromatrizz[3][33] = 9'b111111111;
assign micromatrizz[3][34] = 9'b111111111;
assign micromatrizz[3][35] = 9'b111111111;
assign micromatrizz[3][36] = 9'b111111111;
assign micromatrizz[3][37] = 9'b111111111;
assign micromatrizz[3][38] = 9'b111111111;
assign micromatrizz[3][39] = 9'b111111111;
assign micromatrizz[3][40] = 9'b111111111;
assign micromatrizz[3][41] = 9'b111111111;
assign micromatrizz[3][42] = 9'b111111111;
assign micromatrizz[3][43] = 9'b111111111;
assign micromatrizz[3][44] = 9'b111111111;
assign micromatrizz[3][45] = 9'b111111111;
assign micromatrizz[3][46] = 9'b111111111;
assign micromatrizz[3][47] = 9'b111111111;
assign micromatrizz[3][48] = 9'b111111111;
assign micromatrizz[3][49] = 9'b111111111;
assign micromatrizz[3][50] = 9'b111111111;
assign micromatrizz[3][51] = 9'b111111111;
assign micromatrizz[3][52] = 9'b111111111;
assign micromatrizz[3][53] = 9'b111111111;
assign micromatrizz[3][54] = 9'b111111111;
assign micromatrizz[3][55] = 9'b111111111;
assign micromatrizz[3][56] = 9'b111111111;
assign micromatrizz[3][57] = 9'b111111111;
assign micromatrizz[3][58] = 9'b111111111;
assign micromatrizz[3][59] = 9'b111111111;
assign micromatrizz[3][60] = 9'b111111111;
assign micromatrizz[3][61] = 9'b111111111;
assign micromatrizz[3][62] = 9'b111111111;
assign micromatrizz[3][63] = 9'b111111111;
assign micromatrizz[3][64] = 9'b111111111;
assign micromatrizz[3][65] = 9'b111111111;
assign micromatrizz[3][66] = 9'b111111111;
assign micromatrizz[3][67] = 9'b111111111;
assign micromatrizz[3][68] = 9'b111111111;
assign micromatrizz[3][69] = 9'b111111111;
assign micromatrizz[3][70] = 9'b111111111;
assign micromatrizz[3][71] = 9'b111111111;
assign micromatrizz[3][72] = 9'b111111111;
assign micromatrizz[3][73] = 9'b111111111;
assign micromatrizz[3][74] = 9'b111111111;
assign micromatrizz[3][75] = 9'b111111111;
assign micromatrizz[3][76] = 9'b111111111;
assign micromatrizz[3][77] = 9'b111111111;
assign micromatrizz[3][78] = 9'b111111111;
assign micromatrizz[3][79] = 9'b111111111;
assign micromatrizz[3][80] = 9'b111111111;
assign micromatrizz[3][81] = 9'b111111111;
assign micromatrizz[3][82] = 9'b111111111;
assign micromatrizz[3][83] = 9'b111111111;
assign micromatrizz[3][84] = 9'b111111111;
assign micromatrizz[3][85] = 9'b111111111;
assign micromatrizz[3][86] = 9'b111111111;
assign micromatrizz[3][87] = 9'b111111111;
assign micromatrizz[3][88] = 9'b111111111;
assign micromatrizz[3][89] = 9'b111111111;
assign micromatrizz[3][90] = 9'b111111111;
assign micromatrizz[3][91] = 9'b111111111;
assign micromatrizz[3][92] = 9'b111111111;
assign micromatrizz[3][93] = 9'b111111111;
assign micromatrizz[3][94] = 9'b111111111;
assign micromatrizz[3][95] = 9'b111111111;
assign micromatrizz[3][96] = 9'b111111111;
assign micromatrizz[3][97] = 9'b111111111;
assign micromatrizz[3][98] = 9'b111111111;
assign micromatrizz[3][99] = 9'b111111111;
assign micromatrizz[3][100] = 9'b111111111;
assign micromatrizz[3][101] = 9'b111111111;
assign micromatrizz[3][102] = 9'b111111111;
assign micromatrizz[3][103] = 9'b111111111;
assign micromatrizz[3][104] = 9'b111111111;
assign micromatrizz[3][105] = 9'b111111111;
assign micromatrizz[3][106] = 9'b111111111;
assign micromatrizz[3][107] = 9'b111111111;
assign micromatrizz[3][108] = 9'b111111111;
assign micromatrizz[3][109] = 9'b111111111;
assign micromatrizz[3][110] = 9'b111111111;
assign micromatrizz[3][111] = 9'b111111111;
assign micromatrizz[3][112] = 9'b111111111;
assign micromatrizz[3][113] = 9'b111111111;
assign micromatrizz[3][114] = 9'b111111111;
assign micromatrizz[3][115] = 9'b111111111;
assign micromatrizz[3][116] = 9'b111111111;
assign micromatrizz[3][117] = 9'b111111111;
assign micromatrizz[3][118] = 9'b111111111;
assign micromatrizz[3][119] = 9'b111111111;
assign micromatrizz[3][120] = 9'b111111111;
assign micromatrizz[3][121] = 9'b111111111;
assign micromatrizz[3][122] = 9'b111111111;
assign micromatrizz[3][123] = 9'b111111111;
assign micromatrizz[3][124] = 9'b111111111;
assign micromatrizz[3][125] = 9'b111111111;
assign micromatrizz[3][126] = 9'b111111111;
assign micromatrizz[3][127] = 9'b111111111;
assign micromatrizz[3][128] = 9'b111111111;
assign micromatrizz[3][129] = 9'b111111111;
assign micromatrizz[3][130] = 9'b111111111;
assign micromatrizz[3][131] = 9'b111111111;
assign micromatrizz[3][132] = 9'b111111111;
assign micromatrizz[3][133] = 9'b111111111;
assign micromatrizz[3][134] = 9'b111111111;
assign micromatrizz[3][135] = 9'b111111111;
assign micromatrizz[3][136] = 9'b111111111;
assign micromatrizz[3][137] = 9'b111111111;
assign micromatrizz[3][138] = 9'b111111111;
assign micromatrizz[3][139] = 9'b111111111;
assign micromatrizz[3][140] = 9'b111111111;
assign micromatrizz[3][141] = 9'b111111111;
assign micromatrizz[3][142] = 9'b111111111;
assign micromatrizz[3][143] = 9'b111111111;
assign micromatrizz[3][144] = 9'b111111111;
assign micromatrizz[3][145] = 9'b111111111;
assign micromatrizz[3][146] = 9'b111111111;
assign micromatrizz[3][147] = 9'b111111111;
assign micromatrizz[3][148] = 9'b111111111;
assign micromatrizz[3][149] = 9'b111111111;
assign micromatrizz[3][150] = 9'b111111111;
assign micromatrizz[3][151] = 9'b111111111;
assign micromatrizz[3][152] = 9'b111111111;
assign micromatrizz[3][153] = 9'b111111111;
assign micromatrizz[3][154] = 9'b111111111;
assign micromatrizz[3][155] = 9'b111111111;
assign micromatrizz[3][156] = 9'b111111111;
assign micromatrizz[3][157] = 9'b111111111;
assign micromatrizz[3][158] = 9'b111111111;
assign micromatrizz[3][159] = 9'b111111111;
assign micromatrizz[3][160] = 9'b111111111;
assign micromatrizz[3][161] = 9'b111111111;
assign micromatrizz[3][162] = 9'b111111111;
assign micromatrizz[3][163] = 9'b111111111;
assign micromatrizz[3][164] = 9'b111111111;
assign micromatrizz[3][165] = 9'b111111111;
assign micromatrizz[3][166] = 9'b111111111;
assign micromatrizz[3][167] = 9'b111111111;
assign micromatrizz[3][168] = 9'b111111111;
assign micromatrizz[3][169] = 9'b111111111;
assign micromatrizz[3][170] = 9'b111111111;
assign micromatrizz[3][171] = 9'b111111111;
assign micromatrizz[3][172] = 9'b111111111;
assign micromatrizz[3][173] = 9'b111111111;
assign micromatrizz[3][174] = 9'b111111111;
assign micromatrizz[3][175] = 9'b111111111;
assign micromatrizz[3][176] = 9'b111111111;
assign micromatrizz[3][177] = 9'b111111111;
assign micromatrizz[3][178] = 9'b111111111;
assign micromatrizz[3][179] = 9'b111111111;
assign micromatrizz[3][180] = 9'b111111111;
assign micromatrizz[3][181] = 9'b111111111;
assign micromatrizz[3][182] = 9'b111111111;
assign micromatrizz[3][183] = 9'b111111111;
assign micromatrizz[3][184] = 9'b111111111;
assign micromatrizz[3][185] = 9'b111111111;
assign micromatrizz[3][186] = 9'b111111111;
assign micromatrizz[3][187] = 9'b111111111;
assign micromatrizz[3][188] = 9'b111111111;
assign micromatrizz[3][189] = 9'b111111111;
assign micromatrizz[3][190] = 9'b111111111;
assign micromatrizz[3][191] = 9'b111111111;
assign micromatrizz[3][192] = 9'b111111111;
assign micromatrizz[3][193] = 9'b111111111;
assign micromatrizz[3][194] = 9'b111111111;
assign micromatrizz[3][195] = 9'b111111111;
assign micromatrizz[3][196] = 9'b111111111;
assign micromatrizz[3][197] = 9'b111111111;
assign micromatrizz[3][198] = 9'b111111111;
assign micromatrizz[3][199] = 9'b111111111;
assign micromatrizz[3][200] = 9'b111111111;
assign micromatrizz[3][201] = 9'b111111111;
assign micromatrizz[3][202] = 9'b111111111;
assign micromatrizz[3][203] = 9'b111111111;
assign micromatrizz[3][204] = 9'b111111111;
assign micromatrizz[3][205] = 9'b111111111;
assign micromatrizz[3][206] = 9'b111111111;
assign micromatrizz[3][207] = 9'b111111111;
assign micromatrizz[3][208] = 9'b111111111;
assign micromatrizz[3][209] = 9'b111111111;
assign micromatrizz[3][210] = 9'b111111111;
assign micromatrizz[3][211] = 9'b111111111;
assign micromatrizz[3][212] = 9'b111111111;
assign micromatrizz[3][213] = 9'b111111111;
assign micromatrizz[3][214] = 9'b111111111;
assign micromatrizz[3][215] = 9'b111111111;
assign micromatrizz[3][216] = 9'b111111111;
assign micromatrizz[3][217] = 9'b111111111;
assign micromatrizz[3][218] = 9'b111111111;
assign micromatrizz[3][219] = 9'b111111111;
assign micromatrizz[3][220] = 9'b111111111;
assign micromatrizz[3][221] = 9'b111111111;
assign micromatrizz[3][222] = 9'b111111111;
assign micromatrizz[3][223] = 9'b111111111;
assign micromatrizz[3][224] = 9'b111111111;
assign micromatrizz[3][225] = 9'b111111111;
assign micromatrizz[3][226] = 9'b111111111;
assign micromatrizz[3][227] = 9'b111111111;
assign micromatrizz[3][228] = 9'b111111111;
assign micromatrizz[3][229] = 9'b111111111;
assign micromatrizz[3][230] = 9'b111111111;
assign micromatrizz[3][231] = 9'b111111111;
assign micromatrizz[3][232] = 9'b111111111;
assign micromatrizz[3][233] = 9'b111111111;
assign micromatrizz[3][234] = 9'b111111111;
assign micromatrizz[3][235] = 9'b111111111;
assign micromatrizz[3][236] = 9'b111111111;
assign micromatrizz[3][237] = 9'b111111111;
assign micromatrizz[3][238] = 9'b111111111;
assign micromatrizz[3][239] = 9'b111111111;
assign micromatrizz[3][240] = 9'b111111111;
assign micromatrizz[3][241] = 9'b111111111;
assign micromatrizz[3][242] = 9'b111111111;
assign micromatrizz[3][243] = 9'b111111111;
assign micromatrizz[3][244] = 9'b111111111;
assign micromatrizz[3][245] = 9'b111111111;
assign micromatrizz[3][246] = 9'b111111111;
assign micromatrizz[3][247] = 9'b111111111;
assign micromatrizz[3][248] = 9'b111111111;
assign micromatrizz[3][249] = 9'b111111111;
assign micromatrizz[3][250] = 9'b111111111;
assign micromatrizz[3][251] = 9'b111111111;
assign micromatrizz[3][252] = 9'b111111111;
assign micromatrizz[3][253] = 9'b111111111;
assign micromatrizz[3][254] = 9'b111111111;
assign micromatrizz[3][255] = 9'b111111111;
assign micromatrizz[3][256] = 9'b111111111;
assign micromatrizz[3][257] = 9'b111111111;
assign micromatrizz[3][258] = 9'b111111111;
assign micromatrizz[3][259] = 9'b111111111;
assign micromatrizz[3][260] = 9'b111111111;
assign micromatrizz[3][261] = 9'b111111111;
assign micromatrizz[3][262] = 9'b111111111;
assign micromatrizz[3][263] = 9'b111111111;
assign micromatrizz[3][264] = 9'b111111111;
assign micromatrizz[3][265] = 9'b111111111;
assign micromatrizz[3][266] = 9'b111111111;
assign micromatrizz[3][267] = 9'b111111111;
assign micromatrizz[3][268] = 9'b111111111;
assign micromatrizz[3][269] = 9'b111111111;
assign micromatrizz[3][270] = 9'b111111111;
assign micromatrizz[3][271] = 9'b111111111;
assign micromatrizz[3][272] = 9'b111111111;
assign micromatrizz[3][273] = 9'b111111111;
assign micromatrizz[3][274] = 9'b111111111;
assign micromatrizz[3][275] = 9'b111111111;
assign micromatrizz[3][276] = 9'b111111111;
assign micromatrizz[3][277] = 9'b111111111;
assign micromatrizz[3][278] = 9'b111111111;
assign micromatrizz[3][279] = 9'b111111111;
assign micromatrizz[3][280] = 9'b111111111;
assign micromatrizz[3][281] = 9'b111111111;
assign micromatrizz[3][282] = 9'b111111111;
assign micromatrizz[3][283] = 9'b111111111;
assign micromatrizz[3][284] = 9'b111111111;
assign micromatrizz[3][285] = 9'b111111111;
assign micromatrizz[3][286] = 9'b111111111;
assign micromatrizz[3][287] = 9'b111111111;
assign micromatrizz[3][288] = 9'b111111111;
assign micromatrizz[3][289] = 9'b111111111;
assign micromatrizz[3][290] = 9'b111111111;
assign micromatrizz[3][291] = 9'b111111111;
assign micromatrizz[3][292] = 9'b111111111;
assign micromatrizz[3][293] = 9'b111111111;
assign micromatrizz[3][294] = 9'b111111111;
assign micromatrizz[3][295] = 9'b111111111;
assign micromatrizz[3][296] = 9'b111111111;
assign micromatrizz[3][297] = 9'b111111111;
assign micromatrizz[3][298] = 9'b111111111;
assign micromatrizz[3][299] = 9'b111111111;
assign micromatrizz[3][300] = 9'b111111111;
assign micromatrizz[3][301] = 9'b111111111;
assign micromatrizz[3][302] = 9'b111111111;
assign micromatrizz[3][303] = 9'b111111111;
assign micromatrizz[3][304] = 9'b111111111;
assign micromatrizz[3][305] = 9'b111111111;
assign micromatrizz[3][306] = 9'b111111111;
assign micromatrizz[3][307] = 9'b111111111;
assign micromatrizz[3][308] = 9'b111111111;
assign micromatrizz[3][309] = 9'b111111111;
assign micromatrizz[3][310] = 9'b111111111;
assign micromatrizz[3][311] = 9'b111111111;
assign micromatrizz[3][312] = 9'b111111111;
assign micromatrizz[3][313] = 9'b111111111;
assign micromatrizz[3][314] = 9'b111111111;
assign micromatrizz[3][315] = 9'b111111111;
assign micromatrizz[3][316] = 9'b111111111;
assign micromatrizz[3][317] = 9'b111111111;
assign micromatrizz[3][318] = 9'b111111111;
assign micromatrizz[3][319] = 9'b111111111;
assign micromatrizz[3][320] = 9'b111111111;
assign micromatrizz[3][321] = 9'b111111111;
assign micromatrizz[3][322] = 9'b111111111;
assign micromatrizz[3][323] = 9'b111111111;
assign micromatrizz[3][324] = 9'b111111111;
assign micromatrizz[3][325] = 9'b111111111;
assign micromatrizz[3][326] = 9'b111111111;
assign micromatrizz[3][327] = 9'b111111111;
assign micromatrizz[3][328] = 9'b111111111;
assign micromatrizz[3][329] = 9'b111111111;
assign micromatrizz[3][330] = 9'b111111111;
assign micromatrizz[3][331] = 9'b111111111;
assign micromatrizz[3][332] = 9'b111111111;
assign micromatrizz[3][333] = 9'b111111111;
assign micromatrizz[3][334] = 9'b111111111;
assign micromatrizz[3][335] = 9'b111111111;
assign micromatrizz[3][336] = 9'b111111111;
assign micromatrizz[3][337] = 9'b111111111;
assign micromatrizz[3][338] = 9'b111111111;
assign micromatrizz[3][339] = 9'b111111111;
assign micromatrizz[3][340] = 9'b111111111;
assign micromatrizz[3][341] = 9'b111111111;
assign micromatrizz[3][342] = 9'b111111111;
assign micromatrizz[3][343] = 9'b111111111;
assign micromatrizz[3][344] = 9'b111111111;
assign micromatrizz[3][345] = 9'b111111111;
assign micromatrizz[3][346] = 9'b111111111;
assign micromatrizz[3][347] = 9'b111111111;
assign micromatrizz[3][348] = 9'b111111111;
assign micromatrizz[3][349] = 9'b111111111;
assign micromatrizz[3][350] = 9'b111111111;
assign micromatrizz[3][351] = 9'b111111111;
assign micromatrizz[3][352] = 9'b111111111;
assign micromatrizz[3][353] = 9'b111111111;
assign micromatrizz[3][354] = 9'b111111111;
assign micromatrizz[3][355] = 9'b111111111;
assign micromatrizz[3][356] = 9'b111111111;
assign micromatrizz[3][357] = 9'b111111111;
assign micromatrizz[3][358] = 9'b111111111;
assign micromatrizz[3][359] = 9'b111111111;
assign micromatrizz[3][360] = 9'b111111111;
assign micromatrizz[3][361] = 9'b111111111;
assign micromatrizz[3][362] = 9'b111111111;
assign micromatrizz[3][363] = 9'b111111111;
assign micromatrizz[3][364] = 9'b111111111;
assign micromatrizz[3][365] = 9'b111111111;
assign micromatrizz[3][366] = 9'b111111111;
assign micromatrizz[3][367] = 9'b111111111;
assign micromatrizz[3][368] = 9'b111111111;
assign micromatrizz[3][369] = 9'b111111111;
assign micromatrizz[3][370] = 9'b111111111;
assign micromatrizz[3][371] = 9'b111111111;
assign micromatrizz[3][372] = 9'b111111111;
assign micromatrizz[3][373] = 9'b111111111;
assign micromatrizz[3][374] = 9'b111111111;
assign micromatrizz[3][375] = 9'b111111111;
assign micromatrizz[3][376] = 9'b111111111;
assign micromatrizz[3][377] = 9'b111111111;
assign micromatrizz[3][378] = 9'b111111111;
assign micromatrizz[3][379] = 9'b111111111;
assign micromatrizz[3][380] = 9'b111111111;
assign micromatrizz[3][381] = 9'b111111111;
assign micromatrizz[3][382] = 9'b111111111;
assign micromatrizz[3][383] = 9'b111111111;
assign micromatrizz[3][384] = 9'b111111111;
assign micromatrizz[3][385] = 9'b111111111;
assign micromatrizz[3][386] = 9'b111111111;
assign micromatrizz[3][387] = 9'b111111111;
assign micromatrizz[3][388] = 9'b111111111;
assign micromatrizz[3][389] = 9'b111111111;
assign micromatrizz[3][390] = 9'b111111111;
assign micromatrizz[3][391] = 9'b111111111;
assign micromatrizz[3][392] = 9'b111111111;
assign micromatrizz[3][393] = 9'b111111111;
assign micromatrizz[3][394] = 9'b111111111;
assign micromatrizz[3][395] = 9'b111111111;
assign micromatrizz[3][396] = 9'b111111111;
assign micromatrizz[3][397] = 9'b111111111;
assign micromatrizz[3][398] = 9'b111111111;
assign micromatrizz[3][399] = 9'b111111111;
assign micromatrizz[3][400] = 9'b111111111;
assign micromatrizz[3][401] = 9'b111111111;
assign micromatrizz[3][402] = 9'b111111111;
assign micromatrizz[3][403] = 9'b111111111;
assign micromatrizz[3][404] = 9'b111111111;
assign micromatrizz[3][405] = 9'b111111111;
assign micromatrizz[3][406] = 9'b111111111;
assign micromatrizz[3][407] = 9'b111111111;
assign micromatrizz[3][408] = 9'b111111111;
assign micromatrizz[3][409] = 9'b111111111;
assign micromatrizz[3][410] = 9'b111111111;
assign micromatrizz[3][411] = 9'b111111111;
assign micromatrizz[3][412] = 9'b111111111;
assign micromatrizz[3][413] = 9'b111111111;
assign micromatrizz[3][414] = 9'b111111111;
assign micromatrizz[3][415] = 9'b111111111;
assign micromatrizz[3][416] = 9'b111111111;
assign micromatrizz[3][417] = 9'b111111111;
assign micromatrizz[3][418] = 9'b111111111;
assign micromatrizz[3][419] = 9'b111111111;
assign micromatrizz[3][420] = 9'b111111111;
assign micromatrizz[3][421] = 9'b111111111;
assign micromatrizz[3][422] = 9'b111111111;
assign micromatrizz[3][423] = 9'b111111111;
assign micromatrizz[3][424] = 9'b111111111;
assign micromatrizz[3][425] = 9'b111111111;
assign micromatrizz[3][426] = 9'b111111111;
assign micromatrizz[3][427] = 9'b111111111;
assign micromatrizz[3][428] = 9'b111111111;
assign micromatrizz[3][429] = 9'b111111111;
assign micromatrizz[3][430] = 9'b111111111;
assign micromatrizz[3][431] = 9'b111111111;
assign micromatrizz[3][432] = 9'b111111111;
assign micromatrizz[3][433] = 9'b111111111;
assign micromatrizz[3][434] = 9'b111111111;
assign micromatrizz[3][435] = 9'b111111111;
assign micromatrizz[3][436] = 9'b111111111;
assign micromatrizz[3][437] = 9'b111111111;
assign micromatrizz[3][438] = 9'b111111111;
assign micromatrizz[3][439] = 9'b111111111;
assign micromatrizz[3][440] = 9'b111111111;
assign micromatrizz[3][441] = 9'b111111111;
assign micromatrizz[3][442] = 9'b111111111;
assign micromatrizz[3][443] = 9'b111111111;
assign micromatrizz[3][444] = 9'b111111111;
assign micromatrizz[3][445] = 9'b111111111;
assign micromatrizz[3][446] = 9'b111111111;
assign micromatrizz[3][447] = 9'b111111111;
assign micromatrizz[3][448] = 9'b111111111;
assign micromatrizz[3][449] = 9'b111111111;
assign micromatrizz[3][450] = 9'b111111111;
assign micromatrizz[3][451] = 9'b111111111;
assign micromatrizz[3][452] = 9'b111111111;
assign micromatrizz[3][453] = 9'b111111111;
assign micromatrizz[3][454] = 9'b111111111;
assign micromatrizz[3][455] = 9'b111111111;
assign micromatrizz[3][456] = 9'b111111111;
assign micromatrizz[3][457] = 9'b111111111;
assign micromatrizz[3][458] = 9'b111111111;
assign micromatrizz[3][459] = 9'b111111111;
assign micromatrizz[3][460] = 9'b111111111;
assign micromatrizz[3][461] = 9'b111111111;
assign micromatrizz[3][462] = 9'b111111111;
assign micromatrizz[3][463] = 9'b111111111;
assign micromatrizz[3][464] = 9'b111111111;
assign micromatrizz[3][465] = 9'b111111111;
assign micromatrizz[3][466] = 9'b111111111;
assign micromatrizz[3][467] = 9'b111111111;
assign micromatrizz[3][468] = 9'b111111111;
assign micromatrizz[3][469] = 9'b111111111;
assign micromatrizz[3][470] = 9'b111111111;
assign micromatrizz[3][471] = 9'b111111111;
assign micromatrizz[3][472] = 9'b111111111;
assign micromatrizz[3][473] = 9'b111111111;
assign micromatrizz[3][474] = 9'b111111111;
assign micromatrizz[3][475] = 9'b111111111;
assign micromatrizz[3][476] = 9'b111111111;
assign micromatrizz[3][477] = 9'b111111111;
assign micromatrizz[3][478] = 9'b111111111;
assign micromatrizz[3][479] = 9'b111111111;
assign micromatrizz[3][480] = 9'b111111111;
assign micromatrizz[3][481] = 9'b111111111;
assign micromatrizz[3][482] = 9'b111111111;
assign micromatrizz[3][483] = 9'b111111111;
assign micromatrizz[3][484] = 9'b111111111;
assign micromatrizz[3][485] = 9'b111111111;
assign micromatrizz[3][486] = 9'b111111111;
assign micromatrizz[3][487] = 9'b111111111;
assign micromatrizz[3][488] = 9'b111111111;
assign micromatrizz[3][489] = 9'b111111111;
assign micromatrizz[3][490] = 9'b111111111;
assign micromatrizz[3][491] = 9'b111111111;
assign micromatrizz[3][492] = 9'b111111111;
assign micromatrizz[3][493] = 9'b111111111;
assign micromatrizz[3][494] = 9'b111111111;
assign micromatrizz[3][495] = 9'b111111111;
assign micromatrizz[3][496] = 9'b111111111;
assign micromatrizz[3][497] = 9'b111111111;
assign micromatrizz[3][498] = 9'b111111111;
assign micromatrizz[3][499] = 9'b111111111;
assign micromatrizz[3][500] = 9'b111111111;
assign micromatrizz[3][501] = 9'b111111111;
assign micromatrizz[3][502] = 9'b111111111;
assign micromatrizz[3][503] = 9'b111111111;
assign micromatrizz[3][504] = 9'b111111111;
assign micromatrizz[3][505] = 9'b111111111;
assign micromatrizz[3][506] = 9'b111111111;
assign micromatrizz[3][507] = 9'b111111111;
assign micromatrizz[3][508] = 9'b111111111;
assign micromatrizz[3][509] = 9'b111111111;
assign micromatrizz[3][510] = 9'b111111111;
assign micromatrizz[3][511] = 9'b111111111;
assign micromatrizz[3][512] = 9'b111111111;
assign micromatrizz[3][513] = 9'b111111111;
assign micromatrizz[3][514] = 9'b111111111;
assign micromatrizz[3][515] = 9'b111111111;
assign micromatrizz[3][516] = 9'b111111111;
assign micromatrizz[3][517] = 9'b111111111;
assign micromatrizz[3][518] = 9'b111111111;
assign micromatrizz[3][519] = 9'b111111111;
assign micromatrizz[3][520] = 9'b111111111;
assign micromatrizz[3][521] = 9'b111111111;
assign micromatrizz[3][522] = 9'b111111111;
assign micromatrizz[3][523] = 9'b111111111;
assign micromatrizz[3][524] = 9'b111111111;
assign micromatrizz[3][525] = 9'b111111111;
assign micromatrizz[3][526] = 9'b111111111;
assign micromatrizz[3][527] = 9'b111111111;
assign micromatrizz[3][528] = 9'b111111111;
assign micromatrizz[3][529] = 9'b111111111;
assign micromatrizz[3][530] = 9'b111111111;
assign micromatrizz[3][531] = 9'b111111111;
assign micromatrizz[3][532] = 9'b111111111;
assign micromatrizz[3][533] = 9'b111111111;
assign micromatrizz[3][534] = 9'b111111111;
assign micromatrizz[3][535] = 9'b111111111;
assign micromatrizz[3][536] = 9'b111111111;
assign micromatrizz[3][537] = 9'b111111111;
assign micromatrizz[3][538] = 9'b111111111;
assign micromatrizz[3][539] = 9'b111111111;
assign micromatrizz[3][540] = 9'b111111111;
assign micromatrizz[3][541] = 9'b111111111;
assign micromatrizz[3][542] = 9'b111111111;
assign micromatrizz[3][543] = 9'b111111111;
assign micromatrizz[3][544] = 9'b111111111;
assign micromatrizz[3][545] = 9'b111111111;
assign micromatrizz[3][546] = 9'b111111111;
assign micromatrizz[3][547] = 9'b111111111;
assign micromatrizz[3][548] = 9'b111111111;
assign micromatrizz[3][549] = 9'b111111111;
assign micromatrizz[3][550] = 9'b111111111;
assign micromatrizz[3][551] = 9'b111111111;
assign micromatrizz[3][552] = 9'b111111111;
assign micromatrizz[3][553] = 9'b111111111;
assign micromatrizz[3][554] = 9'b111111111;
assign micromatrizz[3][555] = 9'b111111111;
assign micromatrizz[3][556] = 9'b111111111;
assign micromatrizz[3][557] = 9'b111111111;
assign micromatrizz[3][558] = 9'b111111111;
assign micromatrizz[3][559] = 9'b111111111;
assign micromatrizz[3][560] = 9'b111111111;
assign micromatrizz[3][561] = 9'b111111111;
assign micromatrizz[3][562] = 9'b111111111;
assign micromatrizz[3][563] = 9'b111111111;
assign micromatrizz[3][564] = 9'b111111111;
assign micromatrizz[3][565] = 9'b111111111;
assign micromatrizz[3][566] = 9'b111111111;
assign micromatrizz[3][567] = 9'b111111111;
assign micromatrizz[3][568] = 9'b111111111;
assign micromatrizz[3][569] = 9'b111111111;
assign micromatrizz[3][570] = 9'b111111111;
assign micromatrizz[3][571] = 9'b111111111;
assign micromatrizz[3][572] = 9'b111111111;
assign micromatrizz[3][573] = 9'b111111111;
assign micromatrizz[3][574] = 9'b111111111;
assign micromatrizz[3][575] = 9'b111111111;
assign micromatrizz[3][576] = 9'b111111111;
assign micromatrizz[3][577] = 9'b111111111;
assign micromatrizz[3][578] = 9'b111111111;
assign micromatrizz[3][579] = 9'b111111111;
assign micromatrizz[3][580] = 9'b111111111;
assign micromatrizz[3][581] = 9'b111111111;
assign micromatrizz[3][582] = 9'b111111111;
assign micromatrizz[3][583] = 9'b111111111;
assign micromatrizz[3][584] = 9'b111111111;
assign micromatrizz[3][585] = 9'b111111111;
assign micromatrizz[3][586] = 9'b111111111;
assign micromatrizz[3][587] = 9'b111111111;
assign micromatrizz[3][588] = 9'b111111111;
assign micromatrizz[3][589] = 9'b111111111;
assign micromatrizz[3][590] = 9'b111111111;
assign micromatrizz[3][591] = 9'b111111111;
assign micromatrizz[3][592] = 9'b111111111;
assign micromatrizz[3][593] = 9'b111111111;
assign micromatrizz[3][594] = 9'b111111111;
assign micromatrizz[3][595] = 9'b111111111;
assign micromatrizz[3][596] = 9'b111111111;
assign micromatrizz[3][597] = 9'b111111111;
assign micromatrizz[3][598] = 9'b111111111;
assign micromatrizz[3][599] = 9'b111111111;
assign micromatrizz[3][600] = 9'b111111111;
assign micromatrizz[3][601] = 9'b111111111;
assign micromatrizz[3][602] = 9'b111111111;
assign micromatrizz[3][603] = 9'b111111111;
assign micromatrizz[3][604] = 9'b111111111;
assign micromatrizz[3][605] = 9'b111111111;
assign micromatrizz[3][606] = 9'b111111111;
assign micromatrizz[3][607] = 9'b111111111;
assign micromatrizz[3][608] = 9'b111111111;
assign micromatrizz[3][609] = 9'b111111111;
assign micromatrizz[3][610] = 9'b111111111;
assign micromatrizz[3][611] = 9'b111111111;
assign micromatrizz[3][612] = 9'b111111111;
assign micromatrizz[3][613] = 9'b111111111;
assign micromatrizz[3][614] = 9'b111111111;
assign micromatrizz[3][615] = 9'b111111111;
assign micromatrizz[3][616] = 9'b111111111;
assign micromatrizz[3][617] = 9'b111111111;
assign micromatrizz[3][618] = 9'b111111111;
assign micromatrizz[3][619] = 9'b111111111;
assign micromatrizz[3][620] = 9'b111111111;
assign micromatrizz[3][621] = 9'b111111111;
assign micromatrizz[3][622] = 9'b111111111;
assign micromatrizz[3][623] = 9'b111111111;
assign micromatrizz[3][624] = 9'b111111111;
assign micromatrizz[3][625] = 9'b111111111;
assign micromatrizz[3][626] = 9'b111111111;
assign micromatrizz[3][627] = 9'b111111111;
assign micromatrizz[3][628] = 9'b111111111;
assign micromatrizz[3][629] = 9'b111111111;
assign micromatrizz[3][630] = 9'b111111111;
assign micromatrizz[3][631] = 9'b111111111;
assign micromatrizz[3][632] = 9'b111111111;
assign micromatrizz[3][633] = 9'b111111111;
assign micromatrizz[3][634] = 9'b111111111;
assign micromatrizz[3][635] = 9'b111111111;
assign micromatrizz[3][636] = 9'b111111111;
assign micromatrizz[3][637] = 9'b111111111;
assign micromatrizz[3][638] = 9'b111111111;
assign micromatrizz[3][639] = 9'b111111111;
assign micromatrizz[4][0] = 9'b111111111;
assign micromatrizz[4][1] = 9'b111111111;
assign micromatrizz[4][2] = 9'b111111111;
assign micromatrizz[4][3] = 9'b111111111;
assign micromatrizz[4][4] = 9'b111111111;
assign micromatrizz[4][5] = 9'b111111111;
assign micromatrizz[4][6] = 9'b111111111;
assign micromatrizz[4][7] = 9'b111111111;
assign micromatrizz[4][8] = 9'b111111111;
assign micromatrizz[4][9] = 9'b111111111;
assign micromatrizz[4][10] = 9'b111111111;
assign micromatrizz[4][11] = 9'b111111111;
assign micromatrizz[4][12] = 9'b111111111;
assign micromatrizz[4][13] = 9'b111111111;
assign micromatrizz[4][14] = 9'b111111111;
assign micromatrizz[4][15] = 9'b111111111;
assign micromatrizz[4][16] = 9'b111111111;
assign micromatrizz[4][17] = 9'b111111111;
assign micromatrizz[4][18] = 9'b111111111;
assign micromatrizz[4][19] = 9'b111111111;
assign micromatrizz[4][20] = 9'b111111111;
assign micromatrizz[4][21] = 9'b111111111;
assign micromatrizz[4][22] = 9'b111111111;
assign micromatrizz[4][23] = 9'b111111111;
assign micromatrizz[4][24] = 9'b111111111;
assign micromatrizz[4][25] = 9'b111111111;
assign micromatrizz[4][26] = 9'b111111111;
assign micromatrizz[4][27] = 9'b111111111;
assign micromatrizz[4][28] = 9'b111111111;
assign micromatrizz[4][29] = 9'b111111111;
assign micromatrizz[4][30] = 9'b111111111;
assign micromatrizz[4][31] = 9'b111111111;
assign micromatrizz[4][32] = 9'b111111111;
assign micromatrizz[4][33] = 9'b111111111;
assign micromatrizz[4][34] = 9'b111111111;
assign micromatrizz[4][35] = 9'b111111111;
assign micromatrizz[4][36] = 9'b111111111;
assign micromatrizz[4][37] = 9'b111111111;
assign micromatrizz[4][38] = 9'b111111111;
assign micromatrizz[4][39] = 9'b111111111;
assign micromatrizz[4][40] = 9'b111111111;
assign micromatrizz[4][41] = 9'b111111111;
assign micromatrizz[4][42] = 9'b111111111;
assign micromatrizz[4][43] = 9'b111111111;
assign micromatrizz[4][44] = 9'b111111111;
assign micromatrizz[4][45] = 9'b111111111;
assign micromatrizz[4][46] = 9'b111111111;
assign micromatrizz[4][47] = 9'b111111111;
assign micromatrizz[4][48] = 9'b111111111;
assign micromatrizz[4][49] = 9'b111111111;
assign micromatrizz[4][50] = 9'b111111111;
assign micromatrizz[4][51] = 9'b111111111;
assign micromatrizz[4][52] = 9'b111111111;
assign micromatrizz[4][53] = 9'b111111111;
assign micromatrizz[4][54] = 9'b111111111;
assign micromatrizz[4][55] = 9'b111111111;
assign micromatrizz[4][56] = 9'b111111111;
assign micromatrizz[4][57] = 9'b111111111;
assign micromatrizz[4][58] = 9'b111111111;
assign micromatrizz[4][59] = 9'b111111111;
assign micromatrizz[4][60] = 9'b111111111;
assign micromatrizz[4][61] = 9'b111111111;
assign micromatrizz[4][62] = 9'b111111111;
assign micromatrizz[4][63] = 9'b111111111;
assign micromatrizz[4][64] = 9'b111111111;
assign micromatrizz[4][65] = 9'b111111111;
assign micromatrizz[4][66] = 9'b111111111;
assign micromatrizz[4][67] = 9'b111111111;
assign micromatrizz[4][68] = 9'b111111111;
assign micromatrizz[4][69] = 9'b111111111;
assign micromatrizz[4][70] = 9'b111111111;
assign micromatrizz[4][71] = 9'b111111111;
assign micromatrizz[4][72] = 9'b111111111;
assign micromatrizz[4][73] = 9'b111111111;
assign micromatrizz[4][74] = 9'b111111111;
assign micromatrizz[4][75] = 9'b111111111;
assign micromatrizz[4][76] = 9'b111111111;
assign micromatrizz[4][77] = 9'b111111111;
assign micromatrizz[4][78] = 9'b111111111;
assign micromatrizz[4][79] = 9'b111111111;
assign micromatrizz[4][80] = 9'b111111111;
assign micromatrizz[4][81] = 9'b111111111;
assign micromatrizz[4][82] = 9'b111111111;
assign micromatrizz[4][83] = 9'b111111111;
assign micromatrizz[4][84] = 9'b111111111;
assign micromatrizz[4][85] = 9'b111111111;
assign micromatrizz[4][86] = 9'b111111111;
assign micromatrizz[4][87] = 9'b111111111;
assign micromatrizz[4][88] = 9'b111111111;
assign micromatrizz[4][89] = 9'b111111111;
assign micromatrizz[4][90] = 9'b111111111;
assign micromatrizz[4][91] = 9'b111111111;
assign micromatrizz[4][92] = 9'b111111111;
assign micromatrizz[4][93] = 9'b111111111;
assign micromatrizz[4][94] = 9'b111111111;
assign micromatrizz[4][95] = 9'b111111111;
assign micromatrizz[4][96] = 9'b111111111;
assign micromatrizz[4][97] = 9'b111111111;
assign micromatrizz[4][98] = 9'b111111111;
assign micromatrizz[4][99] = 9'b111111111;
assign micromatrizz[4][100] = 9'b111111111;
assign micromatrizz[4][101] = 9'b111111111;
assign micromatrizz[4][102] = 9'b111111111;
assign micromatrizz[4][103] = 9'b111111111;
assign micromatrizz[4][104] = 9'b111111111;
assign micromatrizz[4][105] = 9'b111111111;
assign micromatrizz[4][106] = 9'b111111111;
assign micromatrizz[4][107] = 9'b111111111;
assign micromatrizz[4][108] = 9'b111111111;
assign micromatrizz[4][109] = 9'b111111111;
assign micromatrizz[4][110] = 9'b111111111;
assign micromatrizz[4][111] = 9'b111111111;
assign micromatrizz[4][112] = 9'b111111111;
assign micromatrizz[4][113] = 9'b111111111;
assign micromatrizz[4][114] = 9'b111111111;
assign micromatrizz[4][115] = 9'b111111111;
assign micromatrizz[4][116] = 9'b111111111;
assign micromatrizz[4][117] = 9'b111111111;
assign micromatrizz[4][118] = 9'b111111111;
assign micromatrizz[4][119] = 9'b111111111;
assign micromatrizz[4][120] = 9'b111111111;
assign micromatrizz[4][121] = 9'b111111111;
assign micromatrizz[4][122] = 9'b111111111;
assign micromatrizz[4][123] = 9'b111111111;
assign micromatrizz[4][124] = 9'b111111111;
assign micromatrizz[4][125] = 9'b111111111;
assign micromatrizz[4][126] = 9'b111111111;
assign micromatrizz[4][127] = 9'b111111111;
assign micromatrizz[4][128] = 9'b111111111;
assign micromatrizz[4][129] = 9'b111111111;
assign micromatrizz[4][130] = 9'b111111111;
assign micromatrizz[4][131] = 9'b111111111;
assign micromatrizz[4][132] = 9'b111111111;
assign micromatrizz[4][133] = 9'b111111111;
assign micromatrizz[4][134] = 9'b111111111;
assign micromatrizz[4][135] = 9'b111111111;
assign micromatrizz[4][136] = 9'b111111111;
assign micromatrizz[4][137] = 9'b111111111;
assign micromatrizz[4][138] = 9'b111111111;
assign micromatrizz[4][139] = 9'b111111111;
assign micromatrizz[4][140] = 9'b111111111;
assign micromatrizz[4][141] = 9'b111111111;
assign micromatrizz[4][142] = 9'b111111111;
assign micromatrizz[4][143] = 9'b111111111;
assign micromatrizz[4][144] = 9'b111111111;
assign micromatrizz[4][145] = 9'b111111111;
assign micromatrizz[4][146] = 9'b111111111;
assign micromatrizz[4][147] = 9'b111111111;
assign micromatrizz[4][148] = 9'b111111111;
assign micromatrizz[4][149] = 9'b111111111;
assign micromatrizz[4][150] = 9'b111111111;
assign micromatrizz[4][151] = 9'b111111111;
assign micromatrizz[4][152] = 9'b111111111;
assign micromatrizz[4][153] = 9'b111111111;
assign micromatrizz[4][154] = 9'b111111111;
assign micromatrizz[4][155] = 9'b111111111;
assign micromatrizz[4][156] = 9'b111111111;
assign micromatrizz[4][157] = 9'b111111111;
assign micromatrizz[4][158] = 9'b111111111;
assign micromatrizz[4][159] = 9'b111111111;
assign micromatrizz[4][160] = 9'b111111111;
assign micromatrizz[4][161] = 9'b111111111;
assign micromatrizz[4][162] = 9'b111111111;
assign micromatrizz[4][163] = 9'b111111111;
assign micromatrizz[4][164] = 9'b111111111;
assign micromatrizz[4][165] = 9'b111111111;
assign micromatrizz[4][166] = 9'b111111111;
assign micromatrizz[4][167] = 9'b111111111;
assign micromatrizz[4][168] = 9'b111111111;
assign micromatrizz[4][169] = 9'b111111111;
assign micromatrizz[4][170] = 9'b111111111;
assign micromatrizz[4][171] = 9'b111111111;
assign micromatrizz[4][172] = 9'b111111111;
assign micromatrizz[4][173] = 9'b111111111;
assign micromatrizz[4][174] = 9'b111111111;
assign micromatrizz[4][175] = 9'b111111111;
assign micromatrizz[4][176] = 9'b111111111;
assign micromatrizz[4][177] = 9'b111111111;
assign micromatrizz[4][178] = 9'b111111111;
assign micromatrizz[4][179] = 9'b111111111;
assign micromatrizz[4][180] = 9'b111111111;
assign micromatrizz[4][181] = 9'b111111111;
assign micromatrizz[4][182] = 9'b111111111;
assign micromatrizz[4][183] = 9'b111111111;
assign micromatrizz[4][184] = 9'b111111111;
assign micromatrizz[4][185] = 9'b111111111;
assign micromatrizz[4][186] = 9'b111111111;
assign micromatrizz[4][187] = 9'b111111111;
assign micromatrizz[4][188] = 9'b111111111;
assign micromatrizz[4][189] = 9'b111111111;
assign micromatrizz[4][190] = 9'b111111111;
assign micromatrizz[4][191] = 9'b111111111;
assign micromatrizz[4][192] = 9'b111111111;
assign micromatrizz[4][193] = 9'b111111111;
assign micromatrizz[4][194] = 9'b111111111;
assign micromatrizz[4][195] = 9'b111111111;
assign micromatrizz[4][196] = 9'b111111111;
assign micromatrizz[4][197] = 9'b111111111;
assign micromatrizz[4][198] = 9'b111111111;
assign micromatrizz[4][199] = 9'b111111111;
assign micromatrizz[4][200] = 9'b111111111;
assign micromatrizz[4][201] = 9'b111111111;
assign micromatrizz[4][202] = 9'b111111111;
assign micromatrizz[4][203] = 9'b111111111;
assign micromatrizz[4][204] = 9'b111111111;
assign micromatrizz[4][205] = 9'b111111111;
assign micromatrizz[4][206] = 9'b111111111;
assign micromatrizz[4][207] = 9'b111111111;
assign micromatrizz[4][208] = 9'b111111111;
assign micromatrizz[4][209] = 9'b111111111;
assign micromatrizz[4][210] = 9'b111111111;
assign micromatrizz[4][211] = 9'b111111111;
assign micromatrizz[4][212] = 9'b111111111;
assign micromatrizz[4][213] = 9'b111111111;
assign micromatrizz[4][214] = 9'b111111111;
assign micromatrizz[4][215] = 9'b111111111;
assign micromatrizz[4][216] = 9'b111111111;
assign micromatrizz[4][217] = 9'b111111111;
assign micromatrizz[4][218] = 9'b111111111;
assign micromatrizz[4][219] = 9'b111111111;
assign micromatrizz[4][220] = 9'b111111111;
assign micromatrizz[4][221] = 9'b111111111;
assign micromatrizz[4][222] = 9'b111111111;
assign micromatrizz[4][223] = 9'b111111111;
assign micromatrizz[4][224] = 9'b111111111;
assign micromatrizz[4][225] = 9'b111111111;
assign micromatrizz[4][226] = 9'b111111111;
assign micromatrizz[4][227] = 9'b111111111;
assign micromatrizz[4][228] = 9'b111111111;
assign micromatrizz[4][229] = 9'b111111111;
assign micromatrizz[4][230] = 9'b111111111;
assign micromatrizz[4][231] = 9'b111111111;
assign micromatrizz[4][232] = 9'b111111111;
assign micromatrizz[4][233] = 9'b111111111;
assign micromatrizz[4][234] = 9'b111111111;
assign micromatrizz[4][235] = 9'b111111111;
assign micromatrizz[4][236] = 9'b111111111;
assign micromatrizz[4][237] = 9'b111111111;
assign micromatrizz[4][238] = 9'b111111111;
assign micromatrizz[4][239] = 9'b111111111;
assign micromatrizz[4][240] = 9'b111111111;
assign micromatrizz[4][241] = 9'b111111111;
assign micromatrizz[4][242] = 9'b111111111;
assign micromatrizz[4][243] = 9'b111111111;
assign micromatrizz[4][244] = 9'b111111111;
assign micromatrizz[4][245] = 9'b111111111;
assign micromatrizz[4][246] = 9'b111111111;
assign micromatrizz[4][247] = 9'b111111111;
assign micromatrizz[4][248] = 9'b111111111;
assign micromatrizz[4][249] = 9'b111111111;
assign micromatrizz[4][250] = 9'b111111111;
assign micromatrizz[4][251] = 9'b111111111;
assign micromatrizz[4][252] = 9'b111111111;
assign micromatrizz[4][253] = 9'b111111111;
assign micromatrizz[4][254] = 9'b111111111;
assign micromatrizz[4][255] = 9'b111111111;
assign micromatrizz[4][256] = 9'b111111111;
assign micromatrizz[4][257] = 9'b111111111;
assign micromatrizz[4][258] = 9'b111111111;
assign micromatrizz[4][259] = 9'b111111111;
assign micromatrizz[4][260] = 9'b111111111;
assign micromatrizz[4][261] = 9'b111111111;
assign micromatrizz[4][262] = 9'b111111111;
assign micromatrizz[4][263] = 9'b111111111;
assign micromatrizz[4][264] = 9'b111111111;
assign micromatrizz[4][265] = 9'b111111111;
assign micromatrizz[4][266] = 9'b111111111;
assign micromatrizz[4][267] = 9'b111111111;
assign micromatrizz[4][268] = 9'b111111111;
assign micromatrizz[4][269] = 9'b111111111;
assign micromatrizz[4][270] = 9'b111111111;
assign micromatrizz[4][271] = 9'b111111111;
assign micromatrizz[4][272] = 9'b111111111;
assign micromatrizz[4][273] = 9'b111111111;
assign micromatrizz[4][274] = 9'b111111111;
assign micromatrizz[4][275] = 9'b111111111;
assign micromatrizz[4][276] = 9'b111111111;
assign micromatrizz[4][277] = 9'b111111111;
assign micromatrizz[4][278] = 9'b111111111;
assign micromatrizz[4][279] = 9'b111111111;
assign micromatrizz[4][280] = 9'b111111111;
assign micromatrizz[4][281] = 9'b111111111;
assign micromatrizz[4][282] = 9'b111111111;
assign micromatrizz[4][283] = 9'b111111111;
assign micromatrizz[4][284] = 9'b111111111;
assign micromatrizz[4][285] = 9'b111111111;
assign micromatrizz[4][286] = 9'b111111111;
assign micromatrizz[4][287] = 9'b111111111;
assign micromatrizz[4][288] = 9'b111111111;
assign micromatrizz[4][289] = 9'b111111111;
assign micromatrizz[4][290] = 9'b111111111;
assign micromatrizz[4][291] = 9'b111111111;
assign micromatrizz[4][292] = 9'b111111111;
assign micromatrizz[4][293] = 9'b111111111;
assign micromatrizz[4][294] = 9'b111111111;
assign micromatrizz[4][295] = 9'b111111111;
assign micromatrizz[4][296] = 9'b111111111;
assign micromatrizz[4][297] = 9'b111111111;
assign micromatrizz[4][298] = 9'b111111111;
assign micromatrizz[4][299] = 9'b111111111;
assign micromatrizz[4][300] = 9'b111111111;
assign micromatrizz[4][301] = 9'b111111111;
assign micromatrizz[4][302] = 9'b111111111;
assign micromatrizz[4][303] = 9'b111111111;
assign micromatrizz[4][304] = 9'b111111111;
assign micromatrizz[4][305] = 9'b111111111;
assign micromatrizz[4][306] = 9'b111111111;
assign micromatrizz[4][307] = 9'b111111111;
assign micromatrizz[4][308] = 9'b111111111;
assign micromatrizz[4][309] = 9'b111111111;
assign micromatrizz[4][310] = 9'b111111111;
assign micromatrizz[4][311] = 9'b111111111;
assign micromatrizz[4][312] = 9'b111111111;
assign micromatrizz[4][313] = 9'b111111111;
assign micromatrizz[4][314] = 9'b111111111;
assign micromatrizz[4][315] = 9'b111111111;
assign micromatrizz[4][316] = 9'b111111111;
assign micromatrizz[4][317] = 9'b111111111;
assign micromatrizz[4][318] = 9'b111111111;
assign micromatrizz[4][319] = 9'b111111111;
assign micromatrizz[4][320] = 9'b111111111;
assign micromatrizz[4][321] = 9'b111111111;
assign micromatrizz[4][322] = 9'b111111111;
assign micromatrizz[4][323] = 9'b111111111;
assign micromatrizz[4][324] = 9'b111111111;
assign micromatrizz[4][325] = 9'b111111111;
assign micromatrizz[4][326] = 9'b111111111;
assign micromatrizz[4][327] = 9'b111111111;
assign micromatrizz[4][328] = 9'b111111111;
assign micromatrizz[4][329] = 9'b111111111;
assign micromatrizz[4][330] = 9'b111111111;
assign micromatrizz[4][331] = 9'b111111111;
assign micromatrizz[4][332] = 9'b111111111;
assign micromatrizz[4][333] = 9'b111111111;
assign micromatrizz[4][334] = 9'b111111111;
assign micromatrizz[4][335] = 9'b111111111;
assign micromatrizz[4][336] = 9'b111111111;
assign micromatrizz[4][337] = 9'b111111111;
assign micromatrizz[4][338] = 9'b111111111;
assign micromatrizz[4][339] = 9'b111111111;
assign micromatrizz[4][340] = 9'b111111111;
assign micromatrizz[4][341] = 9'b111111111;
assign micromatrizz[4][342] = 9'b111111111;
assign micromatrizz[4][343] = 9'b111111111;
assign micromatrizz[4][344] = 9'b111111111;
assign micromatrizz[4][345] = 9'b111111111;
assign micromatrizz[4][346] = 9'b111111111;
assign micromatrizz[4][347] = 9'b111111111;
assign micromatrizz[4][348] = 9'b111111111;
assign micromatrizz[4][349] = 9'b111111111;
assign micromatrizz[4][350] = 9'b111111111;
assign micromatrizz[4][351] = 9'b111111111;
assign micromatrizz[4][352] = 9'b111111111;
assign micromatrizz[4][353] = 9'b111111111;
assign micromatrizz[4][354] = 9'b111111111;
assign micromatrizz[4][355] = 9'b111111111;
assign micromatrizz[4][356] = 9'b111111111;
assign micromatrizz[4][357] = 9'b111111111;
assign micromatrizz[4][358] = 9'b111111111;
assign micromatrizz[4][359] = 9'b111111111;
assign micromatrizz[4][360] = 9'b111111111;
assign micromatrizz[4][361] = 9'b111111111;
assign micromatrizz[4][362] = 9'b111111111;
assign micromatrizz[4][363] = 9'b111111111;
assign micromatrizz[4][364] = 9'b111111111;
assign micromatrizz[4][365] = 9'b111111111;
assign micromatrizz[4][366] = 9'b111111111;
assign micromatrizz[4][367] = 9'b111111111;
assign micromatrizz[4][368] = 9'b111111111;
assign micromatrizz[4][369] = 9'b111111111;
assign micromatrizz[4][370] = 9'b111111111;
assign micromatrizz[4][371] = 9'b111111111;
assign micromatrizz[4][372] = 9'b111111111;
assign micromatrizz[4][373] = 9'b111111111;
assign micromatrizz[4][374] = 9'b111111111;
assign micromatrizz[4][375] = 9'b111111111;
assign micromatrizz[4][376] = 9'b111111111;
assign micromatrizz[4][377] = 9'b111111111;
assign micromatrizz[4][378] = 9'b111111111;
assign micromatrizz[4][379] = 9'b111111111;
assign micromatrizz[4][380] = 9'b111111111;
assign micromatrizz[4][381] = 9'b111111111;
assign micromatrizz[4][382] = 9'b111111111;
assign micromatrizz[4][383] = 9'b111111111;
assign micromatrizz[4][384] = 9'b111111111;
assign micromatrizz[4][385] = 9'b111111111;
assign micromatrizz[4][386] = 9'b111111111;
assign micromatrizz[4][387] = 9'b111111111;
assign micromatrizz[4][388] = 9'b111111111;
assign micromatrizz[4][389] = 9'b111111111;
assign micromatrizz[4][390] = 9'b111111111;
assign micromatrizz[4][391] = 9'b111111111;
assign micromatrizz[4][392] = 9'b111111111;
assign micromatrizz[4][393] = 9'b111111111;
assign micromatrizz[4][394] = 9'b111111111;
assign micromatrizz[4][395] = 9'b111111111;
assign micromatrizz[4][396] = 9'b111111111;
assign micromatrizz[4][397] = 9'b111111111;
assign micromatrizz[4][398] = 9'b111111111;
assign micromatrizz[4][399] = 9'b111111111;
assign micromatrizz[4][400] = 9'b111111111;
assign micromatrizz[4][401] = 9'b111111111;
assign micromatrizz[4][402] = 9'b111111111;
assign micromatrizz[4][403] = 9'b111111111;
assign micromatrizz[4][404] = 9'b111111111;
assign micromatrizz[4][405] = 9'b111111111;
assign micromatrizz[4][406] = 9'b111111111;
assign micromatrizz[4][407] = 9'b111111111;
assign micromatrizz[4][408] = 9'b111111111;
assign micromatrizz[4][409] = 9'b111111111;
assign micromatrizz[4][410] = 9'b111111111;
assign micromatrizz[4][411] = 9'b111111111;
assign micromatrizz[4][412] = 9'b111111111;
assign micromatrizz[4][413] = 9'b111111111;
assign micromatrizz[4][414] = 9'b111111111;
assign micromatrizz[4][415] = 9'b111111111;
assign micromatrizz[4][416] = 9'b111111111;
assign micromatrizz[4][417] = 9'b111111111;
assign micromatrizz[4][418] = 9'b111111111;
assign micromatrizz[4][419] = 9'b111111111;
assign micromatrizz[4][420] = 9'b111111111;
assign micromatrizz[4][421] = 9'b111111111;
assign micromatrizz[4][422] = 9'b111111111;
assign micromatrizz[4][423] = 9'b111111111;
assign micromatrizz[4][424] = 9'b111111111;
assign micromatrizz[4][425] = 9'b111111111;
assign micromatrizz[4][426] = 9'b111111111;
assign micromatrizz[4][427] = 9'b111111111;
assign micromatrizz[4][428] = 9'b111111111;
assign micromatrizz[4][429] = 9'b111111111;
assign micromatrizz[4][430] = 9'b111111111;
assign micromatrizz[4][431] = 9'b111111111;
assign micromatrizz[4][432] = 9'b111111111;
assign micromatrizz[4][433] = 9'b111111111;
assign micromatrizz[4][434] = 9'b111111111;
assign micromatrizz[4][435] = 9'b111111111;
assign micromatrizz[4][436] = 9'b111111111;
assign micromatrizz[4][437] = 9'b111111111;
assign micromatrizz[4][438] = 9'b111111111;
assign micromatrizz[4][439] = 9'b111111111;
assign micromatrizz[4][440] = 9'b111111111;
assign micromatrizz[4][441] = 9'b111111111;
assign micromatrizz[4][442] = 9'b111111111;
assign micromatrizz[4][443] = 9'b111111111;
assign micromatrizz[4][444] = 9'b111111111;
assign micromatrizz[4][445] = 9'b111111111;
assign micromatrizz[4][446] = 9'b111111111;
assign micromatrizz[4][447] = 9'b111111111;
assign micromatrizz[4][448] = 9'b111111111;
assign micromatrizz[4][449] = 9'b111111111;
assign micromatrizz[4][450] = 9'b111111111;
assign micromatrizz[4][451] = 9'b111111111;
assign micromatrizz[4][452] = 9'b111111111;
assign micromatrizz[4][453] = 9'b111111111;
assign micromatrizz[4][454] = 9'b111111111;
assign micromatrizz[4][455] = 9'b111111111;
assign micromatrizz[4][456] = 9'b111111111;
assign micromatrizz[4][457] = 9'b111111111;
assign micromatrizz[4][458] = 9'b111111111;
assign micromatrizz[4][459] = 9'b111111111;
assign micromatrizz[4][460] = 9'b111111111;
assign micromatrizz[4][461] = 9'b111111111;
assign micromatrizz[4][462] = 9'b111111111;
assign micromatrizz[4][463] = 9'b111111111;
assign micromatrizz[4][464] = 9'b111111111;
assign micromatrizz[4][465] = 9'b111111111;
assign micromatrizz[4][466] = 9'b111111111;
assign micromatrizz[4][467] = 9'b111111111;
assign micromatrizz[4][468] = 9'b111111111;
assign micromatrizz[4][469] = 9'b111111111;
assign micromatrizz[4][470] = 9'b111111111;
assign micromatrizz[4][471] = 9'b111111111;
assign micromatrizz[4][472] = 9'b111111111;
assign micromatrizz[4][473] = 9'b111111111;
assign micromatrizz[4][474] = 9'b111111111;
assign micromatrizz[4][475] = 9'b111111111;
assign micromatrizz[4][476] = 9'b111111111;
assign micromatrizz[4][477] = 9'b111111111;
assign micromatrizz[4][478] = 9'b111111111;
assign micromatrizz[4][479] = 9'b111111111;
assign micromatrizz[4][480] = 9'b111111111;
assign micromatrizz[4][481] = 9'b111111111;
assign micromatrizz[4][482] = 9'b111111111;
assign micromatrizz[4][483] = 9'b111111111;
assign micromatrizz[4][484] = 9'b111111111;
assign micromatrizz[4][485] = 9'b111111111;
assign micromatrizz[4][486] = 9'b111111111;
assign micromatrizz[4][487] = 9'b111111111;
assign micromatrizz[4][488] = 9'b111111111;
assign micromatrizz[4][489] = 9'b111111111;
assign micromatrizz[4][490] = 9'b111111111;
assign micromatrizz[4][491] = 9'b111111111;
assign micromatrizz[4][492] = 9'b111111111;
assign micromatrizz[4][493] = 9'b111111111;
assign micromatrizz[4][494] = 9'b111111111;
assign micromatrizz[4][495] = 9'b111111111;
assign micromatrizz[4][496] = 9'b111111111;
assign micromatrizz[4][497] = 9'b111111111;
assign micromatrizz[4][498] = 9'b111111111;
assign micromatrizz[4][499] = 9'b111111111;
assign micromatrizz[4][500] = 9'b111111111;
assign micromatrizz[4][501] = 9'b111111111;
assign micromatrizz[4][502] = 9'b111111111;
assign micromatrizz[4][503] = 9'b111111111;
assign micromatrizz[4][504] = 9'b111111111;
assign micromatrizz[4][505] = 9'b111111111;
assign micromatrizz[4][506] = 9'b111111111;
assign micromatrizz[4][507] = 9'b111111111;
assign micromatrizz[4][508] = 9'b111111111;
assign micromatrizz[4][509] = 9'b111111111;
assign micromatrizz[4][510] = 9'b111111111;
assign micromatrizz[4][511] = 9'b111111111;
assign micromatrizz[4][512] = 9'b111111111;
assign micromatrizz[4][513] = 9'b111111111;
assign micromatrizz[4][514] = 9'b111111111;
assign micromatrizz[4][515] = 9'b111111111;
assign micromatrizz[4][516] = 9'b111111111;
assign micromatrizz[4][517] = 9'b111111111;
assign micromatrizz[4][518] = 9'b111111111;
assign micromatrizz[4][519] = 9'b111111111;
assign micromatrizz[4][520] = 9'b111111111;
assign micromatrizz[4][521] = 9'b111111111;
assign micromatrizz[4][522] = 9'b111111111;
assign micromatrizz[4][523] = 9'b111111111;
assign micromatrizz[4][524] = 9'b111111111;
assign micromatrizz[4][525] = 9'b111111111;
assign micromatrizz[4][526] = 9'b111111111;
assign micromatrizz[4][527] = 9'b111111111;
assign micromatrizz[4][528] = 9'b111111111;
assign micromatrizz[4][529] = 9'b111111111;
assign micromatrizz[4][530] = 9'b111111111;
assign micromatrizz[4][531] = 9'b111111111;
assign micromatrizz[4][532] = 9'b111111111;
assign micromatrizz[4][533] = 9'b111111111;
assign micromatrizz[4][534] = 9'b111111111;
assign micromatrizz[4][535] = 9'b111111111;
assign micromatrizz[4][536] = 9'b111111111;
assign micromatrizz[4][537] = 9'b111111111;
assign micromatrizz[4][538] = 9'b111111111;
assign micromatrizz[4][539] = 9'b111111111;
assign micromatrizz[4][540] = 9'b111111111;
assign micromatrizz[4][541] = 9'b111111111;
assign micromatrizz[4][542] = 9'b111111111;
assign micromatrizz[4][543] = 9'b111111111;
assign micromatrizz[4][544] = 9'b111111111;
assign micromatrizz[4][545] = 9'b111111111;
assign micromatrizz[4][546] = 9'b111111111;
assign micromatrizz[4][547] = 9'b111111111;
assign micromatrizz[4][548] = 9'b111111111;
assign micromatrizz[4][549] = 9'b111111111;
assign micromatrizz[4][550] = 9'b111111111;
assign micromatrizz[4][551] = 9'b111111111;
assign micromatrizz[4][552] = 9'b111111111;
assign micromatrizz[4][553] = 9'b111111111;
assign micromatrizz[4][554] = 9'b111111111;
assign micromatrizz[4][555] = 9'b111111111;
assign micromatrizz[4][556] = 9'b111111111;
assign micromatrizz[4][557] = 9'b111111111;
assign micromatrizz[4][558] = 9'b111111111;
assign micromatrizz[4][559] = 9'b111111111;
assign micromatrizz[4][560] = 9'b111111111;
assign micromatrizz[4][561] = 9'b111111111;
assign micromatrizz[4][562] = 9'b111111111;
assign micromatrizz[4][563] = 9'b111111111;
assign micromatrizz[4][564] = 9'b111111111;
assign micromatrizz[4][565] = 9'b111111111;
assign micromatrizz[4][566] = 9'b111111111;
assign micromatrizz[4][567] = 9'b111111111;
assign micromatrizz[4][568] = 9'b111111111;
assign micromatrizz[4][569] = 9'b111111111;
assign micromatrizz[4][570] = 9'b111111111;
assign micromatrizz[4][571] = 9'b111111111;
assign micromatrizz[4][572] = 9'b111111111;
assign micromatrizz[4][573] = 9'b111111111;
assign micromatrizz[4][574] = 9'b111111111;
assign micromatrizz[4][575] = 9'b111111111;
assign micromatrizz[4][576] = 9'b111111111;
assign micromatrizz[4][577] = 9'b111111111;
assign micromatrizz[4][578] = 9'b111111111;
assign micromatrizz[4][579] = 9'b111111111;
assign micromatrizz[4][580] = 9'b111111111;
assign micromatrizz[4][581] = 9'b111111111;
assign micromatrizz[4][582] = 9'b111111111;
assign micromatrizz[4][583] = 9'b111111111;
assign micromatrizz[4][584] = 9'b111111111;
assign micromatrizz[4][585] = 9'b111111111;
assign micromatrizz[4][586] = 9'b111111111;
assign micromatrizz[4][587] = 9'b111111111;
assign micromatrizz[4][588] = 9'b111111111;
assign micromatrizz[4][589] = 9'b111111111;
assign micromatrizz[4][590] = 9'b111111111;
assign micromatrizz[4][591] = 9'b111111111;
assign micromatrizz[4][592] = 9'b111111111;
assign micromatrizz[4][593] = 9'b111111111;
assign micromatrizz[4][594] = 9'b111111111;
assign micromatrizz[4][595] = 9'b111111111;
assign micromatrizz[4][596] = 9'b111111111;
assign micromatrizz[4][597] = 9'b111111111;
assign micromatrizz[4][598] = 9'b111111111;
assign micromatrizz[4][599] = 9'b111111111;
assign micromatrizz[4][600] = 9'b111111111;
assign micromatrizz[4][601] = 9'b111111111;
assign micromatrizz[4][602] = 9'b111111111;
assign micromatrizz[4][603] = 9'b111111111;
assign micromatrizz[4][604] = 9'b111111111;
assign micromatrizz[4][605] = 9'b111111111;
assign micromatrizz[4][606] = 9'b111111111;
assign micromatrizz[4][607] = 9'b111111111;
assign micromatrizz[4][608] = 9'b111111111;
assign micromatrizz[4][609] = 9'b111111111;
assign micromatrizz[4][610] = 9'b111111111;
assign micromatrizz[4][611] = 9'b111111111;
assign micromatrizz[4][612] = 9'b111111111;
assign micromatrizz[4][613] = 9'b111111111;
assign micromatrizz[4][614] = 9'b111111111;
assign micromatrizz[4][615] = 9'b111111111;
assign micromatrizz[4][616] = 9'b111111111;
assign micromatrizz[4][617] = 9'b111111111;
assign micromatrizz[4][618] = 9'b111111111;
assign micromatrizz[4][619] = 9'b111111111;
assign micromatrizz[4][620] = 9'b111111111;
assign micromatrizz[4][621] = 9'b111111111;
assign micromatrizz[4][622] = 9'b111111111;
assign micromatrizz[4][623] = 9'b111111111;
assign micromatrizz[4][624] = 9'b111111111;
assign micromatrizz[4][625] = 9'b111111111;
assign micromatrizz[4][626] = 9'b111111111;
assign micromatrizz[4][627] = 9'b111111111;
assign micromatrizz[4][628] = 9'b111111111;
assign micromatrizz[4][629] = 9'b111111111;
assign micromatrizz[4][630] = 9'b111111111;
assign micromatrizz[4][631] = 9'b111111111;
assign micromatrizz[4][632] = 9'b111111111;
assign micromatrizz[4][633] = 9'b111111111;
assign micromatrizz[4][634] = 9'b111111111;
assign micromatrizz[4][635] = 9'b111111111;
assign micromatrizz[4][636] = 9'b111111111;
assign micromatrizz[4][637] = 9'b111111111;
assign micromatrizz[4][638] = 9'b111111111;
assign micromatrizz[4][639] = 9'b111111111;
assign micromatrizz[5][0] = 9'b111111111;
assign micromatrizz[5][1] = 9'b111111111;
assign micromatrizz[5][2] = 9'b111111111;
assign micromatrizz[5][3] = 9'b111111111;
assign micromatrizz[5][4] = 9'b111111111;
assign micromatrizz[5][5] = 9'b111111111;
assign micromatrizz[5][6] = 9'b111111111;
assign micromatrizz[5][7] = 9'b111111111;
assign micromatrizz[5][8] = 9'b111111111;
assign micromatrizz[5][9] = 9'b111111111;
assign micromatrizz[5][10] = 9'b111111111;
assign micromatrizz[5][11] = 9'b111111111;
assign micromatrizz[5][12] = 9'b111111111;
assign micromatrizz[5][13] = 9'b111111111;
assign micromatrizz[5][14] = 9'b111111111;
assign micromatrizz[5][15] = 9'b111111111;
assign micromatrizz[5][16] = 9'b111111111;
assign micromatrizz[5][17] = 9'b111111111;
assign micromatrizz[5][18] = 9'b111111111;
assign micromatrizz[5][19] = 9'b111111111;
assign micromatrizz[5][20] = 9'b111111111;
assign micromatrizz[5][21] = 9'b111111111;
assign micromatrizz[5][22] = 9'b111111111;
assign micromatrizz[5][23] = 9'b111111111;
assign micromatrizz[5][24] = 9'b111111111;
assign micromatrizz[5][25] = 9'b111111111;
assign micromatrizz[5][26] = 9'b111111111;
assign micromatrizz[5][27] = 9'b111111111;
assign micromatrizz[5][28] = 9'b111111111;
assign micromatrizz[5][29] = 9'b111111111;
assign micromatrizz[5][30] = 9'b111111111;
assign micromatrizz[5][31] = 9'b111111111;
assign micromatrizz[5][32] = 9'b111111111;
assign micromatrizz[5][33] = 9'b111111111;
assign micromatrizz[5][34] = 9'b111111111;
assign micromatrizz[5][35] = 9'b111111111;
assign micromatrizz[5][36] = 9'b111111111;
assign micromatrizz[5][37] = 9'b111111111;
assign micromatrizz[5][38] = 9'b111111111;
assign micromatrizz[5][39] = 9'b111111111;
assign micromatrizz[5][40] = 9'b111111111;
assign micromatrizz[5][41] = 9'b111111111;
assign micromatrizz[5][42] = 9'b111111111;
assign micromatrizz[5][43] = 9'b111111111;
assign micromatrizz[5][44] = 9'b111111111;
assign micromatrizz[5][45] = 9'b111111111;
assign micromatrizz[5][46] = 9'b111111111;
assign micromatrizz[5][47] = 9'b111111111;
assign micromatrizz[5][48] = 9'b111111111;
assign micromatrizz[5][49] = 9'b111111111;
assign micromatrizz[5][50] = 9'b111111111;
assign micromatrizz[5][51] = 9'b111111111;
assign micromatrizz[5][52] = 9'b111111111;
assign micromatrizz[5][53] = 9'b111111111;
assign micromatrizz[5][54] = 9'b111111111;
assign micromatrizz[5][55] = 9'b111111111;
assign micromatrizz[5][56] = 9'b111111111;
assign micromatrizz[5][57] = 9'b111111111;
assign micromatrizz[5][58] = 9'b111111111;
assign micromatrizz[5][59] = 9'b111111111;
assign micromatrizz[5][60] = 9'b111111111;
assign micromatrizz[5][61] = 9'b111111111;
assign micromatrizz[5][62] = 9'b111111111;
assign micromatrizz[5][63] = 9'b111111111;
assign micromatrizz[5][64] = 9'b111111111;
assign micromatrizz[5][65] = 9'b111111111;
assign micromatrizz[5][66] = 9'b111111111;
assign micromatrizz[5][67] = 9'b111111111;
assign micromatrizz[5][68] = 9'b111111111;
assign micromatrizz[5][69] = 9'b111111111;
assign micromatrizz[5][70] = 9'b111111111;
assign micromatrizz[5][71] = 9'b111111111;
assign micromatrizz[5][72] = 9'b111111111;
assign micromatrizz[5][73] = 9'b111111111;
assign micromatrizz[5][74] = 9'b111111111;
assign micromatrizz[5][75] = 9'b111111111;
assign micromatrizz[5][76] = 9'b111111111;
assign micromatrizz[5][77] = 9'b111111111;
assign micromatrizz[5][78] = 9'b111111111;
assign micromatrizz[5][79] = 9'b111111111;
assign micromatrizz[5][80] = 9'b111111111;
assign micromatrizz[5][81] = 9'b111111111;
assign micromatrizz[5][82] = 9'b111111111;
assign micromatrizz[5][83] = 9'b111111111;
assign micromatrizz[5][84] = 9'b111111111;
assign micromatrizz[5][85] = 9'b111111111;
assign micromatrizz[5][86] = 9'b111111111;
assign micromatrizz[5][87] = 9'b111111111;
assign micromatrizz[5][88] = 9'b111111111;
assign micromatrizz[5][89] = 9'b111111111;
assign micromatrizz[5][90] = 9'b111111111;
assign micromatrizz[5][91] = 9'b111111111;
assign micromatrizz[5][92] = 9'b111111111;
assign micromatrizz[5][93] = 9'b111111111;
assign micromatrizz[5][94] = 9'b111111111;
assign micromatrizz[5][95] = 9'b111111111;
assign micromatrizz[5][96] = 9'b111111111;
assign micromatrizz[5][97] = 9'b111111111;
assign micromatrizz[5][98] = 9'b111111111;
assign micromatrizz[5][99] = 9'b111111111;
assign micromatrizz[5][100] = 9'b111111111;
assign micromatrizz[5][101] = 9'b111111111;
assign micromatrizz[5][102] = 9'b111111111;
assign micromatrizz[5][103] = 9'b111111111;
assign micromatrizz[5][104] = 9'b111111111;
assign micromatrizz[5][105] = 9'b111111111;
assign micromatrizz[5][106] = 9'b111111111;
assign micromatrizz[5][107] = 9'b111111111;
assign micromatrizz[5][108] = 9'b111111111;
assign micromatrizz[5][109] = 9'b111111111;
assign micromatrizz[5][110] = 9'b111111111;
assign micromatrizz[5][111] = 9'b111111111;
assign micromatrizz[5][112] = 9'b111111111;
assign micromatrizz[5][113] = 9'b111111111;
assign micromatrizz[5][114] = 9'b111111111;
assign micromatrizz[5][115] = 9'b111111111;
assign micromatrizz[5][116] = 9'b111111111;
assign micromatrizz[5][117] = 9'b111111111;
assign micromatrizz[5][118] = 9'b111111111;
assign micromatrizz[5][119] = 9'b111111111;
assign micromatrizz[5][120] = 9'b111111111;
assign micromatrizz[5][121] = 9'b111111111;
assign micromatrizz[5][122] = 9'b111111111;
assign micromatrizz[5][123] = 9'b111111111;
assign micromatrizz[5][124] = 9'b111111111;
assign micromatrizz[5][125] = 9'b111111111;
assign micromatrizz[5][126] = 9'b111111111;
assign micromatrizz[5][127] = 9'b111111111;
assign micromatrizz[5][128] = 9'b111111111;
assign micromatrizz[5][129] = 9'b111111111;
assign micromatrizz[5][130] = 9'b111111111;
assign micromatrizz[5][131] = 9'b111111111;
assign micromatrizz[5][132] = 9'b111111111;
assign micromatrizz[5][133] = 9'b111111111;
assign micromatrizz[5][134] = 9'b111111111;
assign micromatrizz[5][135] = 9'b111111111;
assign micromatrizz[5][136] = 9'b111111111;
assign micromatrizz[5][137] = 9'b111111111;
assign micromatrizz[5][138] = 9'b111111111;
assign micromatrizz[5][139] = 9'b111111111;
assign micromatrizz[5][140] = 9'b111111111;
assign micromatrizz[5][141] = 9'b111111111;
assign micromatrizz[5][142] = 9'b111111111;
assign micromatrizz[5][143] = 9'b111111111;
assign micromatrizz[5][144] = 9'b111111111;
assign micromatrizz[5][145] = 9'b111111111;
assign micromatrizz[5][146] = 9'b111111111;
assign micromatrizz[5][147] = 9'b111111111;
assign micromatrizz[5][148] = 9'b111111111;
assign micromatrizz[5][149] = 9'b111111111;
assign micromatrizz[5][150] = 9'b111111111;
assign micromatrizz[5][151] = 9'b111111111;
assign micromatrizz[5][152] = 9'b111111111;
assign micromatrizz[5][153] = 9'b111111111;
assign micromatrizz[5][154] = 9'b111111111;
assign micromatrizz[5][155] = 9'b111111111;
assign micromatrizz[5][156] = 9'b111111111;
assign micromatrizz[5][157] = 9'b111111111;
assign micromatrizz[5][158] = 9'b111111111;
assign micromatrizz[5][159] = 9'b111111111;
assign micromatrizz[5][160] = 9'b111111111;
assign micromatrizz[5][161] = 9'b111111111;
assign micromatrizz[5][162] = 9'b111111111;
assign micromatrizz[5][163] = 9'b111111111;
assign micromatrizz[5][164] = 9'b111111111;
assign micromatrizz[5][165] = 9'b111111111;
assign micromatrizz[5][166] = 9'b111111111;
assign micromatrizz[5][167] = 9'b111111111;
assign micromatrizz[5][168] = 9'b111111111;
assign micromatrizz[5][169] = 9'b111111111;
assign micromatrizz[5][170] = 9'b111111111;
assign micromatrizz[5][171] = 9'b111111111;
assign micromatrizz[5][172] = 9'b111111111;
assign micromatrizz[5][173] = 9'b111111111;
assign micromatrizz[5][174] = 9'b111111111;
assign micromatrizz[5][175] = 9'b111111111;
assign micromatrizz[5][176] = 9'b111111111;
assign micromatrizz[5][177] = 9'b111111111;
assign micromatrizz[5][178] = 9'b111111111;
assign micromatrizz[5][179] = 9'b111111111;
assign micromatrizz[5][180] = 9'b111111111;
assign micromatrizz[5][181] = 9'b111111111;
assign micromatrizz[5][182] = 9'b111111111;
assign micromatrizz[5][183] = 9'b111111111;
assign micromatrizz[5][184] = 9'b111111111;
assign micromatrizz[5][185] = 9'b111111111;
assign micromatrizz[5][186] = 9'b111111111;
assign micromatrizz[5][187] = 9'b111111111;
assign micromatrizz[5][188] = 9'b111111111;
assign micromatrizz[5][189] = 9'b111111111;
assign micromatrizz[5][190] = 9'b111111111;
assign micromatrizz[5][191] = 9'b111111111;
assign micromatrizz[5][192] = 9'b111111111;
assign micromatrizz[5][193] = 9'b111111111;
assign micromatrizz[5][194] = 9'b111111111;
assign micromatrizz[5][195] = 9'b111111111;
assign micromatrizz[5][196] = 9'b111111111;
assign micromatrizz[5][197] = 9'b111111111;
assign micromatrizz[5][198] = 9'b111111111;
assign micromatrizz[5][199] = 9'b111111111;
assign micromatrizz[5][200] = 9'b111111111;
assign micromatrizz[5][201] = 9'b111111111;
assign micromatrizz[5][202] = 9'b111111111;
assign micromatrizz[5][203] = 9'b111111111;
assign micromatrizz[5][204] = 9'b111111111;
assign micromatrizz[5][205] = 9'b111111111;
assign micromatrizz[5][206] = 9'b111111111;
assign micromatrizz[5][207] = 9'b111111111;
assign micromatrizz[5][208] = 9'b111111111;
assign micromatrizz[5][209] = 9'b111111111;
assign micromatrizz[5][210] = 9'b111111111;
assign micromatrizz[5][211] = 9'b111111111;
assign micromatrizz[5][212] = 9'b111111111;
assign micromatrizz[5][213] = 9'b111111111;
assign micromatrizz[5][214] = 9'b111111111;
assign micromatrizz[5][215] = 9'b111111111;
assign micromatrizz[5][216] = 9'b111111111;
assign micromatrizz[5][217] = 9'b111111111;
assign micromatrizz[5][218] = 9'b111111111;
assign micromatrizz[5][219] = 9'b111111111;
assign micromatrizz[5][220] = 9'b111111111;
assign micromatrizz[5][221] = 9'b111111111;
assign micromatrizz[5][222] = 9'b111111111;
assign micromatrizz[5][223] = 9'b111111111;
assign micromatrizz[5][224] = 9'b111111111;
assign micromatrizz[5][225] = 9'b111111111;
assign micromatrizz[5][226] = 9'b111111111;
assign micromatrizz[5][227] = 9'b111111111;
assign micromatrizz[5][228] = 9'b111111111;
assign micromatrizz[5][229] = 9'b111111111;
assign micromatrizz[5][230] = 9'b111111111;
assign micromatrizz[5][231] = 9'b111111111;
assign micromatrizz[5][232] = 9'b111111111;
assign micromatrizz[5][233] = 9'b111111111;
assign micromatrizz[5][234] = 9'b111111111;
assign micromatrizz[5][235] = 9'b111111111;
assign micromatrizz[5][236] = 9'b111111111;
assign micromatrizz[5][237] = 9'b111111111;
assign micromatrizz[5][238] = 9'b111111111;
assign micromatrizz[5][239] = 9'b111111111;
assign micromatrizz[5][240] = 9'b111111111;
assign micromatrizz[5][241] = 9'b111111111;
assign micromatrizz[5][242] = 9'b111111111;
assign micromatrizz[5][243] = 9'b111111111;
assign micromatrizz[5][244] = 9'b111111111;
assign micromatrizz[5][245] = 9'b111111111;
assign micromatrizz[5][246] = 9'b111111111;
assign micromatrizz[5][247] = 9'b111111111;
assign micromatrizz[5][248] = 9'b111111111;
assign micromatrizz[5][249] = 9'b111111111;
assign micromatrizz[5][250] = 9'b111111111;
assign micromatrizz[5][251] = 9'b111111111;
assign micromatrizz[5][252] = 9'b111111111;
assign micromatrizz[5][253] = 9'b111111111;
assign micromatrizz[5][254] = 9'b111111111;
assign micromatrizz[5][255] = 9'b111111111;
assign micromatrizz[5][256] = 9'b111111111;
assign micromatrizz[5][257] = 9'b111111111;
assign micromatrizz[5][258] = 9'b111111111;
assign micromatrizz[5][259] = 9'b111111111;
assign micromatrizz[5][260] = 9'b111111111;
assign micromatrizz[5][261] = 9'b111111111;
assign micromatrizz[5][262] = 9'b111111111;
assign micromatrizz[5][263] = 9'b111111111;
assign micromatrizz[5][264] = 9'b111111111;
assign micromatrizz[5][265] = 9'b111111111;
assign micromatrizz[5][266] = 9'b111111111;
assign micromatrizz[5][267] = 9'b111111111;
assign micromatrizz[5][268] = 9'b111111111;
assign micromatrizz[5][269] = 9'b111111111;
assign micromatrizz[5][270] = 9'b111111111;
assign micromatrizz[5][271] = 9'b111111111;
assign micromatrizz[5][272] = 9'b111111111;
assign micromatrizz[5][273] = 9'b111111111;
assign micromatrizz[5][274] = 9'b111111111;
assign micromatrizz[5][275] = 9'b111111111;
assign micromatrizz[5][276] = 9'b111111111;
assign micromatrizz[5][277] = 9'b111111111;
assign micromatrizz[5][278] = 9'b111111111;
assign micromatrizz[5][279] = 9'b111111111;
assign micromatrizz[5][280] = 9'b111111111;
assign micromatrizz[5][281] = 9'b111111111;
assign micromatrizz[5][282] = 9'b111111111;
assign micromatrizz[5][283] = 9'b111111111;
assign micromatrizz[5][284] = 9'b111111111;
assign micromatrizz[5][285] = 9'b111111111;
assign micromatrizz[5][286] = 9'b111111111;
assign micromatrizz[5][287] = 9'b111111111;
assign micromatrizz[5][288] = 9'b111111111;
assign micromatrizz[5][289] = 9'b111111111;
assign micromatrizz[5][290] = 9'b111111111;
assign micromatrizz[5][291] = 9'b111111111;
assign micromatrizz[5][292] = 9'b111111111;
assign micromatrizz[5][293] = 9'b111111111;
assign micromatrizz[5][294] = 9'b111111111;
assign micromatrizz[5][295] = 9'b111111111;
assign micromatrizz[5][296] = 9'b111111111;
assign micromatrizz[5][297] = 9'b111111111;
assign micromatrizz[5][298] = 9'b111111111;
assign micromatrizz[5][299] = 9'b111111111;
assign micromatrizz[5][300] = 9'b111111111;
assign micromatrizz[5][301] = 9'b111111111;
assign micromatrizz[5][302] = 9'b111111111;
assign micromatrizz[5][303] = 9'b111111111;
assign micromatrizz[5][304] = 9'b111111111;
assign micromatrizz[5][305] = 9'b111111111;
assign micromatrizz[5][306] = 9'b111111111;
assign micromatrizz[5][307] = 9'b111111111;
assign micromatrizz[5][308] = 9'b111111111;
assign micromatrizz[5][309] = 9'b111111111;
assign micromatrizz[5][310] = 9'b111111111;
assign micromatrizz[5][311] = 9'b111111111;
assign micromatrizz[5][312] = 9'b111111111;
assign micromatrizz[5][313] = 9'b111111111;
assign micromatrizz[5][314] = 9'b111111111;
assign micromatrizz[5][315] = 9'b111111111;
assign micromatrizz[5][316] = 9'b111111111;
assign micromatrizz[5][317] = 9'b111111111;
assign micromatrizz[5][318] = 9'b111111111;
assign micromatrizz[5][319] = 9'b111111111;
assign micromatrizz[5][320] = 9'b111111111;
assign micromatrizz[5][321] = 9'b111111111;
assign micromatrizz[5][322] = 9'b111111111;
assign micromatrizz[5][323] = 9'b111111111;
assign micromatrizz[5][324] = 9'b111111111;
assign micromatrizz[5][325] = 9'b111111111;
assign micromatrizz[5][326] = 9'b111111111;
assign micromatrizz[5][327] = 9'b111111111;
assign micromatrizz[5][328] = 9'b111111111;
assign micromatrizz[5][329] = 9'b111111111;
assign micromatrizz[5][330] = 9'b111111111;
assign micromatrizz[5][331] = 9'b111111111;
assign micromatrizz[5][332] = 9'b111111111;
assign micromatrizz[5][333] = 9'b111111111;
assign micromatrizz[5][334] = 9'b111111111;
assign micromatrizz[5][335] = 9'b111111111;
assign micromatrizz[5][336] = 9'b111111111;
assign micromatrizz[5][337] = 9'b111111111;
assign micromatrizz[5][338] = 9'b111111111;
assign micromatrizz[5][339] = 9'b111111111;
assign micromatrizz[5][340] = 9'b111111111;
assign micromatrizz[5][341] = 9'b111111111;
assign micromatrizz[5][342] = 9'b111111111;
assign micromatrizz[5][343] = 9'b111111111;
assign micromatrizz[5][344] = 9'b111111111;
assign micromatrizz[5][345] = 9'b111111111;
assign micromatrizz[5][346] = 9'b111111111;
assign micromatrizz[5][347] = 9'b111111111;
assign micromatrizz[5][348] = 9'b111111111;
assign micromatrizz[5][349] = 9'b111111111;
assign micromatrizz[5][350] = 9'b111111111;
assign micromatrizz[5][351] = 9'b111111111;
assign micromatrizz[5][352] = 9'b111111111;
assign micromatrizz[5][353] = 9'b111111111;
assign micromatrizz[5][354] = 9'b111111111;
assign micromatrizz[5][355] = 9'b111111111;
assign micromatrizz[5][356] = 9'b111111111;
assign micromatrizz[5][357] = 9'b111111111;
assign micromatrizz[5][358] = 9'b111111111;
assign micromatrizz[5][359] = 9'b111111111;
assign micromatrizz[5][360] = 9'b111111111;
assign micromatrizz[5][361] = 9'b111111111;
assign micromatrizz[5][362] = 9'b111111111;
assign micromatrizz[5][363] = 9'b111111111;
assign micromatrizz[5][364] = 9'b111111111;
assign micromatrizz[5][365] = 9'b111111111;
assign micromatrizz[5][366] = 9'b111111111;
assign micromatrizz[5][367] = 9'b111111111;
assign micromatrizz[5][368] = 9'b111111111;
assign micromatrizz[5][369] = 9'b111111111;
assign micromatrizz[5][370] = 9'b111111111;
assign micromatrizz[5][371] = 9'b111111111;
assign micromatrizz[5][372] = 9'b111111111;
assign micromatrizz[5][373] = 9'b111111111;
assign micromatrizz[5][374] = 9'b111111111;
assign micromatrizz[5][375] = 9'b111111111;
assign micromatrizz[5][376] = 9'b111111111;
assign micromatrizz[5][377] = 9'b111111111;
assign micromatrizz[5][378] = 9'b111111111;
assign micromatrizz[5][379] = 9'b111111111;
assign micromatrizz[5][380] = 9'b111111111;
assign micromatrizz[5][381] = 9'b111111111;
assign micromatrizz[5][382] = 9'b111111111;
assign micromatrizz[5][383] = 9'b111111111;
assign micromatrizz[5][384] = 9'b111111111;
assign micromatrizz[5][385] = 9'b111111111;
assign micromatrizz[5][386] = 9'b111111111;
assign micromatrizz[5][387] = 9'b111111111;
assign micromatrizz[5][388] = 9'b111111111;
assign micromatrizz[5][389] = 9'b111111111;
assign micromatrizz[5][390] = 9'b111111111;
assign micromatrizz[5][391] = 9'b111111111;
assign micromatrizz[5][392] = 9'b111111111;
assign micromatrizz[5][393] = 9'b111111111;
assign micromatrizz[5][394] = 9'b111111111;
assign micromatrizz[5][395] = 9'b111111111;
assign micromatrizz[5][396] = 9'b111111111;
assign micromatrizz[5][397] = 9'b111111111;
assign micromatrizz[5][398] = 9'b111111111;
assign micromatrizz[5][399] = 9'b111111111;
assign micromatrizz[5][400] = 9'b111111111;
assign micromatrizz[5][401] = 9'b111111111;
assign micromatrizz[5][402] = 9'b111111111;
assign micromatrizz[5][403] = 9'b111111111;
assign micromatrizz[5][404] = 9'b111111111;
assign micromatrizz[5][405] = 9'b111111111;
assign micromatrizz[5][406] = 9'b111111111;
assign micromatrizz[5][407] = 9'b111111111;
assign micromatrizz[5][408] = 9'b111111111;
assign micromatrizz[5][409] = 9'b111111111;
assign micromatrizz[5][410] = 9'b111111111;
assign micromatrizz[5][411] = 9'b111111111;
assign micromatrizz[5][412] = 9'b111111111;
assign micromatrizz[5][413] = 9'b111111111;
assign micromatrizz[5][414] = 9'b111111111;
assign micromatrizz[5][415] = 9'b111111111;
assign micromatrizz[5][416] = 9'b111111111;
assign micromatrizz[5][417] = 9'b111111111;
assign micromatrizz[5][418] = 9'b111111111;
assign micromatrizz[5][419] = 9'b111111111;
assign micromatrizz[5][420] = 9'b111111111;
assign micromatrizz[5][421] = 9'b111111111;
assign micromatrizz[5][422] = 9'b111111111;
assign micromatrizz[5][423] = 9'b111111111;
assign micromatrizz[5][424] = 9'b111111111;
assign micromatrizz[5][425] = 9'b111111111;
assign micromatrizz[5][426] = 9'b111111111;
assign micromatrizz[5][427] = 9'b111111111;
assign micromatrizz[5][428] = 9'b111111111;
assign micromatrizz[5][429] = 9'b111111111;
assign micromatrizz[5][430] = 9'b111111111;
assign micromatrizz[5][431] = 9'b111111111;
assign micromatrizz[5][432] = 9'b111111111;
assign micromatrizz[5][433] = 9'b111111111;
assign micromatrizz[5][434] = 9'b111111111;
assign micromatrizz[5][435] = 9'b111111111;
assign micromatrizz[5][436] = 9'b111111111;
assign micromatrizz[5][437] = 9'b111111111;
assign micromatrizz[5][438] = 9'b111111111;
assign micromatrizz[5][439] = 9'b111111111;
assign micromatrizz[5][440] = 9'b111111111;
assign micromatrizz[5][441] = 9'b111111111;
assign micromatrizz[5][442] = 9'b111111111;
assign micromatrizz[5][443] = 9'b111111111;
assign micromatrizz[5][444] = 9'b111111111;
assign micromatrizz[5][445] = 9'b111111111;
assign micromatrizz[5][446] = 9'b111111111;
assign micromatrizz[5][447] = 9'b111111111;
assign micromatrizz[5][448] = 9'b111111111;
assign micromatrizz[5][449] = 9'b111111111;
assign micromatrizz[5][450] = 9'b111111111;
assign micromatrizz[5][451] = 9'b111111111;
assign micromatrizz[5][452] = 9'b111111111;
assign micromatrizz[5][453] = 9'b111111111;
assign micromatrizz[5][454] = 9'b111111111;
assign micromatrizz[5][455] = 9'b111111111;
assign micromatrizz[5][456] = 9'b111111111;
assign micromatrizz[5][457] = 9'b111111111;
assign micromatrizz[5][458] = 9'b111111111;
assign micromatrizz[5][459] = 9'b111111111;
assign micromatrizz[5][460] = 9'b111111111;
assign micromatrizz[5][461] = 9'b111111111;
assign micromatrizz[5][462] = 9'b111111111;
assign micromatrizz[5][463] = 9'b111111111;
assign micromatrizz[5][464] = 9'b111111111;
assign micromatrizz[5][465] = 9'b111111111;
assign micromatrizz[5][466] = 9'b111111111;
assign micromatrizz[5][467] = 9'b111111111;
assign micromatrizz[5][468] = 9'b111111111;
assign micromatrizz[5][469] = 9'b111111111;
assign micromatrizz[5][470] = 9'b111111111;
assign micromatrizz[5][471] = 9'b111111111;
assign micromatrizz[5][472] = 9'b111111111;
assign micromatrizz[5][473] = 9'b111111111;
assign micromatrizz[5][474] = 9'b111111111;
assign micromatrizz[5][475] = 9'b111111111;
assign micromatrizz[5][476] = 9'b111111111;
assign micromatrizz[5][477] = 9'b111111111;
assign micromatrizz[5][478] = 9'b111111111;
assign micromatrizz[5][479] = 9'b111111111;
assign micromatrizz[5][480] = 9'b111111111;
assign micromatrizz[5][481] = 9'b111111111;
assign micromatrizz[5][482] = 9'b111111111;
assign micromatrizz[5][483] = 9'b111111111;
assign micromatrizz[5][484] = 9'b111111111;
assign micromatrizz[5][485] = 9'b111111111;
assign micromatrizz[5][486] = 9'b111111111;
assign micromatrizz[5][487] = 9'b111111111;
assign micromatrizz[5][488] = 9'b111111111;
assign micromatrizz[5][489] = 9'b111111111;
assign micromatrizz[5][490] = 9'b111111111;
assign micromatrizz[5][491] = 9'b111111111;
assign micromatrizz[5][492] = 9'b111111111;
assign micromatrizz[5][493] = 9'b111111111;
assign micromatrizz[5][494] = 9'b111111111;
assign micromatrizz[5][495] = 9'b111111111;
assign micromatrizz[5][496] = 9'b111111111;
assign micromatrizz[5][497] = 9'b111111111;
assign micromatrizz[5][498] = 9'b111111111;
assign micromatrizz[5][499] = 9'b111111111;
assign micromatrizz[5][500] = 9'b111111111;
assign micromatrizz[5][501] = 9'b111111111;
assign micromatrizz[5][502] = 9'b111111111;
assign micromatrizz[5][503] = 9'b111111111;
assign micromatrizz[5][504] = 9'b111111111;
assign micromatrizz[5][505] = 9'b111111111;
assign micromatrizz[5][506] = 9'b111111111;
assign micromatrizz[5][507] = 9'b111111111;
assign micromatrizz[5][508] = 9'b111111111;
assign micromatrizz[5][509] = 9'b111111111;
assign micromatrizz[5][510] = 9'b111111111;
assign micromatrizz[5][511] = 9'b111111111;
assign micromatrizz[5][512] = 9'b111111111;
assign micromatrizz[5][513] = 9'b111111111;
assign micromatrizz[5][514] = 9'b111111111;
assign micromatrizz[5][515] = 9'b111111111;
assign micromatrizz[5][516] = 9'b111111111;
assign micromatrizz[5][517] = 9'b111111111;
assign micromatrizz[5][518] = 9'b111111111;
assign micromatrizz[5][519] = 9'b111111111;
assign micromatrizz[5][520] = 9'b111111111;
assign micromatrizz[5][521] = 9'b111111111;
assign micromatrizz[5][522] = 9'b111111111;
assign micromatrizz[5][523] = 9'b111111111;
assign micromatrizz[5][524] = 9'b111111111;
assign micromatrizz[5][525] = 9'b111111111;
assign micromatrizz[5][526] = 9'b111111111;
assign micromatrizz[5][527] = 9'b111111111;
assign micromatrizz[5][528] = 9'b111111111;
assign micromatrizz[5][529] = 9'b111111111;
assign micromatrizz[5][530] = 9'b111111111;
assign micromatrizz[5][531] = 9'b111111111;
assign micromatrizz[5][532] = 9'b111111111;
assign micromatrizz[5][533] = 9'b111111111;
assign micromatrizz[5][534] = 9'b111111111;
assign micromatrizz[5][535] = 9'b111111111;
assign micromatrizz[5][536] = 9'b111111111;
assign micromatrizz[5][537] = 9'b111111111;
assign micromatrizz[5][538] = 9'b111111111;
assign micromatrizz[5][539] = 9'b111111111;
assign micromatrizz[5][540] = 9'b111111111;
assign micromatrizz[5][541] = 9'b111111111;
assign micromatrizz[5][542] = 9'b111111111;
assign micromatrizz[5][543] = 9'b111111111;
assign micromatrizz[5][544] = 9'b111111111;
assign micromatrizz[5][545] = 9'b111111111;
assign micromatrizz[5][546] = 9'b111111111;
assign micromatrizz[5][547] = 9'b111111111;
assign micromatrizz[5][548] = 9'b111111111;
assign micromatrizz[5][549] = 9'b111111111;
assign micromatrizz[5][550] = 9'b111111111;
assign micromatrizz[5][551] = 9'b111111111;
assign micromatrizz[5][552] = 9'b111111111;
assign micromatrizz[5][553] = 9'b111111111;
assign micromatrizz[5][554] = 9'b111111111;
assign micromatrizz[5][555] = 9'b111111111;
assign micromatrizz[5][556] = 9'b111111111;
assign micromatrizz[5][557] = 9'b111111111;
assign micromatrizz[5][558] = 9'b111111111;
assign micromatrizz[5][559] = 9'b111111111;
assign micromatrizz[5][560] = 9'b111111111;
assign micromatrizz[5][561] = 9'b111111111;
assign micromatrizz[5][562] = 9'b111111111;
assign micromatrizz[5][563] = 9'b111111111;
assign micromatrizz[5][564] = 9'b111111111;
assign micromatrizz[5][565] = 9'b111111111;
assign micromatrizz[5][566] = 9'b111111111;
assign micromatrizz[5][567] = 9'b111111111;
assign micromatrizz[5][568] = 9'b111111111;
assign micromatrizz[5][569] = 9'b111111111;
assign micromatrizz[5][570] = 9'b111111111;
assign micromatrizz[5][571] = 9'b111111111;
assign micromatrizz[5][572] = 9'b111111111;
assign micromatrizz[5][573] = 9'b111111111;
assign micromatrizz[5][574] = 9'b111111111;
assign micromatrizz[5][575] = 9'b111111111;
assign micromatrizz[5][576] = 9'b111111111;
assign micromatrizz[5][577] = 9'b111111111;
assign micromatrizz[5][578] = 9'b111111111;
assign micromatrizz[5][579] = 9'b111111111;
assign micromatrizz[5][580] = 9'b111111111;
assign micromatrizz[5][581] = 9'b111111111;
assign micromatrizz[5][582] = 9'b111111111;
assign micromatrizz[5][583] = 9'b111111111;
assign micromatrizz[5][584] = 9'b111111111;
assign micromatrizz[5][585] = 9'b111111111;
assign micromatrizz[5][586] = 9'b111111111;
assign micromatrizz[5][587] = 9'b111111111;
assign micromatrizz[5][588] = 9'b111111111;
assign micromatrizz[5][589] = 9'b111111111;
assign micromatrizz[5][590] = 9'b111111111;
assign micromatrizz[5][591] = 9'b111111111;
assign micromatrizz[5][592] = 9'b111111111;
assign micromatrizz[5][593] = 9'b111111111;
assign micromatrizz[5][594] = 9'b111111111;
assign micromatrizz[5][595] = 9'b111111111;
assign micromatrizz[5][596] = 9'b111111111;
assign micromatrizz[5][597] = 9'b111111111;
assign micromatrizz[5][598] = 9'b111111111;
assign micromatrizz[5][599] = 9'b111111111;
assign micromatrizz[5][600] = 9'b111111111;
assign micromatrizz[5][601] = 9'b111111111;
assign micromatrizz[5][602] = 9'b111111111;
assign micromatrizz[5][603] = 9'b111111111;
assign micromatrizz[5][604] = 9'b111111111;
assign micromatrizz[5][605] = 9'b111111111;
assign micromatrizz[5][606] = 9'b111111111;
assign micromatrizz[5][607] = 9'b111111111;
assign micromatrizz[5][608] = 9'b111111111;
assign micromatrizz[5][609] = 9'b111111111;
assign micromatrizz[5][610] = 9'b111111111;
assign micromatrizz[5][611] = 9'b111111111;
assign micromatrizz[5][612] = 9'b111111111;
assign micromatrizz[5][613] = 9'b111111111;
assign micromatrizz[5][614] = 9'b111111111;
assign micromatrizz[5][615] = 9'b111111111;
assign micromatrizz[5][616] = 9'b111111111;
assign micromatrizz[5][617] = 9'b111111111;
assign micromatrizz[5][618] = 9'b111111111;
assign micromatrizz[5][619] = 9'b111111111;
assign micromatrizz[5][620] = 9'b111111111;
assign micromatrizz[5][621] = 9'b111111111;
assign micromatrizz[5][622] = 9'b111111111;
assign micromatrizz[5][623] = 9'b111111111;
assign micromatrizz[5][624] = 9'b111111111;
assign micromatrizz[5][625] = 9'b111111111;
assign micromatrizz[5][626] = 9'b111111111;
assign micromatrizz[5][627] = 9'b111111111;
assign micromatrizz[5][628] = 9'b111111111;
assign micromatrizz[5][629] = 9'b111111111;
assign micromatrizz[5][630] = 9'b111111111;
assign micromatrizz[5][631] = 9'b111111111;
assign micromatrizz[5][632] = 9'b111111111;
assign micromatrizz[5][633] = 9'b111111111;
assign micromatrizz[5][634] = 9'b111111111;
assign micromatrizz[5][635] = 9'b111111111;
assign micromatrizz[5][636] = 9'b111111111;
assign micromatrizz[5][637] = 9'b111111111;
assign micromatrizz[5][638] = 9'b111111111;
assign micromatrizz[5][639] = 9'b111111111;
assign micromatrizz[6][0] = 9'b111111111;
assign micromatrizz[6][1] = 9'b111111111;
assign micromatrizz[6][2] = 9'b111111111;
assign micromatrizz[6][3] = 9'b111111111;
assign micromatrizz[6][4] = 9'b111111111;
assign micromatrizz[6][5] = 9'b111111111;
assign micromatrizz[6][6] = 9'b111111111;
assign micromatrizz[6][7] = 9'b111111111;
assign micromatrizz[6][8] = 9'b111111111;
assign micromatrizz[6][9] = 9'b111111111;
assign micromatrizz[6][10] = 9'b111111111;
assign micromatrizz[6][11] = 9'b111111111;
assign micromatrizz[6][12] = 9'b111111111;
assign micromatrizz[6][13] = 9'b111111111;
assign micromatrizz[6][14] = 9'b111111111;
assign micromatrizz[6][15] = 9'b111111111;
assign micromatrizz[6][16] = 9'b111111111;
assign micromatrizz[6][17] = 9'b111111111;
assign micromatrizz[6][18] = 9'b111111111;
assign micromatrizz[6][19] = 9'b111111111;
assign micromatrizz[6][20] = 9'b111111111;
assign micromatrizz[6][21] = 9'b111111111;
assign micromatrizz[6][22] = 9'b111111111;
assign micromatrizz[6][23] = 9'b111111111;
assign micromatrizz[6][24] = 9'b111111111;
assign micromatrizz[6][25] = 9'b111111111;
assign micromatrizz[6][26] = 9'b111111111;
assign micromatrizz[6][27] = 9'b111111111;
assign micromatrizz[6][28] = 9'b111111111;
assign micromatrizz[6][29] = 9'b111111111;
assign micromatrizz[6][30] = 9'b111111111;
assign micromatrizz[6][31] = 9'b111111111;
assign micromatrizz[6][32] = 9'b111111111;
assign micromatrizz[6][33] = 9'b111111111;
assign micromatrizz[6][34] = 9'b111111111;
assign micromatrizz[6][35] = 9'b111111111;
assign micromatrizz[6][36] = 9'b111111111;
assign micromatrizz[6][37] = 9'b111111111;
assign micromatrizz[6][38] = 9'b111111111;
assign micromatrizz[6][39] = 9'b111111111;
assign micromatrizz[6][40] = 9'b111111111;
assign micromatrizz[6][41] = 9'b111111111;
assign micromatrizz[6][42] = 9'b111111111;
assign micromatrizz[6][43] = 9'b111111111;
assign micromatrizz[6][44] = 9'b111111111;
assign micromatrizz[6][45] = 9'b111111111;
assign micromatrizz[6][46] = 9'b111111111;
assign micromatrizz[6][47] = 9'b111111111;
assign micromatrizz[6][48] = 9'b111111111;
assign micromatrizz[6][49] = 9'b111111111;
assign micromatrizz[6][50] = 9'b111111111;
assign micromatrizz[6][51] = 9'b111111111;
assign micromatrizz[6][52] = 9'b111111111;
assign micromatrizz[6][53] = 9'b111111111;
assign micromatrizz[6][54] = 9'b111111111;
assign micromatrizz[6][55] = 9'b111111111;
assign micromatrizz[6][56] = 9'b111111111;
assign micromatrizz[6][57] = 9'b111111111;
assign micromatrizz[6][58] = 9'b111111111;
assign micromatrizz[6][59] = 9'b111111111;
assign micromatrizz[6][60] = 9'b111111111;
assign micromatrizz[6][61] = 9'b111111111;
assign micromatrizz[6][62] = 9'b111111111;
assign micromatrizz[6][63] = 9'b111111111;
assign micromatrizz[6][64] = 9'b111111111;
assign micromatrizz[6][65] = 9'b111111111;
assign micromatrizz[6][66] = 9'b111111111;
assign micromatrizz[6][67] = 9'b111111111;
assign micromatrizz[6][68] = 9'b111111111;
assign micromatrizz[6][69] = 9'b111111111;
assign micromatrizz[6][70] = 9'b111111111;
assign micromatrizz[6][71] = 9'b111111111;
assign micromatrizz[6][72] = 9'b111111111;
assign micromatrizz[6][73] = 9'b111111111;
assign micromatrizz[6][74] = 9'b111111111;
assign micromatrizz[6][75] = 9'b111111111;
assign micromatrizz[6][76] = 9'b111111111;
assign micromatrizz[6][77] = 9'b111111111;
assign micromatrizz[6][78] = 9'b111111111;
assign micromatrizz[6][79] = 9'b111111111;
assign micromatrizz[6][80] = 9'b111111111;
assign micromatrizz[6][81] = 9'b111111111;
assign micromatrizz[6][82] = 9'b111111111;
assign micromatrizz[6][83] = 9'b111111111;
assign micromatrizz[6][84] = 9'b111111111;
assign micromatrizz[6][85] = 9'b111111111;
assign micromatrizz[6][86] = 9'b111111111;
assign micromatrizz[6][87] = 9'b111111111;
assign micromatrizz[6][88] = 9'b111111111;
assign micromatrizz[6][89] = 9'b111111111;
assign micromatrizz[6][90] = 9'b111111111;
assign micromatrizz[6][91] = 9'b111111111;
assign micromatrizz[6][92] = 9'b111111111;
assign micromatrizz[6][93] = 9'b111111111;
assign micromatrizz[6][94] = 9'b111111111;
assign micromatrizz[6][95] = 9'b111111111;
assign micromatrizz[6][96] = 9'b111111111;
assign micromatrizz[6][97] = 9'b111111111;
assign micromatrizz[6][98] = 9'b111111111;
assign micromatrizz[6][99] = 9'b111111111;
assign micromatrizz[6][100] = 9'b111111111;
assign micromatrizz[6][101] = 9'b111111111;
assign micromatrizz[6][102] = 9'b111111111;
assign micromatrizz[6][103] = 9'b111111111;
assign micromatrizz[6][104] = 9'b111111111;
assign micromatrizz[6][105] = 9'b111111111;
assign micromatrizz[6][106] = 9'b111111111;
assign micromatrizz[6][107] = 9'b111111111;
assign micromatrizz[6][108] = 9'b111111111;
assign micromatrizz[6][109] = 9'b111111111;
assign micromatrizz[6][110] = 9'b111111111;
assign micromatrizz[6][111] = 9'b111111111;
assign micromatrizz[6][112] = 9'b111111111;
assign micromatrizz[6][113] = 9'b111111111;
assign micromatrizz[6][114] = 9'b111111111;
assign micromatrizz[6][115] = 9'b111111111;
assign micromatrizz[6][116] = 9'b111111111;
assign micromatrizz[6][117] = 9'b111111111;
assign micromatrizz[6][118] = 9'b111111111;
assign micromatrizz[6][119] = 9'b111111111;
assign micromatrizz[6][120] = 9'b111111111;
assign micromatrizz[6][121] = 9'b111111111;
assign micromatrizz[6][122] = 9'b111111111;
assign micromatrizz[6][123] = 9'b111111111;
assign micromatrizz[6][124] = 9'b111111111;
assign micromatrizz[6][125] = 9'b111111111;
assign micromatrizz[6][126] = 9'b111111111;
assign micromatrizz[6][127] = 9'b111111111;
assign micromatrizz[6][128] = 9'b111111111;
assign micromatrizz[6][129] = 9'b111111111;
assign micromatrizz[6][130] = 9'b111111111;
assign micromatrizz[6][131] = 9'b111111111;
assign micromatrizz[6][132] = 9'b111111111;
assign micromatrizz[6][133] = 9'b111111111;
assign micromatrizz[6][134] = 9'b111111111;
assign micromatrizz[6][135] = 9'b111111111;
assign micromatrizz[6][136] = 9'b111111111;
assign micromatrizz[6][137] = 9'b111111111;
assign micromatrizz[6][138] = 9'b111111111;
assign micromatrizz[6][139] = 9'b111111111;
assign micromatrizz[6][140] = 9'b111111111;
assign micromatrizz[6][141] = 9'b111111111;
assign micromatrizz[6][142] = 9'b111111111;
assign micromatrizz[6][143] = 9'b111111111;
assign micromatrizz[6][144] = 9'b111111111;
assign micromatrizz[6][145] = 9'b111111111;
assign micromatrizz[6][146] = 9'b111111111;
assign micromatrizz[6][147] = 9'b111111111;
assign micromatrizz[6][148] = 9'b111111111;
assign micromatrizz[6][149] = 9'b111111111;
assign micromatrizz[6][150] = 9'b111111111;
assign micromatrizz[6][151] = 9'b111111111;
assign micromatrizz[6][152] = 9'b111111111;
assign micromatrizz[6][153] = 9'b111111111;
assign micromatrizz[6][154] = 9'b111111111;
assign micromatrizz[6][155] = 9'b111111111;
assign micromatrizz[6][156] = 9'b111111111;
assign micromatrizz[6][157] = 9'b111111111;
assign micromatrizz[6][158] = 9'b111111111;
assign micromatrizz[6][159] = 9'b111111111;
assign micromatrizz[6][160] = 9'b111111111;
assign micromatrizz[6][161] = 9'b111111111;
assign micromatrizz[6][162] = 9'b111111111;
assign micromatrizz[6][163] = 9'b111111111;
assign micromatrizz[6][164] = 9'b111111111;
assign micromatrizz[6][165] = 9'b111111111;
assign micromatrizz[6][166] = 9'b111111111;
assign micromatrizz[6][167] = 9'b111111111;
assign micromatrizz[6][168] = 9'b111111111;
assign micromatrizz[6][169] = 9'b111111111;
assign micromatrizz[6][170] = 9'b111111111;
assign micromatrizz[6][171] = 9'b111111111;
assign micromatrizz[6][172] = 9'b111111111;
assign micromatrizz[6][173] = 9'b111111111;
assign micromatrizz[6][174] = 9'b111111111;
assign micromatrizz[6][175] = 9'b111111111;
assign micromatrizz[6][176] = 9'b111111111;
assign micromatrizz[6][177] = 9'b111111111;
assign micromatrizz[6][178] = 9'b111111111;
assign micromatrizz[6][179] = 9'b111111111;
assign micromatrizz[6][180] = 9'b111111111;
assign micromatrizz[6][181] = 9'b111111111;
assign micromatrizz[6][182] = 9'b111111111;
assign micromatrizz[6][183] = 9'b111111111;
assign micromatrizz[6][184] = 9'b111111111;
assign micromatrizz[6][185] = 9'b111111111;
assign micromatrizz[6][186] = 9'b111111111;
assign micromatrizz[6][187] = 9'b111111111;
assign micromatrizz[6][188] = 9'b111111111;
assign micromatrizz[6][189] = 9'b111111111;
assign micromatrizz[6][190] = 9'b111111111;
assign micromatrizz[6][191] = 9'b111111111;
assign micromatrizz[6][192] = 9'b111111111;
assign micromatrizz[6][193] = 9'b111111111;
assign micromatrizz[6][194] = 9'b111111111;
assign micromatrizz[6][195] = 9'b111111111;
assign micromatrizz[6][196] = 9'b111111111;
assign micromatrizz[6][197] = 9'b111111111;
assign micromatrizz[6][198] = 9'b111111111;
assign micromatrizz[6][199] = 9'b111111111;
assign micromatrizz[6][200] = 9'b111111111;
assign micromatrizz[6][201] = 9'b111111111;
assign micromatrizz[6][202] = 9'b111111111;
assign micromatrizz[6][203] = 9'b111111111;
assign micromatrizz[6][204] = 9'b111111111;
assign micromatrizz[6][205] = 9'b111111111;
assign micromatrizz[6][206] = 9'b111111111;
assign micromatrizz[6][207] = 9'b111111111;
assign micromatrizz[6][208] = 9'b111111111;
assign micromatrizz[6][209] = 9'b111111111;
assign micromatrizz[6][210] = 9'b111111111;
assign micromatrizz[6][211] = 9'b111111111;
assign micromatrizz[6][212] = 9'b111111111;
assign micromatrizz[6][213] = 9'b111111111;
assign micromatrizz[6][214] = 9'b111111111;
assign micromatrizz[6][215] = 9'b111111111;
assign micromatrizz[6][216] = 9'b111111111;
assign micromatrizz[6][217] = 9'b111111111;
assign micromatrizz[6][218] = 9'b111111111;
assign micromatrizz[6][219] = 9'b111111111;
assign micromatrizz[6][220] = 9'b111111111;
assign micromatrizz[6][221] = 9'b111111111;
assign micromatrizz[6][222] = 9'b111111111;
assign micromatrizz[6][223] = 9'b111111111;
assign micromatrizz[6][224] = 9'b111111111;
assign micromatrizz[6][225] = 9'b111111111;
assign micromatrizz[6][226] = 9'b111111111;
assign micromatrizz[6][227] = 9'b111111111;
assign micromatrizz[6][228] = 9'b111111111;
assign micromatrizz[6][229] = 9'b111111111;
assign micromatrizz[6][230] = 9'b111111111;
assign micromatrizz[6][231] = 9'b111111111;
assign micromatrizz[6][232] = 9'b111111111;
assign micromatrizz[6][233] = 9'b111111111;
assign micromatrizz[6][234] = 9'b111111111;
assign micromatrizz[6][235] = 9'b111111111;
assign micromatrizz[6][236] = 9'b111111111;
assign micromatrizz[6][237] = 9'b111111111;
assign micromatrizz[6][238] = 9'b111111111;
assign micromatrizz[6][239] = 9'b111111111;
assign micromatrizz[6][240] = 9'b111111111;
assign micromatrizz[6][241] = 9'b111111111;
assign micromatrizz[6][242] = 9'b111111111;
assign micromatrizz[6][243] = 9'b111111111;
assign micromatrizz[6][244] = 9'b111111111;
assign micromatrizz[6][245] = 9'b111111111;
assign micromatrizz[6][246] = 9'b111111111;
assign micromatrizz[6][247] = 9'b111111111;
assign micromatrizz[6][248] = 9'b111111111;
assign micromatrizz[6][249] = 9'b111111111;
assign micromatrizz[6][250] = 9'b111111111;
assign micromatrizz[6][251] = 9'b111111111;
assign micromatrizz[6][252] = 9'b111111111;
assign micromatrizz[6][253] = 9'b111111111;
assign micromatrizz[6][254] = 9'b111111111;
assign micromatrizz[6][255] = 9'b111111111;
assign micromatrizz[6][256] = 9'b111111111;
assign micromatrizz[6][257] = 9'b111111111;
assign micromatrizz[6][258] = 9'b111111111;
assign micromatrizz[6][259] = 9'b111111111;
assign micromatrizz[6][260] = 9'b111111111;
assign micromatrizz[6][261] = 9'b111111111;
assign micromatrizz[6][262] = 9'b111111111;
assign micromatrizz[6][263] = 9'b111111111;
assign micromatrizz[6][264] = 9'b111111111;
assign micromatrizz[6][265] = 9'b111111111;
assign micromatrizz[6][266] = 9'b111111111;
assign micromatrizz[6][267] = 9'b111111111;
assign micromatrizz[6][268] = 9'b111111111;
assign micromatrizz[6][269] = 9'b111111111;
assign micromatrizz[6][270] = 9'b111111111;
assign micromatrizz[6][271] = 9'b111111111;
assign micromatrizz[6][272] = 9'b111111111;
assign micromatrizz[6][273] = 9'b111111111;
assign micromatrizz[6][274] = 9'b111111111;
assign micromatrizz[6][275] = 9'b111111111;
assign micromatrizz[6][276] = 9'b111111111;
assign micromatrizz[6][277] = 9'b111111111;
assign micromatrizz[6][278] = 9'b111111111;
assign micromatrizz[6][279] = 9'b111111111;
assign micromatrizz[6][280] = 9'b111111111;
assign micromatrizz[6][281] = 9'b111111111;
assign micromatrizz[6][282] = 9'b111111111;
assign micromatrizz[6][283] = 9'b111111111;
assign micromatrizz[6][284] = 9'b111111111;
assign micromatrizz[6][285] = 9'b111111111;
assign micromatrizz[6][286] = 9'b111111111;
assign micromatrizz[6][287] = 9'b111111111;
assign micromatrizz[6][288] = 9'b111111111;
assign micromatrizz[6][289] = 9'b111111111;
assign micromatrizz[6][290] = 9'b111111111;
assign micromatrizz[6][291] = 9'b111111111;
assign micromatrizz[6][292] = 9'b111111111;
assign micromatrizz[6][293] = 9'b111111111;
assign micromatrizz[6][294] = 9'b111111111;
assign micromatrizz[6][295] = 9'b111111111;
assign micromatrizz[6][296] = 9'b111111111;
assign micromatrizz[6][297] = 9'b111111111;
assign micromatrizz[6][298] = 9'b111111111;
assign micromatrizz[6][299] = 9'b111111111;
assign micromatrizz[6][300] = 9'b111111111;
assign micromatrizz[6][301] = 9'b111111111;
assign micromatrizz[6][302] = 9'b111111111;
assign micromatrizz[6][303] = 9'b111111111;
assign micromatrizz[6][304] = 9'b111111111;
assign micromatrizz[6][305] = 9'b111111111;
assign micromatrizz[6][306] = 9'b111111111;
assign micromatrizz[6][307] = 9'b111111111;
assign micromatrizz[6][308] = 9'b111111111;
assign micromatrizz[6][309] = 9'b111111111;
assign micromatrizz[6][310] = 9'b111111111;
assign micromatrizz[6][311] = 9'b111111111;
assign micromatrizz[6][312] = 9'b111111111;
assign micromatrizz[6][313] = 9'b111111111;
assign micromatrizz[6][314] = 9'b111111111;
assign micromatrizz[6][315] = 9'b111111111;
assign micromatrizz[6][316] = 9'b111111111;
assign micromatrizz[6][317] = 9'b111111111;
assign micromatrizz[6][318] = 9'b111111111;
assign micromatrizz[6][319] = 9'b111111111;
assign micromatrizz[6][320] = 9'b111111111;
assign micromatrizz[6][321] = 9'b111111111;
assign micromatrizz[6][322] = 9'b111111111;
assign micromatrizz[6][323] = 9'b111111111;
assign micromatrizz[6][324] = 9'b111111111;
assign micromatrizz[6][325] = 9'b111111111;
assign micromatrizz[6][326] = 9'b111111111;
assign micromatrizz[6][327] = 9'b111111111;
assign micromatrizz[6][328] = 9'b111111111;
assign micromatrizz[6][329] = 9'b111111111;
assign micromatrizz[6][330] = 9'b111111111;
assign micromatrizz[6][331] = 9'b111111111;
assign micromatrizz[6][332] = 9'b111111111;
assign micromatrizz[6][333] = 9'b111111111;
assign micromatrizz[6][334] = 9'b111111111;
assign micromatrizz[6][335] = 9'b111111111;
assign micromatrizz[6][336] = 9'b111111111;
assign micromatrizz[6][337] = 9'b111111111;
assign micromatrizz[6][338] = 9'b111111111;
assign micromatrizz[6][339] = 9'b111111111;
assign micromatrizz[6][340] = 9'b111111111;
assign micromatrizz[6][341] = 9'b111111111;
assign micromatrizz[6][342] = 9'b111111111;
assign micromatrizz[6][343] = 9'b111111111;
assign micromatrizz[6][344] = 9'b111111111;
assign micromatrizz[6][345] = 9'b111111111;
assign micromatrizz[6][346] = 9'b111111111;
assign micromatrizz[6][347] = 9'b111111111;
assign micromatrizz[6][348] = 9'b111111111;
assign micromatrizz[6][349] = 9'b111111111;
assign micromatrizz[6][350] = 9'b111111111;
assign micromatrizz[6][351] = 9'b111111111;
assign micromatrizz[6][352] = 9'b111111111;
assign micromatrizz[6][353] = 9'b111111111;
assign micromatrizz[6][354] = 9'b111111111;
assign micromatrizz[6][355] = 9'b111111111;
assign micromatrizz[6][356] = 9'b111111111;
assign micromatrizz[6][357] = 9'b111111111;
assign micromatrizz[6][358] = 9'b111111111;
assign micromatrizz[6][359] = 9'b111111111;
assign micromatrizz[6][360] = 9'b111111111;
assign micromatrizz[6][361] = 9'b111111111;
assign micromatrizz[6][362] = 9'b111111111;
assign micromatrizz[6][363] = 9'b111111111;
assign micromatrizz[6][364] = 9'b111111111;
assign micromatrizz[6][365] = 9'b111111111;
assign micromatrizz[6][366] = 9'b111111111;
assign micromatrizz[6][367] = 9'b111111111;
assign micromatrizz[6][368] = 9'b111111111;
assign micromatrizz[6][369] = 9'b111111111;
assign micromatrizz[6][370] = 9'b111111111;
assign micromatrizz[6][371] = 9'b111111111;
assign micromatrizz[6][372] = 9'b111111111;
assign micromatrizz[6][373] = 9'b111111111;
assign micromatrizz[6][374] = 9'b111111111;
assign micromatrizz[6][375] = 9'b111111111;
assign micromatrizz[6][376] = 9'b111111111;
assign micromatrizz[6][377] = 9'b111111111;
assign micromatrizz[6][378] = 9'b111111111;
assign micromatrizz[6][379] = 9'b111111111;
assign micromatrizz[6][380] = 9'b111111111;
assign micromatrizz[6][381] = 9'b111111111;
assign micromatrizz[6][382] = 9'b111111111;
assign micromatrizz[6][383] = 9'b111111111;
assign micromatrizz[6][384] = 9'b111111111;
assign micromatrizz[6][385] = 9'b111111111;
assign micromatrizz[6][386] = 9'b111111111;
assign micromatrizz[6][387] = 9'b111111111;
assign micromatrizz[6][388] = 9'b111111111;
assign micromatrizz[6][389] = 9'b111111111;
assign micromatrizz[6][390] = 9'b111111111;
assign micromatrizz[6][391] = 9'b111111111;
assign micromatrizz[6][392] = 9'b111111111;
assign micromatrizz[6][393] = 9'b111111111;
assign micromatrizz[6][394] = 9'b111111111;
assign micromatrizz[6][395] = 9'b111111111;
assign micromatrizz[6][396] = 9'b111111111;
assign micromatrizz[6][397] = 9'b111111111;
assign micromatrizz[6][398] = 9'b111111111;
assign micromatrizz[6][399] = 9'b111111111;
assign micromatrizz[6][400] = 9'b111111111;
assign micromatrizz[6][401] = 9'b111111111;
assign micromatrizz[6][402] = 9'b111111111;
assign micromatrizz[6][403] = 9'b111111111;
assign micromatrizz[6][404] = 9'b111111111;
assign micromatrizz[6][405] = 9'b111111111;
assign micromatrizz[6][406] = 9'b111111111;
assign micromatrizz[6][407] = 9'b111111111;
assign micromatrizz[6][408] = 9'b111111111;
assign micromatrizz[6][409] = 9'b111111111;
assign micromatrizz[6][410] = 9'b111111111;
assign micromatrizz[6][411] = 9'b111111111;
assign micromatrizz[6][412] = 9'b111111111;
assign micromatrizz[6][413] = 9'b111111111;
assign micromatrizz[6][414] = 9'b111111111;
assign micromatrizz[6][415] = 9'b111111111;
assign micromatrizz[6][416] = 9'b111111111;
assign micromatrizz[6][417] = 9'b111111111;
assign micromatrizz[6][418] = 9'b111111111;
assign micromatrizz[6][419] = 9'b111111111;
assign micromatrizz[6][420] = 9'b111111111;
assign micromatrizz[6][421] = 9'b111111111;
assign micromatrizz[6][422] = 9'b111111111;
assign micromatrizz[6][423] = 9'b111111111;
assign micromatrizz[6][424] = 9'b111111111;
assign micromatrizz[6][425] = 9'b111111111;
assign micromatrizz[6][426] = 9'b111111111;
assign micromatrizz[6][427] = 9'b111111111;
assign micromatrizz[6][428] = 9'b111111111;
assign micromatrizz[6][429] = 9'b111111111;
assign micromatrizz[6][430] = 9'b111111111;
assign micromatrizz[6][431] = 9'b111111111;
assign micromatrizz[6][432] = 9'b111111111;
assign micromatrizz[6][433] = 9'b111111111;
assign micromatrizz[6][434] = 9'b111111111;
assign micromatrizz[6][435] = 9'b111111111;
assign micromatrizz[6][436] = 9'b111111111;
assign micromatrizz[6][437] = 9'b111111111;
assign micromatrizz[6][438] = 9'b111111111;
assign micromatrizz[6][439] = 9'b111111111;
assign micromatrizz[6][440] = 9'b111111111;
assign micromatrizz[6][441] = 9'b111111111;
assign micromatrizz[6][442] = 9'b111111111;
assign micromatrizz[6][443] = 9'b111111111;
assign micromatrizz[6][444] = 9'b111111111;
assign micromatrizz[6][445] = 9'b111111111;
assign micromatrizz[6][446] = 9'b111111111;
assign micromatrizz[6][447] = 9'b111111111;
assign micromatrizz[6][448] = 9'b111111111;
assign micromatrizz[6][449] = 9'b111111111;
assign micromatrizz[6][450] = 9'b111111111;
assign micromatrizz[6][451] = 9'b111111111;
assign micromatrizz[6][452] = 9'b111111111;
assign micromatrizz[6][453] = 9'b111111111;
assign micromatrizz[6][454] = 9'b111111111;
assign micromatrizz[6][455] = 9'b111111111;
assign micromatrizz[6][456] = 9'b111111111;
assign micromatrizz[6][457] = 9'b111111111;
assign micromatrizz[6][458] = 9'b111111111;
assign micromatrizz[6][459] = 9'b111111111;
assign micromatrizz[6][460] = 9'b111111111;
assign micromatrizz[6][461] = 9'b111111111;
assign micromatrizz[6][462] = 9'b111111111;
assign micromatrizz[6][463] = 9'b111111111;
assign micromatrizz[6][464] = 9'b111111111;
assign micromatrizz[6][465] = 9'b111111111;
assign micromatrizz[6][466] = 9'b111111111;
assign micromatrizz[6][467] = 9'b111111111;
assign micromatrizz[6][468] = 9'b111111111;
assign micromatrizz[6][469] = 9'b111111111;
assign micromatrizz[6][470] = 9'b111111111;
assign micromatrizz[6][471] = 9'b111111111;
assign micromatrizz[6][472] = 9'b111111111;
assign micromatrizz[6][473] = 9'b111111111;
assign micromatrizz[6][474] = 9'b111111111;
assign micromatrizz[6][475] = 9'b111111111;
assign micromatrizz[6][476] = 9'b111111111;
assign micromatrizz[6][477] = 9'b111111111;
assign micromatrizz[6][478] = 9'b111111111;
assign micromatrizz[6][479] = 9'b111111111;
assign micromatrizz[6][480] = 9'b111111111;
assign micromatrizz[6][481] = 9'b111111111;
assign micromatrizz[6][482] = 9'b111111111;
assign micromatrizz[6][483] = 9'b111111111;
assign micromatrizz[6][484] = 9'b111111111;
assign micromatrizz[6][485] = 9'b111111111;
assign micromatrizz[6][486] = 9'b111111111;
assign micromatrizz[6][487] = 9'b111111111;
assign micromatrizz[6][488] = 9'b111111111;
assign micromatrizz[6][489] = 9'b111111111;
assign micromatrizz[6][490] = 9'b111111111;
assign micromatrizz[6][491] = 9'b111111111;
assign micromatrizz[6][492] = 9'b111111111;
assign micromatrizz[6][493] = 9'b111111111;
assign micromatrizz[6][494] = 9'b111111111;
assign micromatrizz[6][495] = 9'b111111111;
assign micromatrizz[6][496] = 9'b111111111;
assign micromatrizz[6][497] = 9'b111111111;
assign micromatrizz[6][498] = 9'b111111111;
assign micromatrizz[6][499] = 9'b111111111;
assign micromatrizz[6][500] = 9'b111111111;
assign micromatrizz[6][501] = 9'b111111111;
assign micromatrizz[6][502] = 9'b111111111;
assign micromatrizz[6][503] = 9'b111111111;
assign micromatrizz[6][504] = 9'b111111111;
assign micromatrizz[6][505] = 9'b111111111;
assign micromatrizz[6][506] = 9'b111111111;
assign micromatrizz[6][507] = 9'b111111111;
assign micromatrizz[6][508] = 9'b111111111;
assign micromatrizz[6][509] = 9'b111111111;
assign micromatrizz[6][510] = 9'b111111111;
assign micromatrizz[6][511] = 9'b111111111;
assign micromatrizz[6][512] = 9'b111111111;
assign micromatrizz[6][513] = 9'b111111111;
assign micromatrizz[6][514] = 9'b111111111;
assign micromatrizz[6][515] = 9'b111111111;
assign micromatrizz[6][516] = 9'b111111111;
assign micromatrizz[6][517] = 9'b111111111;
assign micromatrizz[6][518] = 9'b111111111;
assign micromatrizz[6][519] = 9'b111111111;
assign micromatrizz[6][520] = 9'b111111111;
assign micromatrizz[6][521] = 9'b111111111;
assign micromatrizz[6][522] = 9'b111111111;
assign micromatrizz[6][523] = 9'b111111111;
assign micromatrizz[6][524] = 9'b111111111;
assign micromatrizz[6][525] = 9'b111111111;
assign micromatrizz[6][526] = 9'b111111111;
assign micromatrizz[6][527] = 9'b111111111;
assign micromatrizz[6][528] = 9'b111111111;
assign micromatrizz[6][529] = 9'b111111111;
assign micromatrizz[6][530] = 9'b111111111;
assign micromatrizz[6][531] = 9'b111111111;
assign micromatrizz[6][532] = 9'b111111111;
assign micromatrizz[6][533] = 9'b111111111;
assign micromatrizz[6][534] = 9'b111111111;
assign micromatrizz[6][535] = 9'b111111111;
assign micromatrizz[6][536] = 9'b111111111;
assign micromatrizz[6][537] = 9'b111111111;
assign micromatrizz[6][538] = 9'b111111111;
assign micromatrizz[6][539] = 9'b111111111;
assign micromatrizz[6][540] = 9'b111111111;
assign micromatrizz[6][541] = 9'b111111111;
assign micromatrizz[6][542] = 9'b111111111;
assign micromatrizz[6][543] = 9'b111111111;
assign micromatrizz[6][544] = 9'b111111111;
assign micromatrizz[6][545] = 9'b111111111;
assign micromatrizz[6][546] = 9'b111111111;
assign micromatrizz[6][547] = 9'b111111111;
assign micromatrizz[6][548] = 9'b111111111;
assign micromatrizz[6][549] = 9'b111111111;
assign micromatrizz[6][550] = 9'b111111111;
assign micromatrizz[6][551] = 9'b111111111;
assign micromatrizz[6][552] = 9'b111111111;
assign micromatrizz[6][553] = 9'b111111111;
assign micromatrizz[6][554] = 9'b111111111;
assign micromatrizz[6][555] = 9'b111111111;
assign micromatrizz[6][556] = 9'b111111111;
assign micromatrizz[6][557] = 9'b111111111;
assign micromatrizz[6][558] = 9'b111111111;
assign micromatrizz[6][559] = 9'b111111111;
assign micromatrizz[6][560] = 9'b111111111;
assign micromatrizz[6][561] = 9'b111111111;
assign micromatrizz[6][562] = 9'b111111111;
assign micromatrizz[6][563] = 9'b111111111;
assign micromatrizz[6][564] = 9'b111111111;
assign micromatrizz[6][565] = 9'b111111111;
assign micromatrizz[6][566] = 9'b111111111;
assign micromatrizz[6][567] = 9'b111111111;
assign micromatrizz[6][568] = 9'b111111111;
assign micromatrizz[6][569] = 9'b111111111;
assign micromatrizz[6][570] = 9'b111111111;
assign micromatrizz[6][571] = 9'b111111111;
assign micromatrizz[6][572] = 9'b111111111;
assign micromatrizz[6][573] = 9'b111111111;
assign micromatrizz[6][574] = 9'b111111111;
assign micromatrizz[6][575] = 9'b111111111;
assign micromatrizz[6][576] = 9'b111111111;
assign micromatrizz[6][577] = 9'b111111111;
assign micromatrizz[6][578] = 9'b111111111;
assign micromatrizz[6][579] = 9'b111111111;
assign micromatrizz[6][580] = 9'b111111111;
assign micromatrizz[6][581] = 9'b111111111;
assign micromatrizz[6][582] = 9'b111111111;
assign micromatrizz[6][583] = 9'b111111111;
assign micromatrizz[6][584] = 9'b111111111;
assign micromatrizz[6][585] = 9'b111111111;
assign micromatrizz[6][586] = 9'b111111111;
assign micromatrizz[6][587] = 9'b111111111;
assign micromatrizz[6][588] = 9'b111111111;
assign micromatrizz[6][589] = 9'b111111111;
assign micromatrizz[6][590] = 9'b111111111;
assign micromatrizz[6][591] = 9'b111111111;
assign micromatrizz[6][592] = 9'b111111111;
assign micromatrizz[6][593] = 9'b111111111;
assign micromatrizz[6][594] = 9'b111111111;
assign micromatrizz[6][595] = 9'b111111111;
assign micromatrizz[6][596] = 9'b111111111;
assign micromatrizz[6][597] = 9'b111111111;
assign micromatrizz[6][598] = 9'b111111111;
assign micromatrizz[6][599] = 9'b111111111;
assign micromatrizz[6][600] = 9'b111111111;
assign micromatrizz[6][601] = 9'b111111111;
assign micromatrizz[6][602] = 9'b111111111;
assign micromatrizz[6][603] = 9'b111111111;
assign micromatrizz[6][604] = 9'b111111111;
assign micromatrizz[6][605] = 9'b111111111;
assign micromatrizz[6][606] = 9'b111111111;
assign micromatrizz[6][607] = 9'b111111111;
assign micromatrizz[6][608] = 9'b111111111;
assign micromatrizz[6][609] = 9'b111111111;
assign micromatrizz[6][610] = 9'b111111111;
assign micromatrizz[6][611] = 9'b111111111;
assign micromatrizz[6][612] = 9'b111111111;
assign micromatrizz[6][613] = 9'b111111111;
assign micromatrizz[6][614] = 9'b111111111;
assign micromatrizz[6][615] = 9'b111111111;
assign micromatrizz[6][616] = 9'b111111111;
assign micromatrizz[6][617] = 9'b111111111;
assign micromatrizz[6][618] = 9'b111111111;
assign micromatrizz[6][619] = 9'b111111111;
assign micromatrizz[6][620] = 9'b111111111;
assign micromatrizz[6][621] = 9'b111111111;
assign micromatrizz[6][622] = 9'b111111111;
assign micromatrizz[6][623] = 9'b111111111;
assign micromatrizz[6][624] = 9'b111111111;
assign micromatrizz[6][625] = 9'b111111111;
assign micromatrizz[6][626] = 9'b111111111;
assign micromatrizz[6][627] = 9'b111111111;
assign micromatrizz[6][628] = 9'b111111111;
assign micromatrizz[6][629] = 9'b111111111;
assign micromatrizz[6][630] = 9'b111111111;
assign micromatrizz[6][631] = 9'b111111111;
assign micromatrizz[6][632] = 9'b111111111;
assign micromatrizz[6][633] = 9'b111111111;
assign micromatrizz[6][634] = 9'b111111111;
assign micromatrizz[6][635] = 9'b111111111;
assign micromatrizz[6][636] = 9'b111111111;
assign micromatrizz[6][637] = 9'b111111111;
assign micromatrizz[6][638] = 9'b111111111;
assign micromatrizz[6][639] = 9'b111111111;
assign micromatrizz[7][0] = 9'b111111111;
assign micromatrizz[7][1] = 9'b111111111;
assign micromatrizz[7][2] = 9'b111111111;
assign micromatrizz[7][3] = 9'b111111111;
assign micromatrizz[7][4] = 9'b111111111;
assign micromatrizz[7][5] = 9'b111111111;
assign micromatrizz[7][6] = 9'b111111111;
assign micromatrizz[7][7] = 9'b111111111;
assign micromatrizz[7][8] = 9'b111111111;
assign micromatrizz[7][9] = 9'b111111111;
assign micromatrizz[7][10] = 9'b111111111;
assign micromatrizz[7][11] = 9'b111111111;
assign micromatrizz[7][12] = 9'b111111111;
assign micromatrizz[7][13] = 9'b111111111;
assign micromatrizz[7][14] = 9'b111111111;
assign micromatrizz[7][15] = 9'b111111111;
assign micromatrizz[7][16] = 9'b111111111;
assign micromatrizz[7][17] = 9'b111111111;
assign micromatrizz[7][18] = 9'b111111111;
assign micromatrizz[7][19] = 9'b111111111;
assign micromatrizz[7][20] = 9'b111111111;
assign micromatrizz[7][21] = 9'b111111111;
assign micromatrizz[7][22] = 9'b111111111;
assign micromatrizz[7][23] = 9'b111111111;
assign micromatrizz[7][24] = 9'b111111111;
assign micromatrizz[7][25] = 9'b111111111;
assign micromatrizz[7][26] = 9'b111111111;
assign micromatrizz[7][27] = 9'b111111111;
assign micromatrizz[7][28] = 9'b111111111;
assign micromatrizz[7][29] = 9'b111111111;
assign micromatrizz[7][30] = 9'b111111111;
assign micromatrizz[7][31] = 9'b111111111;
assign micromatrizz[7][32] = 9'b111111111;
assign micromatrizz[7][33] = 9'b111111111;
assign micromatrizz[7][34] = 9'b111111111;
assign micromatrizz[7][35] = 9'b111111111;
assign micromatrizz[7][36] = 9'b111111111;
assign micromatrizz[7][37] = 9'b111111111;
assign micromatrizz[7][38] = 9'b111111111;
assign micromatrizz[7][39] = 9'b111111111;
assign micromatrizz[7][40] = 9'b111111111;
assign micromatrizz[7][41] = 9'b111111111;
assign micromatrizz[7][42] = 9'b111111111;
assign micromatrizz[7][43] = 9'b111111111;
assign micromatrizz[7][44] = 9'b111111111;
assign micromatrizz[7][45] = 9'b111111111;
assign micromatrizz[7][46] = 9'b111111111;
assign micromatrizz[7][47] = 9'b111111111;
assign micromatrizz[7][48] = 9'b111111111;
assign micromatrizz[7][49] = 9'b111111111;
assign micromatrizz[7][50] = 9'b111111111;
assign micromatrizz[7][51] = 9'b111111111;
assign micromatrizz[7][52] = 9'b111111111;
assign micromatrizz[7][53] = 9'b111111111;
assign micromatrizz[7][54] = 9'b111111111;
assign micromatrizz[7][55] = 9'b111111111;
assign micromatrizz[7][56] = 9'b111111111;
assign micromatrizz[7][57] = 9'b111111111;
assign micromatrizz[7][58] = 9'b111111111;
assign micromatrizz[7][59] = 9'b111111111;
assign micromatrizz[7][60] = 9'b111111111;
assign micromatrizz[7][61] = 9'b111111111;
assign micromatrizz[7][62] = 9'b111111111;
assign micromatrizz[7][63] = 9'b111111111;
assign micromatrizz[7][64] = 9'b111111111;
assign micromatrizz[7][65] = 9'b111111111;
assign micromatrizz[7][66] = 9'b111111111;
assign micromatrizz[7][67] = 9'b111111111;
assign micromatrizz[7][68] = 9'b111111111;
assign micromatrizz[7][69] = 9'b111111111;
assign micromatrizz[7][70] = 9'b111111111;
assign micromatrizz[7][71] = 9'b111111111;
assign micromatrizz[7][72] = 9'b111111111;
assign micromatrizz[7][73] = 9'b111111111;
assign micromatrizz[7][74] = 9'b111111111;
assign micromatrizz[7][75] = 9'b111111111;
assign micromatrizz[7][76] = 9'b111111111;
assign micromatrizz[7][77] = 9'b111111111;
assign micromatrizz[7][78] = 9'b111111111;
assign micromatrizz[7][79] = 9'b111111111;
assign micromatrizz[7][80] = 9'b111111111;
assign micromatrizz[7][81] = 9'b111111111;
assign micromatrizz[7][82] = 9'b111111111;
assign micromatrizz[7][83] = 9'b111111111;
assign micromatrizz[7][84] = 9'b111111111;
assign micromatrizz[7][85] = 9'b111111111;
assign micromatrizz[7][86] = 9'b111111111;
assign micromatrizz[7][87] = 9'b111111111;
assign micromatrizz[7][88] = 9'b111111111;
assign micromatrizz[7][89] = 9'b111111111;
assign micromatrizz[7][90] = 9'b111111111;
assign micromatrizz[7][91] = 9'b111111111;
assign micromatrizz[7][92] = 9'b111111111;
assign micromatrizz[7][93] = 9'b111111111;
assign micromatrizz[7][94] = 9'b111111111;
assign micromatrizz[7][95] = 9'b111111111;
assign micromatrizz[7][96] = 9'b111111111;
assign micromatrizz[7][97] = 9'b111111111;
assign micromatrizz[7][98] = 9'b111111111;
assign micromatrizz[7][99] = 9'b111111111;
assign micromatrizz[7][100] = 9'b111111111;
assign micromatrizz[7][101] = 9'b111111111;
assign micromatrizz[7][102] = 9'b111111111;
assign micromatrizz[7][103] = 9'b111111111;
assign micromatrizz[7][104] = 9'b111111111;
assign micromatrizz[7][105] = 9'b111111111;
assign micromatrizz[7][106] = 9'b111111111;
assign micromatrizz[7][107] = 9'b111111111;
assign micromatrizz[7][108] = 9'b111111111;
assign micromatrizz[7][109] = 9'b111111111;
assign micromatrizz[7][110] = 9'b111111111;
assign micromatrizz[7][111] = 9'b111111111;
assign micromatrizz[7][112] = 9'b111111111;
assign micromatrizz[7][113] = 9'b111111111;
assign micromatrizz[7][114] = 9'b111111111;
assign micromatrizz[7][115] = 9'b111111111;
assign micromatrizz[7][116] = 9'b111111111;
assign micromatrizz[7][117] = 9'b111111111;
assign micromatrizz[7][118] = 9'b111111111;
assign micromatrizz[7][119] = 9'b111111111;
assign micromatrizz[7][120] = 9'b111111111;
assign micromatrizz[7][121] = 9'b111111111;
assign micromatrizz[7][122] = 9'b111111111;
assign micromatrizz[7][123] = 9'b111111111;
assign micromatrizz[7][124] = 9'b111111111;
assign micromatrizz[7][125] = 9'b111111111;
assign micromatrizz[7][126] = 9'b111111111;
assign micromatrizz[7][127] = 9'b111111111;
assign micromatrizz[7][128] = 9'b111111111;
assign micromatrizz[7][129] = 9'b111111111;
assign micromatrizz[7][130] = 9'b111111111;
assign micromatrizz[7][131] = 9'b111111111;
assign micromatrizz[7][132] = 9'b111111111;
assign micromatrizz[7][133] = 9'b111111111;
assign micromatrizz[7][134] = 9'b111111111;
assign micromatrizz[7][135] = 9'b111111111;
assign micromatrizz[7][136] = 9'b111111111;
assign micromatrizz[7][137] = 9'b111111111;
assign micromatrizz[7][138] = 9'b111111111;
assign micromatrizz[7][139] = 9'b111111111;
assign micromatrizz[7][140] = 9'b111111111;
assign micromatrizz[7][141] = 9'b111111111;
assign micromatrizz[7][142] = 9'b111111111;
assign micromatrizz[7][143] = 9'b111111111;
assign micromatrizz[7][144] = 9'b111111111;
assign micromatrizz[7][145] = 9'b111111111;
assign micromatrizz[7][146] = 9'b111111111;
assign micromatrizz[7][147] = 9'b111111111;
assign micromatrizz[7][148] = 9'b111111111;
assign micromatrizz[7][149] = 9'b111111111;
assign micromatrizz[7][150] = 9'b111111111;
assign micromatrizz[7][151] = 9'b111111111;
assign micromatrizz[7][152] = 9'b111111111;
assign micromatrizz[7][153] = 9'b111111111;
assign micromatrizz[7][154] = 9'b111111111;
assign micromatrizz[7][155] = 9'b111111111;
assign micromatrizz[7][156] = 9'b111111111;
assign micromatrizz[7][157] = 9'b111111111;
assign micromatrizz[7][158] = 9'b111111111;
assign micromatrizz[7][159] = 9'b111111111;
assign micromatrizz[7][160] = 9'b111111111;
assign micromatrizz[7][161] = 9'b111111111;
assign micromatrizz[7][162] = 9'b111111111;
assign micromatrizz[7][163] = 9'b111111111;
assign micromatrizz[7][164] = 9'b111111111;
assign micromatrizz[7][165] = 9'b111111111;
assign micromatrizz[7][166] = 9'b111111111;
assign micromatrizz[7][167] = 9'b111111111;
assign micromatrizz[7][168] = 9'b111111111;
assign micromatrizz[7][169] = 9'b111111111;
assign micromatrizz[7][170] = 9'b111111111;
assign micromatrizz[7][171] = 9'b111111111;
assign micromatrizz[7][172] = 9'b111111111;
assign micromatrizz[7][173] = 9'b111111111;
assign micromatrizz[7][174] = 9'b111111111;
assign micromatrizz[7][175] = 9'b111111111;
assign micromatrizz[7][176] = 9'b111111111;
assign micromatrizz[7][177] = 9'b111111111;
assign micromatrizz[7][178] = 9'b111111111;
assign micromatrizz[7][179] = 9'b111111111;
assign micromatrizz[7][180] = 9'b111111111;
assign micromatrizz[7][181] = 9'b111111111;
assign micromatrizz[7][182] = 9'b111111111;
assign micromatrizz[7][183] = 9'b111111111;
assign micromatrizz[7][184] = 9'b111111111;
assign micromatrizz[7][185] = 9'b111111111;
assign micromatrizz[7][186] = 9'b111111111;
assign micromatrizz[7][187] = 9'b111111111;
assign micromatrizz[7][188] = 9'b111111111;
assign micromatrizz[7][189] = 9'b111111111;
assign micromatrizz[7][190] = 9'b111111111;
assign micromatrizz[7][191] = 9'b111111111;
assign micromatrizz[7][192] = 9'b111111111;
assign micromatrizz[7][193] = 9'b111111111;
assign micromatrizz[7][194] = 9'b111111111;
assign micromatrizz[7][195] = 9'b111111111;
assign micromatrizz[7][196] = 9'b111111111;
assign micromatrizz[7][197] = 9'b111111111;
assign micromatrizz[7][198] = 9'b111111111;
assign micromatrizz[7][199] = 9'b111111111;
assign micromatrizz[7][200] = 9'b111111111;
assign micromatrizz[7][201] = 9'b111111111;
assign micromatrizz[7][202] = 9'b111111111;
assign micromatrizz[7][203] = 9'b111111111;
assign micromatrizz[7][204] = 9'b111111111;
assign micromatrizz[7][205] = 9'b111111111;
assign micromatrizz[7][206] = 9'b111111111;
assign micromatrizz[7][207] = 9'b111111111;
assign micromatrizz[7][208] = 9'b111111111;
assign micromatrizz[7][209] = 9'b111111111;
assign micromatrizz[7][210] = 9'b111111111;
assign micromatrizz[7][211] = 9'b111111111;
assign micromatrizz[7][212] = 9'b111111111;
assign micromatrizz[7][213] = 9'b111111111;
assign micromatrizz[7][214] = 9'b111111111;
assign micromatrizz[7][215] = 9'b111111111;
assign micromatrizz[7][216] = 9'b111111111;
assign micromatrizz[7][217] = 9'b111111111;
assign micromatrizz[7][218] = 9'b111111111;
assign micromatrizz[7][219] = 9'b111111111;
assign micromatrizz[7][220] = 9'b111111111;
assign micromatrizz[7][221] = 9'b111111111;
assign micromatrizz[7][222] = 9'b111111111;
assign micromatrizz[7][223] = 9'b111111111;
assign micromatrizz[7][224] = 9'b111111111;
assign micromatrizz[7][225] = 9'b111111111;
assign micromatrizz[7][226] = 9'b111111111;
assign micromatrizz[7][227] = 9'b111111111;
assign micromatrizz[7][228] = 9'b111111111;
assign micromatrizz[7][229] = 9'b111111111;
assign micromatrizz[7][230] = 9'b111111111;
assign micromatrizz[7][231] = 9'b111111111;
assign micromatrizz[7][232] = 9'b111111111;
assign micromatrizz[7][233] = 9'b111111111;
assign micromatrizz[7][234] = 9'b111111111;
assign micromatrizz[7][235] = 9'b111111111;
assign micromatrizz[7][236] = 9'b111111111;
assign micromatrizz[7][237] = 9'b111111111;
assign micromatrizz[7][238] = 9'b111111111;
assign micromatrizz[7][239] = 9'b111111111;
assign micromatrizz[7][240] = 9'b111111111;
assign micromatrizz[7][241] = 9'b111111111;
assign micromatrizz[7][242] = 9'b111111111;
assign micromatrizz[7][243] = 9'b111111111;
assign micromatrizz[7][244] = 9'b111111111;
assign micromatrizz[7][245] = 9'b111111111;
assign micromatrizz[7][246] = 9'b111111111;
assign micromatrizz[7][247] = 9'b111111111;
assign micromatrizz[7][248] = 9'b111111111;
assign micromatrizz[7][249] = 9'b111111111;
assign micromatrizz[7][250] = 9'b111111111;
assign micromatrizz[7][251] = 9'b111111111;
assign micromatrizz[7][252] = 9'b111111111;
assign micromatrizz[7][253] = 9'b111111111;
assign micromatrizz[7][254] = 9'b111111111;
assign micromatrizz[7][255] = 9'b111111111;
assign micromatrizz[7][256] = 9'b111111111;
assign micromatrizz[7][257] = 9'b111111111;
assign micromatrizz[7][258] = 9'b111111111;
assign micromatrizz[7][259] = 9'b111111111;
assign micromatrizz[7][260] = 9'b111111111;
assign micromatrizz[7][261] = 9'b111111111;
assign micromatrizz[7][262] = 9'b111111111;
assign micromatrizz[7][263] = 9'b111111111;
assign micromatrizz[7][264] = 9'b111111111;
assign micromatrizz[7][265] = 9'b111111111;
assign micromatrizz[7][266] = 9'b111111111;
assign micromatrizz[7][267] = 9'b111111111;
assign micromatrizz[7][268] = 9'b111111111;
assign micromatrizz[7][269] = 9'b111111111;
assign micromatrizz[7][270] = 9'b111111111;
assign micromatrizz[7][271] = 9'b111111111;
assign micromatrizz[7][272] = 9'b111111111;
assign micromatrizz[7][273] = 9'b111111111;
assign micromatrizz[7][274] = 9'b111111111;
assign micromatrizz[7][275] = 9'b111111111;
assign micromatrizz[7][276] = 9'b111111111;
assign micromatrizz[7][277] = 9'b111111111;
assign micromatrizz[7][278] = 9'b111111111;
assign micromatrizz[7][279] = 9'b111111111;
assign micromatrizz[7][280] = 9'b111111111;
assign micromatrizz[7][281] = 9'b111111111;
assign micromatrizz[7][282] = 9'b111111111;
assign micromatrizz[7][283] = 9'b111111111;
assign micromatrizz[7][284] = 9'b111111111;
assign micromatrizz[7][285] = 9'b111111111;
assign micromatrizz[7][286] = 9'b111111111;
assign micromatrizz[7][287] = 9'b111111111;
assign micromatrizz[7][288] = 9'b111111111;
assign micromatrizz[7][289] = 9'b111111111;
assign micromatrizz[7][290] = 9'b111111111;
assign micromatrizz[7][291] = 9'b111111111;
assign micromatrizz[7][292] = 9'b111111111;
assign micromatrizz[7][293] = 9'b111111111;
assign micromatrizz[7][294] = 9'b111111111;
assign micromatrizz[7][295] = 9'b111111111;
assign micromatrizz[7][296] = 9'b111111111;
assign micromatrizz[7][297] = 9'b111111111;
assign micromatrizz[7][298] = 9'b111111111;
assign micromatrizz[7][299] = 9'b111111111;
assign micromatrizz[7][300] = 9'b111111111;
assign micromatrizz[7][301] = 9'b111111111;
assign micromatrizz[7][302] = 9'b111111111;
assign micromatrizz[7][303] = 9'b111111111;
assign micromatrizz[7][304] = 9'b111111111;
assign micromatrizz[7][305] = 9'b111111111;
assign micromatrizz[7][306] = 9'b111111111;
assign micromatrizz[7][307] = 9'b111111111;
assign micromatrizz[7][308] = 9'b111111111;
assign micromatrizz[7][309] = 9'b111111111;
assign micromatrizz[7][310] = 9'b111111111;
assign micromatrizz[7][311] = 9'b111111111;
assign micromatrizz[7][312] = 9'b111111111;
assign micromatrizz[7][313] = 9'b111111111;
assign micromatrizz[7][314] = 9'b111111111;
assign micromatrizz[7][315] = 9'b111111111;
assign micromatrizz[7][316] = 9'b111111111;
assign micromatrizz[7][317] = 9'b111111111;
assign micromatrizz[7][318] = 9'b111111111;
assign micromatrizz[7][319] = 9'b111111111;
assign micromatrizz[7][320] = 9'b111111111;
assign micromatrizz[7][321] = 9'b111111111;
assign micromatrizz[7][322] = 9'b111111111;
assign micromatrizz[7][323] = 9'b111111111;
assign micromatrizz[7][324] = 9'b111111111;
assign micromatrizz[7][325] = 9'b111111111;
assign micromatrizz[7][326] = 9'b111111111;
assign micromatrizz[7][327] = 9'b111111111;
assign micromatrizz[7][328] = 9'b111111111;
assign micromatrizz[7][329] = 9'b111111111;
assign micromatrizz[7][330] = 9'b111111111;
assign micromatrizz[7][331] = 9'b111111111;
assign micromatrizz[7][332] = 9'b111111111;
assign micromatrizz[7][333] = 9'b111111111;
assign micromatrizz[7][334] = 9'b111111111;
assign micromatrizz[7][335] = 9'b111111111;
assign micromatrizz[7][336] = 9'b111111111;
assign micromatrizz[7][337] = 9'b111111111;
assign micromatrizz[7][338] = 9'b111111111;
assign micromatrizz[7][339] = 9'b111111111;
assign micromatrizz[7][340] = 9'b111111111;
assign micromatrizz[7][341] = 9'b111111111;
assign micromatrizz[7][342] = 9'b111111111;
assign micromatrizz[7][343] = 9'b111111111;
assign micromatrizz[7][344] = 9'b111111111;
assign micromatrizz[7][345] = 9'b111111111;
assign micromatrizz[7][346] = 9'b111111111;
assign micromatrizz[7][347] = 9'b111111111;
assign micromatrizz[7][348] = 9'b111111111;
assign micromatrizz[7][349] = 9'b111111111;
assign micromatrizz[7][350] = 9'b111111111;
assign micromatrizz[7][351] = 9'b111111111;
assign micromatrizz[7][352] = 9'b111111111;
assign micromatrizz[7][353] = 9'b111111111;
assign micromatrizz[7][354] = 9'b111111111;
assign micromatrizz[7][355] = 9'b111111111;
assign micromatrizz[7][356] = 9'b111111111;
assign micromatrizz[7][357] = 9'b111111111;
assign micromatrizz[7][358] = 9'b111111111;
assign micromatrizz[7][359] = 9'b111111111;
assign micromatrizz[7][360] = 9'b111111111;
assign micromatrizz[7][361] = 9'b111111111;
assign micromatrizz[7][362] = 9'b111111111;
assign micromatrizz[7][363] = 9'b111111111;
assign micromatrizz[7][364] = 9'b111111111;
assign micromatrizz[7][365] = 9'b111111111;
assign micromatrizz[7][366] = 9'b111111111;
assign micromatrizz[7][367] = 9'b111111111;
assign micromatrizz[7][368] = 9'b111111111;
assign micromatrizz[7][369] = 9'b111111111;
assign micromatrizz[7][370] = 9'b111111111;
assign micromatrizz[7][371] = 9'b111111111;
assign micromatrizz[7][372] = 9'b111111111;
assign micromatrizz[7][373] = 9'b111111111;
assign micromatrizz[7][374] = 9'b111111111;
assign micromatrizz[7][375] = 9'b111111111;
assign micromatrizz[7][376] = 9'b111111111;
assign micromatrizz[7][377] = 9'b111111111;
assign micromatrizz[7][378] = 9'b111111111;
assign micromatrizz[7][379] = 9'b111111111;
assign micromatrizz[7][380] = 9'b111111111;
assign micromatrizz[7][381] = 9'b111111111;
assign micromatrizz[7][382] = 9'b111111111;
assign micromatrizz[7][383] = 9'b111111111;
assign micromatrizz[7][384] = 9'b111111111;
assign micromatrizz[7][385] = 9'b111111111;
assign micromatrizz[7][386] = 9'b111111111;
assign micromatrizz[7][387] = 9'b111111111;
assign micromatrizz[7][388] = 9'b111111111;
assign micromatrizz[7][389] = 9'b111111111;
assign micromatrizz[7][390] = 9'b111111111;
assign micromatrizz[7][391] = 9'b111111111;
assign micromatrizz[7][392] = 9'b111111111;
assign micromatrizz[7][393] = 9'b111111111;
assign micromatrizz[7][394] = 9'b111111111;
assign micromatrizz[7][395] = 9'b111111111;
assign micromatrizz[7][396] = 9'b111111111;
assign micromatrizz[7][397] = 9'b111111111;
assign micromatrizz[7][398] = 9'b111111111;
assign micromatrizz[7][399] = 9'b111111111;
assign micromatrizz[7][400] = 9'b111111111;
assign micromatrizz[7][401] = 9'b111111111;
assign micromatrizz[7][402] = 9'b111111111;
assign micromatrizz[7][403] = 9'b111111111;
assign micromatrizz[7][404] = 9'b111111111;
assign micromatrizz[7][405] = 9'b111111111;
assign micromatrizz[7][406] = 9'b111111111;
assign micromatrizz[7][407] = 9'b111111111;
assign micromatrizz[7][408] = 9'b111111111;
assign micromatrizz[7][409] = 9'b111111111;
assign micromatrizz[7][410] = 9'b111111111;
assign micromatrizz[7][411] = 9'b111111111;
assign micromatrizz[7][412] = 9'b111111111;
assign micromatrizz[7][413] = 9'b111111111;
assign micromatrizz[7][414] = 9'b111111111;
assign micromatrizz[7][415] = 9'b111111111;
assign micromatrizz[7][416] = 9'b111111111;
assign micromatrizz[7][417] = 9'b111111111;
assign micromatrizz[7][418] = 9'b111111111;
assign micromatrizz[7][419] = 9'b111111111;
assign micromatrizz[7][420] = 9'b111111111;
assign micromatrizz[7][421] = 9'b111111111;
assign micromatrizz[7][422] = 9'b111111111;
assign micromatrizz[7][423] = 9'b111111111;
assign micromatrizz[7][424] = 9'b111111111;
assign micromatrizz[7][425] = 9'b111111111;
assign micromatrizz[7][426] = 9'b111111111;
assign micromatrizz[7][427] = 9'b111111111;
assign micromatrizz[7][428] = 9'b111111111;
assign micromatrizz[7][429] = 9'b111111111;
assign micromatrizz[7][430] = 9'b111111111;
assign micromatrizz[7][431] = 9'b111111111;
assign micromatrizz[7][432] = 9'b111111111;
assign micromatrizz[7][433] = 9'b111111111;
assign micromatrizz[7][434] = 9'b111111111;
assign micromatrizz[7][435] = 9'b111111111;
assign micromatrizz[7][436] = 9'b111111111;
assign micromatrizz[7][437] = 9'b111111111;
assign micromatrizz[7][438] = 9'b111111111;
assign micromatrizz[7][439] = 9'b111111111;
assign micromatrizz[7][440] = 9'b111111111;
assign micromatrizz[7][441] = 9'b111111111;
assign micromatrizz[7][442] = 9'b111111111;
assign micromatrizz[7][443] = 9'b111111111;
assign micromatrizz[7][444] = 9'b111111111;
assign micromatrizz[7][445] = 9'b111111111;
assign micromatrizz[7][446] = 9'b111111111;
assign micromatrizz[7][447] = 9'b111111111;
assign micromatrizz[7][448] = 9'b111111111;
assign micromatrizz[7][449] = 9'b111111111;
assign micromatrizz[7][450] = 9'b111111111;
assign micromatrizz[7][451] = 9'b111111111;
assign micromatrizz[7][452] = 9'b111111111;
assign micromatrizz[7][453] = 9'b111111111;
assign micromatrizz[7][454] = 9'b111111111;
assign micromatrizz[7][455] = 9'b111111111;
assign micromatrizz[7][456] = 9'b111111111;
assign micromatrizz[7][457] = 9'b111111111;
assign micromatrizz[7][458] = 9'b111111111;
assign micromatrizz[7][459] = 9'b111111111;
assign micromatrizz[7][460] = 9'b111111111;
assign micromatrizz[7][461] = 9'b111111111;
assign micromatrizz[7][462] = 9'b111111111;
assign micromatrizz[7][463] = 9'b111111111;
assign micromatrizz[7][464] = 9'b111111111;
assign micromatrizz[7][465] = 9'b111111111;
assign micromatrizz[7][466] = 9'b111111111;
assign micromatrizz[7][467] = 9'b111111111;
assign micromatrizz[7][468] = 9'b111111111;
assign micromatrizz[7][469] = 9'b111111111;
assign micromatrizz[7][470] = 9'b111111111;
assign micromatrizz[7][471] = 9'b111111111;
assign micromatrizz[7][472] = 9'b111111111;
assign micromatrizz[7][473] = 9'b111111111;
assign micromatrizz[7][474] = 9'b111111111;
assign micromatrizz[7][475] = 9'b111111111;
assign micromatrizz[7][476] = 9'b111111111;
assign micromatrizz[7][477] = 9'b111111111;
assign micromatrizz[7][478] = 9'b111111111;
assign micromatrizz[7][479] = 9'b111111111;
assign micromatrizz[7][480] = 9'b111111111;
assign micromatrizz[7][481] = 9'b111111111;
assign micromatrizz[7][482] = 9'b111111111;
assign micromatrizz[7][483] = 9'b111111111;
assign micromatrizz[7][484] = 9'b111111111;
assign micromatrizz[7][485] = 9'b111111111;
assign micromatrizz[7][486] = 9'b111111111;
assign micromatrizz[7][487] = 9'b111111111;
assign micromatrizz[7][488] = 9'b111111111;
assign micromatrizz[7][489] = 9'b111111111;
assign micromatrizz[7][490] = 9'b111111111;
assign micromatrizz[7][491] = 9'b111111111;
assign micromatrizz[7][492] = 9'b111111111;
assign micromatrizz[7][493] = 9'b111111111;
assign micromatrizz[7][494] = 9'b111111111;
assign micromatrizz[7][495] = 9'b111111111;
assign micromatrizz[7][496] = 9'b111111111;
assign micromatrizz[7][497] = 9'b111111111;
assign micromatrizz[7][498] = 9'b111111111;
assign micromatrizz[7][499] = 9'b111111111;
assign micromatrizz[7][500] = 9'b111111111;
assign micromatrizz[7][501] = 9'b111111111;
assign micromatrizz[7][502] = 9'b111111111;
assign micromatrizz[7][503] = 9'b111111111;
assign micromatrizz[7][504] = 9'b111111111;
assign micromatrizz[7][505] = 9'b111111111;
assign micromatrizz[7][506] = 9'b111111111;
assign micromatrizz[7][507] = 9'b111111111;
assign micromatrizz[7][508] = 9'b111111111;
assign micromatrizz[7][509] = 9'b111111111;
assign micromatrizz[7][510] = 9'b111111111;
assign micromatrizz[7][511] = 9'b111111111;
assign micromatrizz[7][512] = 9'b111111111;
assign micromatrizz[7][513] = 9'b111111111;
assign micromatrizz[7][514] = 9'b111111111;
assign micromatrizz[7][515] = 9'b111111111;
assign micromatrizz[7][516] = 9'b111111111;
assign micromatrizz[7][517] = 9'b111111111;
assign micromatrizz[7][518] = 9'b111111111;
assign micromatrizz[7][519] = 9'b111111111;
assign micromatrizz[7][520] = 9'b111111111;
assign micromatrizz[7][521] = 9'b111111111;
assign micromatrizz[7][522] = 9'b111111111;
assign micromatrizz[7][523] = 9'b111111111;
assign micromatrizz[7][524] = 9'b111111111;
assign micromatrizz[7][525] = 9'b111111111;
assign micromatrizz[7][526] = 9'b111111111;
assign micromatrizz[7][527] = 9'b111111111;
assign micromatrizz[7][528] = 9'b111111111;
assign micromatrizz[7][529] = 9'b111111111;
assign micromatrizz[7][530] = 9'b111111111;
assign micromatrizz[7][531] = 9'b111111111;
assign micromatrizz[7][532] = 9'b111111111;
assign micromatrizz[7][533] = 9'b111111111;
assign micromatrizz[7][534] = 9'b111111111;
assign micromatrizz[7][535] = 9'b111111111;
assign micromatrizz[7][536] = 9'b111111111;
assign micromatrizz[7][537] = 9'b111111111;
assign micromatrizz[7][538] = 9'b111111111;
assign micromatrizz[7][539] = 9'b111111111;
assign micromatrizz[7][540] = 9'b111111111;
assign micromatrizz[7][541] = 9'b111111111;
assign micromatrizz[7][542] = 9'b111111111;
assign micromatrizz[7][543] = 9'b111111111;
assign micromatrizz[7][544] = 9'b111111111;
assign micromatrizz[7][545] = 9'b111111111;
assign micromatrizz[7][546] = 9'b111111111;
assign micromatrizz[7][547] = 9'b111111111;
assign micromatrizz[7][548] = 9'b111111111;
assign micromatrizz[7][549] = 9'b111111111;
assign micromatrizz[7][550] = 9'b111111111;
assign micromatrizz[7][551] = 9'b111111111;
assign micromatrizz[7][552] = 9'b111111111;
assign micromatrizz[7][553] = 9'b111111111;
assign micromatrizz[7][554] = 9'b111111111;
assign micromatrizz[7][555] = 9'b111111111;
assign micromatrizz[7][556] = 9'b111111111;
assign micromatrizz[7][557] = 9'b111111111;
assign micromatrizz[7][558] = 9'b111111111;
assign micromatrizz[7][559] = 9'b111111111;
assign micromatrizz[7][560] = 9'b111111111;
assign micromatrizz[7][561] = 9'b111111111;
assign micromatrizz[7][562] = 9'b111111111;
assign micromatrizz[7][563] = 9'b111111111;
assign micromatrizz[7][564] = 9'b111111111;
assign micromatrizz[7][565] = 9'b111111111;
assign micromatrizz[7][566] = 9'b111111111;
assign micromatrizz[7][567] = 9'b111111111;
assign micromatrizz[7][568] = 9'b111111111;
assign micromatrizz[7][569] = 9'b111111111;
assign micromatrizz[7][570] = 9'b111111111;
assign micromatrizz[7][571] = 9'b111111111;
assign micromatrizz[7][572] = 9'b111111111;
assign micromatrizz[7][573] = 9'b111111111;
assign micromatrizz[7][574] = 9'b111111111;
assign micromatrizz[7][575] = 9'b111111111;
assign micromatrizz[7][576] = 9'b111111111;
assign micromatrizz[7][577] = 9'b111111111;
assign micromatrizz[7][578] = 9'b111111111;
assign micromatrizz[7][579] = 9'b111111111;
assign micromatrizz[7][580] = 9'b111111111;
assign micromatrizz[7][581] = 9'b111111111;
assign micromatrizz[7][582] = 9'b111111111;
assign micromatrizz[7][583] = 9'b111111111;
assign micromatrizz[7][584] = 9'b111111111;
assign micromatrizz[7][585] = 9'b111111111;
assign micromatrizz[7][586] = 9'b111111111;
assign micromatrizz[7][587] = 9'b111111111;
assign micromatrizz[7][588] = 9'b111111111;
assign micromatrizz[7][589] = 9'b111111111;
assign micromatrizz[7][590] = 9'b111111111;
assign micromatrizz[7][591] = 9'b111111111;
assign micromatrizz[7][592] = 9'b111111111;
assign micromatrizz[7][593] = 9'b111111111;
assign micromatrizz[7][594] = 9'b111111111;
assign micromatrizz[7][595] = 9'b111111111;
assign micromatrizz[7][596] = 9'b111111111;
assign micromatrizz[7][597] = 9'b111111111;
assign micromatrizz[7][598] = 9'b111111111;
assign micromatrizz[7][599] = 9'b111111111;
assign micromatrizz[7][600] = 9'b111111111;
assign micromatrizz[7][601] = 9'b111111111;
assign micromatrizz[7][602] = 9'b111111111;
assign micromatrizz[7][603] = 9'b111111111;
assign micromatrizz[7][604] = 9'b111111111;
assign micromatrizz[7][605] = 9'b111111111;
assign micromatrizz[7][606] = 9'b111111111;
assign micromatrizz[7][607] = 9'b111111111;
assign micromatrizz[7][608] = 9'b111111111;
assign micromatrizz[7][609] = 9'b111111111;
assign micromatrizz[7][610] = 9'b111111111;
assign micromatrizz[7][611] = 9'b111111111;
assign micromatrizz[7][612] = 9'b111111111;
assign micromatrizz[7][613] = 9'b111111111;
assign micromatrizz[7][614] = 9'b111111111;
assign micromatrizz[7][615] = 9'b111111111;
assign micromatrizz[7][616] = 9'b111111111;
assign micromatrizz[7][617] = 9'b111111111;
assign micromatrizz[7][618] = 9'b111111111;
assign micromatrizz[7][619] = 9'b111111111;
assign micromatrizz[7][620] = 9'b111111111;
assign micromatrizz[7][621] = 9'b111111111;
assign micromatrizz[7][622] = 9'b111111111;
assign micromatrizz[7][623] = 9'b111111111;
assign micromatrizz[7][624] = 9'b111111111;
assign micromatrizz[7][625] = 9'b111111111;
assign micromatrizz[7][626] = 9'b111111111;
assign micromatrizz[7][627] = 9'b111111111;
assign micromatrizz[7][628] = 9'b111111111;
assign micromatrizz[7][629] = 9'b111111111;
assign micromatrizz[7][630] = 9'b111111111;
assign micromatrizz[7][631] = 9'b111111111;
assign micromatrizz[7][632] = 9'b111111111;
assign micromatrizz[7][633] = 9'b111111111;
assign micromatrizz[7][634] = 9'b111111111;
assign micromatrizz[7][635] = 9'b111111111;
assign micromatrizz[7][636] = 9'b111111111;
assign micromatrizz[7][637] = 9'b111111111;
assign micromatrizz[7][638] = 9'b111111111;
assign micromatrizz[7][639] = 9'b111111111;
assign micromatrizz[8][0] = 9'b111111111;
assign micromatrizz[8][1] = 9'b111111111;
assign micromatrizz[8][2] = 9'b111111111;
assign micromatrizz[8][3] = 9'b111111111;
assign micromatrizz[8][4] = 9'b111111111;
assign micromatrizz[8][5] = 9'b111111111;
assign micromatrizz[8][6] = 9'b111111111;
assign micromatrizz[8][7] = 9'b111111111;
assign micromatrizz[8][8] = 9'b111111111;
assign micromatrizz[8][9] = 9'b111111111;
assign micromatrizz[8][10] = 9'b111111111;
assign micromatrizz[8][11] = 9'b111111111;
assign micromatrizz[8][12] = 9'b111111111;
assign micromatrizz[8][13] = 9'b111111111;
assign micromatrizz[8][14] = 9'b111111111;
assign micromatrizz[8][15] = 9'b111111111;
assign micromatrizz[8][16] = 9'b111111111;
assign micromatrizz[8][17] = 9'b111111111;
assign micromatrizz[8][18] = 9'b111111111;
assign micromatrizz[8][19] = 9'b111111111;
assign micromatrizz[8][20] = 9'b111111111;
assign micromatrizz[8][21] = 9'b111111111;
assign micromatrizz[8][22] = 9'b111111111;
assign micromatrizz[8][23] = 9'b111111111;
assign micromatrizz[8][24] = 9'b111111111;
assign micromatrizz[8][25] = 9'b111111111;
assign micromatrizz[8][26] = 9'b111111111;
assign micromatrizz[8][27] = 9'b111111111;
assign micromatrizz[8][28] = 9'b111111111;
assign micromatrizz[8][29] = 9'b111111111;
assign micromatrizz[8][30] = 9'b111111111;
assign micromatrizz[8][31] = 9'b111111111;
assign micromatrizz[8][32] = 9'b111111111;
assign micromatrizz[8][33] = 9'b111111111;
assign micromatrizz[8][34] = 9'b111111111;
assign micromatrizz[8][35] = 9'b111111111;
assign micromatrizz[8][36] = 9'b111111111;
assign micromatrizz[8][37] = 9'b111111111;
assign micromatrizz[8][38] = 9'b111111111;
assign micromatrizz[8][39] = 9'b111111111;
assign micromatrizz[8][40] = 9'b111111111;
assign micromatrizz[8][41] = 9'b111111111;
assign micromatrizz[8][42] = 9'b111111111;
assign micromatrizz[8][43] = 9'b111111111;
assign micromatrizz[8][44] = 9'b111111111;
assign micromatrizz[8][45] = 9'b111111111;
assign micromatrizz[8][46] = 9'b111111111;
assign micromatrizz[8][47] = 9'b111111111;
assign micromatrizz[8][48] = 9'b111111111;
assign micromatrizz[8][49] = 9'b111111111;
assign micromatrizz[8][50] = 9'b111111111;
assign micromatrizz[8][51] = 9'b111111111;
assign micromatrizz[8][52] = 9'b111111111;
assign micromatrizz[8][53] = 9'b111111111;
assign micromatrizz[8][54] = 9'b111111111;
assign micromatrizz[8][55] = 9'b111111111;
assign micromatrizz[8][56] = 9'b111111111;
assign micromatrizz[8][57] = 9'b111111111;
assign micromatrizz[8][58] = 9'b111111111;
assign micromatrizz[8][59] = 9'b111111111;
assign micromatrizz[8][60] = 9'b111111111;
assign micromatrizz[8][61] = 9'b111111111;
assign micromatrizz[8][62] = 9'b111111111;
assign micromatrizz[8][63] = 9'b111111111;
assign micromatrizz[8][64] = 9'b111111111;
assign micromatrizz[8][65] = 9'b111111111;
assign micromatrizz[8][66] = 9'b111111111;
assign micromatrizz[8][67] = 9'b111111111;
assign micromatrizz[8][68] = 9'b111111111;
assign micromatrizz[8][69] = 9'b111111111;
assign micromatrizz[8][70] = 9'b111111111;
assign micromatrizz[8][71] = 9'b111111111;
assign micromatrizz[8][72] = 9'b111111111;
assign micromatrizz[8][73] = 9'b111111111;
assign micromatrizz[8][74] = 9'b111111111;
assign micromatrizz[8][75] = 9'b111111111;
assign micromatrizz[8][76] = 9'b111111111;
assign micromatrizz[8][77] = 9'b111111111;
assign micromatrizz[8][78] = 9'b111111111;
assign micromatrizz[8][79] = 9'b111111111;
assign micromatrizz[8][80] = 9'b111111111;
assign micromatrizz[8][81] = 9'b111111111;
assign micromatrizz[8][82] = 9'b111111111;
assign micromatrizz[8][83] = 9'b111111111;
assign micromatrizz[8][84] = 9'b111111111;
assign micromatrizz[8][85] = 9'b111111111;
assign micromatrizz[8][86] = 9'b111111111;
assign micromatrizz[8][87] = 9'b111111111;
assign micromatrizz[8][88] = 9'b111111111;
assign micromatrizz[8][89] = 9'b111111111;
assign micromatrizz[8][90] = 9'b111111111;
assign micromatrizz[8][91] = 9'b111111111;
assign micromatrizz[8][92] = 9'b111111111;
assign micromatrizz[8][93] = 9'b111111111;
assign micromatrizz[8][94] = 9'b111111111;
assign micromatrizz[8][95] = 9'b111111111;
assign micromatrizz[8][96] = 9'b111111111;
assign micromatrizz[8][97] = 9'b111111111;
assign micromatrizz[8][98] = 9'b111111111;
assign micromatrizz[8][99] = 9'b111111111;
assign micromatrizz[8][100] = 9'b111111111;
assign micromatrizz[8][101] = 9'b111111111;
assign micromatrizz[8][102] = 9'b111111111;
assign micromatrizz[8][103] = 9'b111111111;
assign micromatrizz[8][104] = 9'b111111111;
assign micromatrizz[8][105] = 9'b111111111;
assign micromatrizz[8][106] = 9'b111111111;
assign micromatrizz[8][107] = 9'b111111111;
assign micromatrizz[8][108] = 9'b111111111;
assign micromatrizz[8][109] = 9'b111111111;
assign micromatrizz[8][110] = 9'b111111111;
assign micromatrizz[8][111] = 9'b111111111;
assign micromatrizz[8][112] = 9'b111111111;
assign micromatrizz[8][113] = 9'b111111111;
assign micromatrizz[8][114] = 9'b111111111;
assign micromatrizz[8][115] = 9'b111111111;
assign micromatrizz[8][116] = 9'b111111111;
assign micromatrizz[8][117] = 9'b111111111;
assign micromatrizz[8][118] = 9'b111111111;
assign micromatrizz[8][119] = 9'b111111111;
assign micromatrizz[8][120] = 9'b111111111;
assign micromatrizz[8][121] = 9'b111111111;
assign micromatrizz[8][122] = 9'b111111111;
assign micromatrizz[8][123] = 9'b111111111;
assign micromatrizz[8][124] = 9'b111111111;
assign micromatrizz[8][125] = 9'b111111111;
assign micromatrizz[8][126] = 9'b111111111;
assign micromatrizz[8][127] = 9'b111111111;
assign micromatrizz[8][128] = 9'b111111111;
assign micromatrizz[8][129] = 9'b111111111;
assign micromatrizz[8][130] = 9'b111111111;
assign micromatrizz[8][131] = 9'b111111111;
assign micromatrizz[8][132] = 9'b111111111;
assign micromatrizz[8][133] = 9'b111111111;
assign micromatrizz[8][134] = 9'b111111111;
assign micromatrizz[8][135] = 9'b111111111;
assign micromatrizz[8][136] = 9'b111111111;
assign micromatrizz[8][137] = 9'b111111111;
assign micromatrizz[8][138] = 9'b111111111;
assign micromatrizz[8][139] = 9'b111111111;
assign micromatrizz[8][140] = 9'b111111111;
assign micromatrizz[8][141] = 9'b111111111;
assign micromatrizz[8][142] = 9'b111111111;
assign micromatrizz[8][143] = 9'b111111111;
assign micromatrizz[8][144] = 9'b111111111;
assign micromatrizz[8][145] = 9'b111111111;
assign micromatrizz[8][146] = 9'b111111111;
assign micromatrizz[8][147] = 9'b111111111;
assign micromatrizz[8][148] = 9'b111111111;
assign micromatrizz[8][149] = 9'b111111111;
assign micromatrizz[8][150] = 9'b111111111;
assign micromatrizz[8][151] = 9'b111111111;
assign micromatrizz[8][152] = 9'b111111111;
assign micromatrizz[8][153] = 9'b111111111;
assign micromatrizz[8][154] = 9'b111111111;
assign micromatrizz[8][155] = 9'b111111111;
assign micromatrizz[8][156] = 9'b111111111;
assign micromatrizz[8][157] = 9'b111111111;
assign micromatrizz[8][158] = 9'b111111111;
assign micromatrizz[8][159] = 9'b111111111;
assign micromatrizz[8][160] = 9'b111111111;
assign micromatrizz[8][161] = 9'b111111111;
assign micromatrizz[8][162] = 9'b111111111;
assign micromatrizz[8][163] = 9'b111111111;
assign micromatrizz[8][164] = 9'b111111111;
assign micromatrizz[8][165] = 9'b111111111;
assign micromatrizz[8][166] = 9'b111111111;
assign micromatrizz[8][167] = 9'b111111111;
assign micromatrizz[8][168] = 9'b111111111;
assign micromatrizz[8][169] = 9'b111111111;
assign micromatrizz[8][170] = 9'b111111111;
assign micromatrizz[8][171] = 9'b111111111;
assign micromatrizz[8][172] = 9'b111111111;
assign micromatrizz[8][173] = 9'b111111111;
assign micromatrizz[8][174] = 9'b111111111;
assign micromatrizz[8][175] = 9'b111111111;
assign micromatrizz[8][176] = 9'b111111111;
assign micromatrizz[8][177] = 9'b111111111;
assign micromatrizz[8][178] = 9'b111111111;
assign micromatrizz[8][179] = 9'b111111111;
assign micromatrizz[8][180] = 9'b111111111;
assign micromatrizz[8][181] = 9'b111111111;
assign micromatrizz[8][182] = 9'b111111111;
assign micromatrizz[8][183] = 9'b111111111;
assign micromatrizz[8][184] = 9'b111111111;
assign micromatrizz[8][185] = 9'b111111111;
assign micromatrizz[8][186] = 9'b111111111;
assign micromatrizz[8][187] = 9'b111111111;
assign micromatrizz[8][188] = 9'b111111111;
assign micromatrizz[8][189] = 9'b111111111;
assign micromatrizz[8][190] = 9'b111111111;
assign micromatrizz[8][191] = 9'b111111111;
assign micromatrizz[8][192] = 9'b111111111;
assign micromatrizz[8][193] = 9'b111111111;
assign micromatrizz[8][194] = 9'b111111111;
assign micromatrizz[8][195] = 9'b111111111;
assign micromatrizz[8][196] = 9'b111111111;
assign micromatrizz[8][197] = 9'b111111111;
assign micromatrizz[8][198] = 9'b111111111;
assign micromatrizz[8][199] = 9'b111111111;
assign micromatrizz[8][200] = 9'b111111111;
assign micromatrizz[8][201] = 9'b111111111;
assign micromatrizz[8][202] = 9'b111111111;
assign micromatrizz[8][203] = 9'b111111111;
assign micromatrizz[8][204] = 9'b111111111;
assign micromatrizz[8][205] = 9'b111111111;
assign micromatrizz[8][206] = 9'b111111111;
assign micromatrizz[8][207] = 9'b111111111;
assign micromatrizz[8][208] = 9'b111111111;
assign micromatrizz[8][209] = 9'b111111111;
assign micromatrizz[8][210] = 9'b111111111;
assign micromatrizz[8][211] = 9'b111111111;
assign micromatrizz[8][212] = 9'b111111111;
assign micromatrizz[8][213] = 9'b111111111;
assign micromatrizz[8][214] = 9'b111111111;
assign micromatrizz[8][215] = 9'b111111111;
assign micromatrizz[8][216] = 9'b111111111;
assign micromatrizz[8][217] = 9'b111111111;
assign micromatrizz[8][218] = 9'b111111111;
assign micromatrizz[8][219] = 9'b111111111;
assign micromatrizz[8][220] = 9'b111111111;
assign micromatrizz[8][221] = 9'b111111111;
assign micromatrizz[8][222] = 9'b111111111;
assign micromatrizz[8][223] = 9'b111111111;
assign micromatrizz[8][224] = 9'b111111111;
assign micromatrizz[8][225] = 9'b111111111;
assign micromatrizz[8][226] = 9'b111111111;
assign micromatrizz[8][227] = 9'b111111111;
assign micromatrizz[8][228] = 9'b111111111;
assign micromatrizz[8][229] = 9'b111111111;
assign micromatrizz[8][230] = 9'b111111111;
assign micromatrizz[8][231] = 9'b111111111;
assign micromatrizz[8][232] = 9'b111111111;
assign micromatrizz[8][233] = 9'b111111111;
assign micromatrizz[8][234] = 9'b111111111;
assign micromatrizz[8][235] = 9'b111111111;
assign micromatrizz[8][236] = 9'b111111111;
assign micromatrizz[8][237] = 9'b111111111;
assign micromatrizz[8][238] = 9'b111111111;
assign micromatrizz[8][239] = 9'b111111111;
assign micromatrizz[8][240] = 9'b111111111;
assign micromatrizz[8][241] = 9'b111111111;
assign micromatrizz[8][242] = 9'b111111111;
assign micromatrizz[8][243] = 9'b111111111;
assign micromatrizz[8][244] = 9'b111111111;
assign micromatrizz[8][245] = 9'b111111111;
assign micromatrizz[8][246] = 9'b111111111;
assign micromatrizz[8][247] = 9'b111111111;
assign micromatrizz[8][248] = 9'b111111111;
assign micromatrizz[8][249] = 9'b111111111;
assign micromatrizz[8][250] = 9'b111111111;
assign micromatrizz[8][251] = 9'b111111111;
assign micromatrizz[8][252] = 9'b111111111;
assign micromatrizz[8][253] = 9'b111111111;
assign micromatrizz[8][254] = 9'b111111111;
assign micromatrizz[8][255] = 9'b111111111;
assign micromatrizz[8][256] = 9'b111111111;
assign micromatrizz[8][257] = 9'b111111111;
assign micromatrizz[8][258] = 9'b111111111;
assign micromatrizz[8][259] = 9'b111111111;
assign micromatrizz[8][260] = 9'b111111111;
assign micromatrizz[8][261] = 9'b111111111;
assign micromatrizz[8][262] = 9'b111111111;
assign micromatrizz[8][263] = 9'b111111111;
assign micromatrizz[8][264] = 9'b111111111;
assign micromatrizz[8][265] = 9'b111111111;
assign micromatrizz[8][266] = 9'b111111111;
assign micromatrizz[8][267] = 9'b111111111;
assign micromatrizz[8][268] = 9'b111111111;
assign micromatrizz[8][269] = 9'b111111111;
assign micromatrizz[8][270] = 9'b111111111;
assign micromatrizz[8][271] = 9'b111111111;
assign micromatrizz[8][272] = 9'b111111111;
assign micromatrizz[8][273] = 9'b111111111;
assign micromatrizz[8][274] = 9'b111111111;
assign micromatrizz[8][275] = 9'b111111111;
assign micromatrizz[8][276] = 9'b111111111;
assign micromatrizz[8][277] = 9'b111111111;
assign micromatrizz[8][278] = 9'b111111111;
assign micromatrizz[8][279] = 9'b111111111;
assign micromatrizz[8][280] = 9'b111111111;
assign micromatrizz[8][281] = 9'b111111111;
assign micromatrizz[8][282] = 9'b111111111;
assign micromatrizz[8][283] = 9'b111111111;
assign micromatrizz[8][284] = 9'b111111111;
assign micromatrizz[8][285] = 9'b111111111;
assign micromatrizz[8][286] = 9'b111111111;
assign micromatrizz[8][287] = 9'b111111111;
assign micromatrizz[8][288] = 9'b111111111;
assign micromatrizz[8][289] = 9'b111111111;
assign micromatrizz[8][290] = 9'b111111111;
assign micromatrizz[8][291] = 9'b111111111;
assign micromatrizz[8][292] = 9'b111111111;
assign micromatrizz[8][293] = 9'b111111111;
assign micromatrizz[8][294] = 9'b111111111;
assign micromatrizz[8][295] = 9'b111111111;
assign micromatrizz[8][296] = 9'b111111111;
assign micromatrizz[8][297] = 9'b111111111;
assign micromatrizz[8][298] = 9'b111111111;
assign micromatrizz[8][299] = 9'b111111111;
assign micromatrizz[8][300] = 9'b111111111;
assign micromatrizz[8][301] = 9'b111111111;
assign micromatrizz[8][302] = 9'b111111111;
assign micromatrizz[8][303] = 9'b111111111;
assign micromatrizz[8][304] = 9'b111111111;
assign micromatrizz[8][305] = 9'b111111111;
assign micromatrizz[8][306] = 9'b111111111;
assign micromatrizz[8][307] = 9'b111111111;
assign micromatrizz[8][308] = 9'b111111111;
assign micromatrizz[8][309] = 9'b111111111;
assign micromatrizz[8][310] = 9'b111111111;
assign micromatrizz[8][311] = 9'b111111111;
assign micromatrizz[8][312] = 9'b111111111;
assign micromatrizz[8][313] = 9'b111111111;
assign micromatrizz[8][314] = 9'b111111111;
assign micromatrizz[8][315] = 9'b111111111;
assign micromatrizz[8][316] = 9'b111111111;
assign micromatrizz[8][317] = 9'b111111111;
assign micromatrizz[8][318] = 9'b111111111;
assign micromatrizz[8][319] = 9'b111111111;
assign micromatrizz[8][320] = 9'b111111111;
assign micromatrizz[8][321] = 9'b111111111;
assign micromatrizz[8][322] = 9'b111111111;
assign micromatrizz[8][323] = 9'b111111111;
assign micromatrizz[8][324] = 9'b111111111;
assign micromatrizz[8][325] = 9'b111111111;
assign micromatrizz[8][326] = 9'b111111111;
assign micromatrizz[8][327] = 9'b111111111;
assign micromatrizz[8][328] = 9'b111111111;
assign micromatrizz[8][329] = 9'b111111111;
assign micromatrizz[8][330] = 9'b111111111;
assign micromatrizz[8][331] = 9'b111111111;
assign micromatrizz[8][332] = 9'b111111111;
assign micromatrizz[8][333] = 9'b111111111;
assign micromatrizz[8][334] = 9'b111111111;
assign micromatrizz[8][335] = 9'b111111111;
assign micromatrizz[8][336] = 9'b111111111;
assign micromatrizz[8][337] = 9'b111111111;
assign micromatrizz[8][338] = 9'b111111111;
assign micromatrizz[8][339] = 9'b111111111;
assign micromatrizz[8][340] = 9'b111111111;
assign micromatrizz[8][341] = 9'b111111111;
assign micromatrizz[8][342] = 9'b111111111;
assign micromatrizz[8][343] = 9'b111111111;
assign micromatrizz[8][344] = 9'b111111111;
assign micromatrizz[8][345] = 9'b111111111;
assign micromatrizz[8][346] = 9'b111111111;
assign micromatrizz[8][347] = 9'b111111111;
assign micromatrizz[8][348] = 9'b111111111;
assign micromatrizz[8][349] = 9'b111111111;
assign micromatrizz[8][350] = 9'b111111111;
assign micromatrizz[8][351] = 9'b111111111;
assign micromatrizz[8][352] = 9'b111111111;
assign micromatrizz[8][353] = 9'b111111111;
assign micromatrizz[8][354] = 9'b111111111;
assign micromatrizz[8][355] = 9'b111111111;
assign micromatrizz[8][356] = 9'b111111111;
assign micromatrizz[8][357] = 9'b111111111;
assign micromatrizz[8][358] = 9'b111111111;
assign micromatrizz[8][359] = 9'b111111111;
assign micromatrizz[8][360] = 9'b111111111;
assign micromatrizz[8][361] = 9'b111111111;
assign micromatrizz[8][362] = 9'b111111111;
assign micromatrizz[8][363] = 9'b111111111;
assign micromatrizz[8][364] = 9'b111111111;
assign micromatrizz[8][365] = 9'b111111111;
assign micromatrizz[8][366] = 9'b111111111;
assign micromatrizz[8][367] = 9'b111111111;
assign micromatrizz[8][368] = 9'b111111111;
assign micromatrizz[8][369] = 9'b111111111;
assign micromatrizz[8][370] = 9'b111111111;
assign micromatrizz[8][371] = 9'b111111111;
assign micromatrizz[8][372] = 9'b111111111;
assign micromatrizz[8][373] = 9'b111111111;
assign micromatrizz[8][374] = 9'b111111111;
assign micromatrizz[8][375] = 9'b111111111;
assign micromatrizz[8][376] = 9'b111111111;
assign micromatrizz[8][377] = 9'b111111111;
assign micromatrizz[8][378] = 9'b111111111;
assign micromatrizz[8][379] = 9'b111111111;
assign micromatrizz[8][380] = 9'b111111111;
assign micromatrizz[8][381] = 9'b111111111;
assign micromatrizz[8][382] = 9'b111111111;
assign micromatrizz[8][383] = 9'b111111111;
assign micromatrizz[8][384] = 9'b111111111;
assign micromatrizz[8][385] = 9'b111111111;
assign micromatrizz[8][386] = 9'b111111111;
assign micromatrizz[8][387] = 9'b111111111;
assign micromatrizz[8][388] = 9'b111111111;
assign micromatrizz[8][389] = 9'b111111111;
assign micromatrizz[8][390] = 9'b111111111;
assign micromatrizz[8][391] = 9'b111111111;
assign micromatrizz[8][392] = 9'b111111111;
assign micromatrizz[8][393] = 9'b111111111;
assign micromatrizz[8][394] = 9'b111111111;
assign micromatrizz[8][395] = 9'b111111111;
assign micromatrizz[8][396] = 9'b111111111;
assign micromatrizz[8][397] = 9'b111111111;
assign micromatrizz[8][398] = 9'b111111111;
assign micromatrizz[8][399] = 9'b111111111;
assign micromatrizz[8][400] = 9'b111111111;
assign micromatrizz[8][401] = 9'b111111111;
assign micromatrizz[8][402] = 9'b111111111;
assign micromatrizz[8][403] = 9'b111111111;
assign micromatrizz[8][404] = 9'b111111111;
assign micromatrizz[8][405] = 9'b111111111;
assign micromatrizz[8][406] = 9'b111111111;
assign micromatrizz[8][407] = 9'b111111111;
assign micromatrizz[8][408] = 9'b111111111;
assign micromatrizz[8][409] = 9'b111111111;
assign micromatrizz[8][410] = 9'b111111111;
assign micromatrizz[8][411] = 9'b111111111;
assign micromatrizz[8][412] = 9'b111111111;
assign micromatrizz[8][413] = 9'b111111111;
assign micromatrizz[8][414] = 9'b111111111;
assign micromatrizz[8][415] = 9'b111111111;
assign micromatrizz[8][416] = 9'b111111111;
assign micromatrizz[8][417] = 9'b111111111;
assign micromatrizz[8][418] = 9'b111111111;
assign micromatrizz[8][419] = 9'b111111111;
assign micromatrizz[8][420] = 9'b111111111;
assign micromatrizz[8][421] = 9'b111111111;
assign micromatrizz[8][422] = 9'b111111111;
assign micromatrizz[8][423] = 9'b111111111;
assign micromatrizz[8][424] = 9'b111111111;
assign micromatrizz[8][425] = 9'b111111111;
assign micromatrizz[8][426] = 9'b111111111;
assign micromatrizz[8][427] = 9'b111111111;
assign micromatrizz[8][428] = 9'b111111111;
assign micromatrizz[8][429] = 9'b111111111;
assign micromatrizz[8][430] = 9'b111111111;
assign micromatrizz[8][431] = 9'b111111111;
assign micromatrizz[8][432] = 9'b111111111;
assign micromatrizz[8][433] = 9'b111111111;
assign micromatrizz[8][434] = 9'b111111111;
assign micromatrizz[8][435] = 9'b111111111;
assign micromatrizz[8][436] = 9'b111111111;
assign micromatrizz[8][437] = 9'b111111111;
assign micromatrizz[8][438] = 9'b111111111;
assign micromatrizz[8][439] = 9'b111111111;
assign micromatrizz[8][440] = 9'b111111111;
assign micromatrizz[8][441] = 9'b111111111;
assign micromatrizz[8][442] = 9'b111111111;
assign micromatrizz[8][443] = 9'b111111111;
assign micromatrizz[8][444] = 9'b111111111;
assign micromatrizz[8][445] = 9'b111111111;
assign micromatrizz[8][446] = 9'b111111111;
assign micromatrizz[8][447] = 9'b111111111;
assign micromatrizz[8][448] = 9'b111111111;
assign micromatrizz[8][449] = 9'b111111111;
assign micromatrizz[8][450] = 9'b111111111;
assign micromatrizz[8][451] = 9'b111111111;
assign micromatrizz[8][452] = 9'b111111111;
assign micromatrizz[8][453] = 9'b111111111;
assign micromatrizz[8][454] = 9'b111111111;
assign micromatrizz[8][455] = 9'b111111111;
assign micromatrizz[8][456] = 9'b111111111;
assign micromatrizz[8][457] = 9'b111111111;
assign micromatrizz[8][458] = 9'b111111111;
assign micromatrizz[8][459] = 9'b111111111;
assign micromatrizz[8][460] = 9'b111111111;
assign micromatrizz[8][461] = 9'b111111111;
assign micromatrizz[8][462] = 9'b111111111;
assign micromatrizz[8][463] = 9'b111111111;
assign micromatrizz[8][464] = 9'b111111111;
assign micromatrizz[8][465] = 9'b111111111;
assign micromatrizz[8][466] = 9'b111111111;
assign micromatrizz[8][467] = 9'b111111111;
assign micromatrizz[8][468] = 9'b111111111;
assign micromatrizz[8][469] = 9'b111111111;
assign micromatrizz[8][470] = 9'b111111111;
assign micromatrizz[8][471] = 9'b111111111;
assign micromatrizz[8][472] = 9'b111111111;
assign micromatrizz[8][473] = 9'b111111111;
assign micromatrizz[8][474] = 9'b111111111;
assign micromatrizz[8][475] = 9'b111111111;
assign micromatrizz[8][476] = 9'b111111111;
assign micromatrizz[8][477] = 9'b111111111;
assign micromatrizz[8][478] = 9'b111111111;
assign micromatrizz[8][479] = 9'b111111111;
assign micromatrizz[8][480] = 9'b111111111;
assign micromatrizz[8][481] = 9'b111111111;
assign micromatrizz[8][482] = 9'b111111111;
assign micromatrizz[8][483] = 9'b111111111;
assign micromatrizz[8][484] = 9'b111111111;
assign micromatrizz[8][485] = 9'b111111111;
assign micromatrizz[8][486] = 9'b111111111;
assign micromatrizz[8][487] = 9'b111111111;
assign micromatrizz[8][488] = 9'b111111111;
assign micromatrizz[8][489] = 9'b111111111;
assign micromatrizz[8][490] = 9'b111111111;
assign micromatrizz[8][491] = 9'b111111111;
assign micromatrizz[8][492] = 9'b111111111;
assign micromatrizz[8][493] = 9'b111111111;
assign micromatrizz[8][494] = 9'b111111111;
assign micromatrizz[8][495] = 9'b111111111;
assign micromatrizz[8][496] = 9'b111111111;
assign micromatrizz[8][497] = 9'b111111111;
assign micromatrizz[8][498] = 9'b111111111;
assign micromatrizz[8][499] = 9'b111111111;
assign micromatrizz[8][500] = 9'b111111111;
assign micromatrizz[8][501] = 9'b111111111;
assign micromatrizz[8][502] = 9'b111111111;
assign micromatrizz[8][503] = 9'b111111111;
assign micromatrizz[8][504] = 9'b111111111;
assign micromatrizz[8][505] = 9'b111111111;
assign micromatrizz[8][506] = 9'b111111111;
assign micromatrizz[8][507] = 9'b111111111;
assign micromatrizz[8][508] = 9'b111111111;
assign micromatrizz[8][509] = 9'b111111111;
assign micromatrizz[8][510] = 9'b111111111;
assign micromatrizz[8][511] = 9'b111111111;
assign micromatrizz[8][512] = 9'b111111111;
assign micromatrizz[8][513] = 9'b111111111;
assign micromatrizz[8][514] = 9'b111111111;
assign micromatrizz[8][515] = 9'b111111111;
assign micromatrizz[8][516] = 9'b111111111;
assign micromatrizz[8][517] = 9'b111111111;
assign micromatrizz[8][518] = 9'b111111111;
assign micromatrizz[8][519] = 9'b111111111;
assign micromatrizz[8][520] = 9'b111111111;
assign micromatrizz[8][521] = 9'b111111111;
assign micromatrizz[8][522] = 9'b111111111;
assign micromatrizz[8][523] = 9'b111111111;
assign micromatrizz[8][524] = 9'b111111111;
assign micromatrizz[8][525] = 9'b111111111;
assign micromatrizz[8][526] = 9'b111111111;
assign micromatrizz[8][527] = 9'b111111111;
assign micromatrizz[8][528] = 9'b111111111;
assign micromatrizz[8][529] = 9'b111111111;
assign micromatrizz[8][530] = 9'b111111111;
assign micromatrizz[8][531] = 9'b111111111;
assign micromatrizz[8][532] = 9'b111111111;
assign micromatrizz[8][533] = 9'b111111111;
assign micromatrizz[8][534] = 9'b111111111;
assign micromatrizz[8][535] = 9'b111111111;
assign micromatrizz[8][536] = 9'b111111111;
assign micromatrizz[8][537] = 9'b111111111;
assign micromatrizz[8][538] = 9'b111111111;
assign micromatrizz[8][539] = 9'b111111111;
assign micromatrizz[8][540] = 9'b111111111;
assign micromatrizz[8][541] = 9'b111111111;
assign micromatrizz[8][542] = 9'b111111111;
assign micromatrizz[8][543] = 9'b111111111;
assign micromatrizz[8][544] = 9'b111111111;
assign micromatrizz[8][545] = 9'b111111111;
assign micromatrizz[8][546] = 9'b111111111;
assign micromatrizz[8][547] = 9'b111111111;
assign micromatrizz[8][548] = 9'b111111111;
assign micromatrizz[8][549] = 9'b111111111;
assign micromatrizz[8][550] = 9'b111111111;
assign micromatrizz[8][551] = 9'b111111111;
assign micromatrizz[8][552] = 9'b111111111;
assign micromatrizz[8][553] = 9'b111111111;
assign micromatrizz[8][554] = 9'b111111111;
assign micromatrizz[8][555] = 9'b111111111;
assign micromatrizz[8][556] = 9'b111111111;
assign micromatrizz[8][557] = 9'b111111111;
assign micromatrizz[8][558] = 9'b111111111;
assign micromatrizz[8][559] = 9'b111111111;
assign micromatrizz[8][560] = 9'b111111111;
assign micromatrizz[8][561] = 9'b111111111;
assign micromatrizz[8][562] = 9'b111111111;
assign micromatrizz[8][563] = 9'b111111111;
assign micromatrizz[8][564] = 9'b111111111;
assign micromatrizz[8][565] = 9'b111111111;
assign micromatrizz[8][566] = 9'b111111111;
assign micromatrizz[8][567] = 9'b111111111;
assign micromatrizz[8][568] = 9'b111111111;
assign micromatrizz[8][569] = 9'b111111111;
assign micromatrizz[8][570] = 9'b111111111;
assign micromatrizz[8][571] = 9'b111111111;
assign micromatrizz[8][572] = 9'b111111111;
assign micromatrizz[8][573] = 9'b111111111;
assign micromatrizz[8][574] = 9'b111111111;
assign micromatrizz[8][575] = 9'b111111111;
assign micromatrizz[8][576] = 9'b111111111;
assign micromatrizz[8][577] = 9'b111111111;
assign micromatrizz[8][578] = 9'b111111111;
assign micromatrizz[8][579] = 9'b111111111;
assign micromatrizz[8][580] = 9'b111111111;
assign micromatrizz[8][581] = 9'b111111111;
assign micromatrizz[8][582] = 9'b111111111;
assign micromatrizz[8][583] = 9'b111111111;
assign micromatrizz[8][584] = 9'b111111111;
assign micromatrizz[8][585] = 9'b111111111;
assign micromatrizz[8][586] = 9'b111111111;
assign micromatrizz[8][587] = 9'b111111111;
assign micromatrizz[8][588] = 9'b111111111;
assign micromatrizz[8][589] = 9'b111111111;
assign micromatrizz[8][590] = 9'b111111111;
assign micromatrizz[8][591] = 9'b111111111;
assign micromatrizz[8][592] = 9'b111111111;
assign micromatrizz[8][593] = 9'b111111111;
assign micromatrizz[8][594] = 9'b111111111;
assign micromatrizz[8][595] = 9'b111111111;
assign micromatrizz[8][596] = 9'b111111111;
assign micromatrizz[8][597] = 9'b111111111;
assign micromatrizz[8][598] = 9'b111111111;
assign micromatrizz[8][599] = 9'b111111111;
assign micromatrizz[8][600] = 9'b111111111;
assign micromatrizz[8][601] = 9'b111111111;
assign micromatrizz[8][602] = 9'b111111111;
assign micromatrizz[8][603] = 9'b111111111;
assign micromatrizz[8][604] = 9'b111111111;
assign micromatrizz[8][605] = 9'b111111111;
assign micromatrizz[8][606] = 9'b111111111;
assign micromatrizz[8][607] = 9'b111111111;
assign micromatrizz[8][608] = 9'b111111111;
assign micromatrizz[8][609] = 9'b111111111;
assign micromatrizz[8][610] = 9'b111111111;
assign micromatrizz[8][611] = 9'b111111111;
assign micromatrizz[8][612] = 9'b111111111;
assign micromatrizz[8][613] = 9'b111111111;
assign micromatrizz[8][614] = 9'b111111111;
assign micromatrizz[8][615] = 9'b111111111;
assign micromatrizz[8][616] = 9'b111111111;
assign micromatrizz[8][617] = 9'b111111111;
assign micromatrizz[8][618] = 9'b111111111;
assign micromatrizz[8][619] = 9'b111111111;
assign micromatrizz[8][620] = 9'b111111111;
assign micromatrizz[8][621] = 9'b111111111;
assign micromatrizz[8][622] = 9'b111111111;
assign micromatrizz[8][623] = 9'b111111111;
assign micromatrizz[8][624] = 9'b111111111;
assign micromatrizz[8][625] = 9'b111111111;
assign micromatrizz[8][626] = 9'b111111111;
assign micromatrizz[8][627] = 9'b111111111;
assign micromatrizz[8][628] = 9'b111111111;
assign micromatrizz[8][629] = 9'b111111111;
assign micromatrizz[8][630] = 9'b111111111;
assign micromatrizz[8][631] = 9'b111111111;
assign micromatrizz[8][632] = 9'b111111111;
assign micromatrizz[8][633] = 9'b111111111;
assign micromatrizz[8][634] = 9'b111111111;
assign micromatrizz[8][635] = 9'b111111111;
assign micromatrizz[8][636] = 9'b111111111;
assign micromatrizz[8][637] = 9'b111111111;
assign micromatrizz[8][638] = 9'b111111111;
assign micromatrizz[8][639] = 9'b111111111;
assign micromatrizz[9][0] = 9'b111111111;
assign micromatrizz[9][1] = 9'b111111111;
assign micromatrizz[9][2] = 9'b111111111;
assign micromatrizz[9][3] = 9'b111111111;
assign micromatrizz[9][4] = 9'b111111111;
assign micromatrizz[9][5] = 9'b111111111;
assign micromatrizz[9][6] = 9'b111111111;
assign micromatrizz[9][7] = 9'b111111111;
assign micromatrizz[9][8] = 9'b111111111;
assign micromatrizz[9][9] = 9'b111111111;
assign micromatrizz[9][10] = 9'b111111111;
assign micromatrizz[9][11] = 9'b111111111;
assign micromatrizz[9][12] = 9'b111111111;
assign micromatrizz[9][13] = 9'b111111111;
assign micromatrizz[9][14] = 9'b111111111;
assign micromatrizz[9][15] = 9'b111111111;
assign micromatrizz[9][16] = 9'b111111111;
assign micromatrizz[9][17] = 9'b111111111;
assign micromatrizz[9][18] = 9'b111111111;
assign micromatrizz[9][19] = 9'b111111111;
assign micromatrizz[9][20] = 9'b111111111;
assign micromatrizz[9][21] = 9'b111111111;
assign micromatrizz[9][22] = 9'b111111111;
assign micromatrizz[9][23] = 9'b111111111;
assign micromatrizz[9][24] = 9'b111111111;
assign micromatrizz[9][25] = 9'b111111111;
assign micromatrizz[9][26] = 9'b111111111;
assign micromatrizz[9][27] = 9'b111111111;
assign micromatrizz[9][28] = 9'b111111111;
assign micromatrizz[9][29] = 9'b111111111;
assign micromatrizz[9][30] = 9'b111111111;
assign micromatrizz[9][31] = 9'b111111111;
assign micromatrizz[9][32] = 9'b111111111;
assign micromatrizz[9][33] = 9'b111111111;
assign micromatrizz[9][34] = 9'b111111111;
assign micromatrizz[9][35] = 9'b111111111;
assign micromatrizz[9][36] = 9'b111111111;
assign micromatrizz[9][37] = 9'b111111111;
assign micromatrizz[9][38] = 9'b111111111;
assign micromatrizz[9][39] = 9'b111111111;
assign micromatrizz[9][40] = 9'b111111111;
assign micromatrizz[9][41] = 9'b111111111;
assign micromatrizz[9][42] = 9'b111111111;
assign micromatrizz[9][43] = 9'b111111111;
assign micromatrizz[9][44] = 9'b111111111;
assign micromatrizz[9][45] = 9'b111111111;
assign micromatrizz[9][46] = 9'b111111111;
assign micromatrizz[9][47] = 9'b111111111;
assign micromatrizz[9][48] = 9'b111111111;
assign micromatrizz[9][49] = 9'b111111111;
assign micromatrizz[9][50] = 9'b111111111;
assign micromatrizz[9][51] = 9'b111111111;
assign micromatrizz[9][52] = 9'b111111111;
assign micromatrizz[9][53] = 9'b111111111;
assign micromatrizz[9][54] = 9'b111111111;
assign micromatrizz[9][55] = 9'b111111111;
assign micromatrizz[9][56] = 9'b111111111;
assign micromatrizz[9][57] = 9'b111111111;
assign micromatrizz[9][58] = 9'b111111111;
assign micromatrizz[9][59] = 9'b111111111;
assign micromatrizz[9][60] = 9'b111111111;
assign micromatrizz[9][61] = 9'b111111111;
assign micromatrizz[9][62] = 9'b111111111;
assign micromatrizz[9][63] = 9'b111111111;
assign micromatrizz[9][64] = 9'b111111111;
assign micromatrizz[9][65] = 9'b111111111;
assign micromatrizz[9][66] = 9'b111111111;
assign micromatrizz[9][67] = 9'b111111111;
assign micromatrizz[9][68] = 9'b111111111;
assign micromatrizz[9][69] = 9'b111111111;
assign micromatrizz[9][70] = 9'b111111111;
assign micromatrizz[9][71] = 9'b111111111;
assign micromatrizz[9][72] = 9'b111111111;
assign micromatrizz[9][73] = 9'b111111111;
assign micromatrizz[9][74] = 9'b111111111;
assign micromatrizz[9][75] = 9'b111111111;
assign micromatrizz[9][76] = 9'b111111111;
assign micromatrizz[9][77] = 9'b111111111;
assign micromatrizz[9][78] = 9'b111111111;
assign micromatrizz[9][79] = 9'b111111111;
assign micromatrizz[9][80] = 9'b111111111;
assign micromatrizz[9][81] = 9'b111111111;
assign micromatrizz[9][82] = 9'b111111111;
assign micromatrizz[9][83] = 9'b111111111;
assign micromatrizz[9][84] = 9'b111111111;
assign micromatrizz[9][85] = 9'b111111111;
assign micromatrizz[9][86] = 9'b111111111;
assign micromatrizz[9][87] = 9'b111111111;
assign micromatrizz[9][88] = 9'b111111111;
assign micromatrizz[9][89] = 9'b111111111;
assign micromatrizz[9][90] = 9'b111111111;
assign micromatrizz[9][91] = 9'b111111111;
assign micromatrizz[9][92] = 9'b111111111;
assign micromatrizz[9][93] = 9'b111111111;
assign micromatrizz[9][94] = 9'b111111111;
assign micromatrizz[9][95] = 9'b111111111;
assign micromatrizz[9][96] = 9'b111111111;
assign micromatrizz[9][97] = 9'b111111111;
assign micromatrizz[9][98] = 9'b111111111;
assign micromatrizz[9][99] = 9'b111111111;
assign micromatrizz[9][100] = 9'b111111111;
assign micromatrizz[9][101] = 9'b111111111;
assign micromatrizz[9][102] = 9'b111111111;
assign micromatrizz[9][103] = 9'b111111111;
assign micromatrizz[9][104] = 9'b111111111;
assign micromatrizz[9][105] = 9'b111111111;
assign micromatrizz[9][106] = 9'b111111111;
assign micromatrizz[9][107] = 9'b111111111;
assign micromatrizz[9][108] = 9'b111111111;
assign micromatrizz[9][109] = 9'b111111111;
assign micromatrizz[9][110] = 9'b111111111;
assign micromatrizz[9][111] = 9'b111111111;
assign micromatrizz[9][112] = 9'b111111111;
assign micromatrizz[9][113] = 9'b111111111;
assign micromatrizz[9][114] = 9'b111111111;
assign micromatrizz[9][115] = 9'b111111111;
assign micromatrizz[9][116] = 9'b111111111;
assign micromatrizz[9][117] = 9'b111111111;
assign micromatrizz[9][118] = 9'b111111111;
assign micromatrizz[9][119] = 9'b111111111;
assign micromatrizz[9][120] = 9'b111111111;
assign micromatrizz[9][121] = 9'b111111111;
assign micromatrizz[9][122] = 9'b111111111;
assign micromatrizz[9][123] = 9'b111111111;
assign micromatrizz[9][124] = 9'b111111111;
assign micromatrizz[9][125] = 9'b111111111;
assign micromatrizz[9][126] = 9'b111111111;
assign micromatrizz[9][127] = 9'b111111111;
assign micromatrizz[9][128] = 9'b111111111;
assign micromatrizz[9][129] = 9'b111111111;
assign micromatrizz[9][130] = 9'b111111111;
assign micromatrizz[9][131] = 9'b111111111;
assign micromatrizz[9][132] = 9'b111111111;
assign micromatrizz[9][133] = 9'b111111111;
assign micromatrizz[9][134] = 9'b111111111;
assign micromatrizz[9][135] = 9'b111111111;
assign micromatrizz[9][136] = 9'b111111111;
assign micromatrizz[9][137] = 9'b111111111;
assign micromatrizz[9][138] = 9'b111111111;
assign micromatrizz[9][139] = 9'b111111111;
assign micromatrizz[9][140] = 9'b111111111;
assign micromatrizz[9][141] = 9'b111111111;
assign micromatrizz[9][142] = 9'b111111111;
assign micromatrizz[9][143] = 9'b111111111;
assign micromatrizz[9][144] = 9'b111111111;
assign micromatrizz[9][145] = 9'b111111111;
assign micromatrizz[9][146] = 9'b111111111;
assign micromatrizz[9][147] = 9'b111111111;
assign micromatrizz[9][148] = 9'b111111111;
assign micromatrizz[9][149] = 9'b111111111;
assign micromatrizz[9][150] = 9'b111111111;
assign micromatrizz[9][151] = 9'b111111111;
assign micromatrizz[9][152] = 9'b111111111;
assign micromatrizz[9][153] = 9'b111111111;
assign micromatrizz[9][154] = 9'b111111111;
assign micromatrizz[9][155] = 9'b111111111;
assign micromatrizz[9][156] = 9'b111111111;
assign micromatrizz[9][157] = 9'b111111111;
assign micromatrizz[9][158] = 9'b111111111;
assign micromatrizz[9][159] = 9'b111111111;
assign micromatrizz[9][160] = 9'b111111111;
assign micromatrizz[9][161] = 9'b111111111;
assign micromatrizz[9][162] = 9'b111111111;
assign micromatrizz[9][163] = 9'b111111111;
assign micromatrizz[9][164] = 9'b111111111;
assign micromatrizz[9][165] = 9'b111111111;
assign micromatrizz[9][166] = 9'b111111111;
assign micromatrizz[9][167] = 9'b111111111;
assign micromatrizz[9][168] = 9'b111111111;
assign micromatrizz[9][169] = 9'b111111111;
assign micromatrizz[9][170] = 9'b111111111;
assign micromatrizz[9][171] = 9'b111111111;
assign micromatrizz[9][172] = 9'b111111111;
assign micromatrizz[9][173] = 9'b111111111;
assign micromatrizz[9][174] = 9'b111111111;
assign micromatrizz[9][175] = 9'b111111111;
assign micromatrizz[9][176] = 9'b111111111;
assign micromatrizz[9][177] = 9'b111111111;
assign micromatrizz[9][178] = 9'b111111111;
assign micromatrizz[9][179] = 9'b111111111;
assign micromatrizz[9][180] = 9'b111111111;
assign micromatrizz[9][181] = 9'b111111111;
assign micromatrizz[9][182] = 9'b111111111;
assign micromatrizz[9][183] = 9'b111111111;
assign micromatrizz[9][184] = 9'b111111111;
assign micromatrizz[9][185] = 9'b111111111;
assign micromatrizz[9][186] = 9'b111111111;
assign micromatrizz[9][187] = 9'b111111111;
assign micromatrizz[9][188] = 9'b111111111;
assign micromatrizz[9][189] = 9'b111111111;
assign micromatrizz[9][190] = 9'b111111111;
assign micromatrizz[9][191] = 9'b111111111;
assign micromatrizz[9][192] = 9'b111111111;
assign micromatrizz[9][193] = 9'b111111111;
assign micromatrizz[9][194] = 9'b111111111;
assign micromatrizz[9][195] = 9'b111111111;
assign micromatrizz[9][196] = 9'b111111111;
assign micromatrizz[9][197] = 9'b111111111;
assign micromatrizz[9][198] = 9'b111111111;
assign micromatrizz[9][199] = 9'b111111111;
assign micromatrizz[9][200] = 9'b111111111;
assign micromatrizz[9][201] = 9'b111111111;
assign micromatrizz[9][202] = 9'b111111111;
assign micromatrizz[9][203] = 9'b111111111;
assign micromatrizz[9][204] = 9'b111111111;
assign micromatrizz[9][205] = 9'b111111111;
assign micromatrizz[9][206] = 9'b111111111;
assign micromatrizz[9][207] = 9'b111111111;
assign micromatrizz[9][208] = 9'b111111111;
assign micromatrizz[9][209] = 9'b111111111;
assign micromatrizz[9][210] = 9'b111111111;
assign micromatrizz[9][211] = 9'b111111111;
assign micromatrizz[9][212] = 9'b111111111;
assign micromatrizz[9][213] = 9'b111111111;
assign micromatrizz[9][214] = 9'b111111111;
assign micromatrizz[9][215] = 9'b111111111;
assign micromatrizz[9][216] = 9'b111111111;
assign micromatrizz[9][217] = 9'b111111111;
assign micromatrizz[9][218] = 9'b111111111;
assign micromatrizz[9][219] = 9'b111111111;
assign micromatrizz[9][220] = 9'b111111111;
assign micromatrizz[9][221] = 9'b111111111;
assign micromatrizz[9][222] = 9'b111111111;
assign micromatrizz[9][223] = 9'b111111111;
assign micromatrizz[9][224] = 9'b111111111;
assign micromatrizz[9][225] = 9'b111111111;
assign micromatrizz[9][226] = 9'b111111111;
assign micromatrizz[9][227] = 9'b111111111;
assign micromatrizz[9][228] = 9'b111111111;
assign micromatrizz[9][229] = 9'b111111111;
assign micromatrizz[9][230] = 9'b111111111;
assign micromatrizz[9][231] = 9'b111111111;
assign micromatrizz[9][232] = 9'b111111111;
assign micromatrizz[9][233] = 9'b111111111;
assign micromatrizz[9][234] = 9'b111111111;
assign micromatrizz[9][235] = 9'b111111111;
assign micromatrizz[9][236] = 9'b111111111;
assign micromatrizz[9][237] = 9'b111111111;
assign micromatrizz[9][238] = 9'b111111111;
assign micromatrizz[9][239] = 9'b111111111;
assign micromatrizz[9][240] = 9'b111111111;
assign micromatrizz[9][241] = 9'b111111111;
assign micromatrizz[9][242] = 9'b111111111;
assign micromatrizz[9][243] = 9'b111111111;
assign micromatrizz[9][244] = 9'b111111111;
assign micromatrizz[9][245] = 9'b111111111;
assign micromatrizz[9][246] = 9'b111111111;
assign micromatrizz[9][247] = 9'b111111111;
assign micromatrizz[9][248] = 9'b111111111;
assign micromatrizz[9][249] = 9'b111111111;
assign micromatrizz[9][250] = 9'b111111111;
assign micromatrizz[9][251] = 9'b111111111;
assign micromatrizz[9][252] = 9'b111111111;
assign micromatrizz[9][253] = 9'b111111111;
assign micromatrizz[9][254] = 9'b111111111;
assign micromatrizz[9][255] = 9'b111111111;
assign micromatrizz[9][256] = 9'b111111111;
assign micromatrizz[9][257] = 9'b111111111;
assign micromatrizz[9][258] = 9'b111111111;
assign micromatrizz[9][259] = 9'b111111111;
assign micromatrizz[9][260] = 9'b111111111;
assign micromatrizz[9][261] = 9'b111111111;
assign micromatrizz[9][262] = 9'b111111111;
assign micromatrizz[9][263] = 9'b111111111;
assign micromatrizz[9][264] = 9'b111111111;
assign micromatrizz[9][265] = 9'b111111111;
assign micromatrizz[9][266] = 9'b111111111;
assign micromatrizz[9][267] = 9'b111111111;
assign micromatrizz[9][268] = 9'b111111111;
assign micromatrizz[9][269] = 9'b111111111;
assign micromatrizz[9][270] = 9'b111111111;
assign micromatrizz[9][271] = 9'b111111111;
assign micromatrizz[9][272] = 9'b111111111;
assign micromatrizz[9][273] = 9'b111111111;
assign micromatrizz[9][274] = 9'b111111111;
assign micromatrizz[9][275] = 9'b111111111;
assign micromatrizz[9][276] = 9'b111111111;
assign micromatrizz[9][277] = 9'b111111111;
assign micromatrizz[9][278] = 9'b111111111;
assign micromatrizz[9][279] = 9'b111111111;
assign micromatrizz[9][280] = 9'b111111111;
assign micromatrizz[9][281] = 9'b111111111;
assign micromatrizz[9][282] = 9'b111111111;
assign micromatrizz[9][283] = 9'b111111111;
assign micromatrizz[9][284] = 9'b111111111;
assign micromatrizz[9][285] = 9'b111111111;
assign micromatrizz[9][286] = 9'b111111111;
assign micromatrizz[9][287] = 9'b111111111;
assign micromatrizz[9][288] = 9'b111111111;
assign micromatrizz[9][289] = 9'b111111111;
assign micromatrizz[9][290] = 9'b111111111;
assign micromatrizz[9][291] = 9'b111111111;
assign micromatrizz[9][292] = 9'b111111111;
assign micromatrizz[9][293] = 9'b111111111;
assign micromatrizz[9][294] = 9'b111111111;
assign micromatrizz[9][295] = 9'b111111111;
assign micromatrizz[9][296] = 9'b111111111;
assign micromatrizz[9][297] = 9'b111111111;
assign micromatrizz[9][298] = 9'b111111111;
assign micromatrizz[9][299] = 9'b111111111;
assign micromatrizz[9][300] = 9'b111111111;
assign micromatrizz[9][301] = 9'b111111111;
assign micromatrizz[9][302] = 9'b111111111;
assign micromatrizz[9][303] = 9'b111111111;
assign micromatrizz[9][304] = 9'b111111111;
assign micromatrizz[9][305] = 9'b111111111;
assign micromatrizz[9][306] = 9'b111111111;
assign micromatrizz[9][307] = 9'b111111111;
assign micromatrizz[9][308] = 9'b111111111;
assign micromatrizz[9][309] = 9'b111111111;
assign micromatrizz[9][310] = 9'b111111111;
assign micromatrizz[9][311] = 9'b111111111;
assign micromatrizz[9][312] = 9'b111111111;
assign micromatrizz[9][313] = 9'b111111111;
assign micromatrizz[9][314] = 9'b111111111;
assign micromatrizz[9][315] = 9'b111111111;
assign micromatrizz[9][316] = 9'b111111111;
assign micromatrizz[9][317] = 9'b111111111;
assign micromatrizz[9][318] = 9'b111111111;
assign micromatrizz[9][319] = 9'b111111111;
assign micromatrizz[9][320] = 9'b111111111;
assign micromatrizz[9][321] = 9'b111111111;
assign micromatrizz[9][322] = 9'b111111111;
assign micromatrizz[9][323] = 9'b111111111;
assign micromatrizz[9][324] = 9'b111111111;
assign micromatrizz[9][325] = 9'b111111111;
assign micromatrizz[9][326] = 9'b111111111;
assign micromatrizz[9][327] = 9'b111111111;
assign micromatrizz[9][328] = 9'b111111111;
assign micromatrizz[9][329] = 9'b111111111;
assign micromatrizz[9][330] = 9'b111111111;
assign micromatrizz[9][331] = 9'b111111111;
assign micromatrizz[9][332] = 9'b111111111;
assign micromatrizz[9][333] = 9'b111111111;
assign micromatrizz[9][334] = 9'b111111111;
assign micromatrizz[9][335] = 9'b111111111;
assign micromatrizz[9][336] = 9'b111111111;
assign micromatrizz[9][337] = 9'b111111111;
assign micromatrizz[9][338] = 9'b111111111;
assign micromatrizz[9][339] = 9'b111111111;
assign micromatrizz[9][340] = 9'b111111111;
assign micromatrizz[9][341] = 9'b111111111;
assign micromatrizz[9][342] = 9'b111111111;
assign micromatrizz[9][343] = 9'b111111111;
assign micromatrizz[9][344] = 9'b111111111;
assign micromatrizz[9][345] = 9'b111111111;
assign micromatrizz[9][346] = 9'b111111111;
assign micromatrizz[9][347] = 9'b111111111;
assign micromatrizz[9][348] = 9'b111111111;
assign micromatrizz[9][349] = 9'b111111111;
assign micromatrizz[9][350] = 9'b111111111;
assign micromatrizz[9][351] = 9'b111111111;
assign micromatrizz[9][352] = 9'b111111111;
assign micromatrizz[9][353] = 9'b111111111;
assign micromatrizz[9][354] = 9'b111111111;
assign micromatrizz[9][355] = 9'b111111111;
assign micromatrizz[9][356] = 9'b111111111;
assign micromatrizz[9][357] = 9'b111111111;
assign micromatrizz[9][358] = 9'b111111111;
assign micromatrizz[9][359] = 9'b111111111;
assign micromatrizz[9][360] = 9'b111111111;
assign micromatrizz[9][361] = 9'b111111111;
assign micromatrizz[9][362] = 9'b111111111;
assign micromatrizz[9][363] = 9'b111111111;
assign micromatrizz[9][364] = 9'b111111111;
assign micromatrizz[9][365] = 9'b111111111;
assign micromatrizz[9][366] = 9'b111111111;
assign micromatrizz[9][367] = 9'b111111111;
assign micromatrizz[9][368] = 9'b111111111;
assign micromatrizz[9][369] = 9'b111111111;
assign micromatrizz[9][370] = 9'b111111111;
assign micromatrizz[9][371] = 9'b111111111;
assign micromatrizz[9][372] = 9'b111111111;
assign micromatrizz[9][373] = 9'b111111111;
assign micromatrizz[9][374] = 9'b111111111;
assign micromatrizz[9][375] = 9'b111111111;
assign micromatrizz[9][376] = 9'b111111111;
assign micromatrizz[9][377] = 9'b111111111;
assign micromatrizz[9][378] = 9'b111111111;
assign micromatrizz[9][379] = 9'b111111111;
assign micromatrizz[9][380] = 9'b111111111;
assign micromatrizz[9][381] = 9'b111111111;
assign micromatrizz[9][382] = 9'b111111111;
assign micromatrizz[9][383] = 9'b111111111;
assign micromatrizz[9][384] = 9'b111111111;
assign micromatrizz[9][385] = 9'b111111111;
assign micromatrizz[9][386] = 9'b111111111;
assign micromatrizz[9][387] = 9'b111111111;
assign micromatrizz[9][388] = 9'b111111111;
assign micromatrizz[9][389] = 9'b111111111;
assign micromatrizz[9][390] = 9'b111111111;
assign micromatrizz[9][391] = 9'b111111111;
assign micromatrizz[9][392] = 9'b111111111;
assign micromatrizz[9][393] = 9'b111111111;
assign micromatrizz[9][394] = 9'b111111111;
assign micromatrizz[9][395] = 9'b111111111;
assign micromatrizz[9][396] = 9'b111111111;
assign micromatrizz[9][397] = 9'b111111111;
assign micromatrizz[9][398] = 9'b111111111;
assign micromatrizz[9][399] = 9'b111111111;
assign micromatrizz[9][400] = 9'b111111111;
assign micromatrizz[9][401] = 9'b111111111;
assign micromatrizz[9][402] = 9'b111111111;
assign micromatrizz[9][403] = 9'b111111111;
assign micromatrizz[9][404] = 9'b111111111;
assign micromatrizz[9][405] = 9'b111111111;
assign micromatrizz[9][406] = 9'b111111111;
assign micromatrizz[9][407] = 9'b111111111;
assign micromatrizz[9][408] = 9'b111111111;
assign micromatrizz[9][409] = 9'b111111111;
assign micromatrizz[9][410] = 9'b111111111;
assign micromatrizz[9][411] = 9'b111111111;
assign micromatrizz[9][412] = 9'b111111111;
assign micromatrizz[9][413] = 9'b111111111;
assign micromatrizz[9][414] = 9'b111111111;
assign micromatrizz[9][415] = 9'b111111111;
assign micromatrizz[9][416] = 9'b111111111;
assign micromatrizz[9][417] = 9'b111111111;
assign micromatrizz[9][418] = 9'b111111111;
assign micromatrizz[9][419] = 9'b111111111;
assign micromatrizz[9][420] = 9'b111111111;
assign micromatrizz[9][421] = 9'b111111111;
assign micromatrizz[9][422] = 9'b111111111;
assign micromatrizz[9][423] = 9'b111111111;
assign micromatrizz[9][424] = 9'b111111111;
assign micromatrizz[9][425] = 9'b111111111;
assign micromatrizz[9][426] = 9'b111111111;
assign micromatrizz[9][427] = 9'b111111111;
assign micromatrizz[9][428] = 9'b111111111;
assign micromatrizz[9][429] = 9'b111111111;
assign micromatrizz[9][430] = 9'b111111111;
assign micromatrizz[9][431] = 9'b111111111;
assign micromatrizz[9][432] = 9'b111111111;
assign micromatrizz[9][433] = 9'b111111111;
assign micromatrizz[9][434] = 9'b111111111;
assign micromatrizz[9][435] = 9'b111111111;
assign micromatrizz[9][436] = 9'b111111111;
assign micromatrizz[9][437] = 9'b111111111;
assign micromatrizz[9][438] = 9'b111111111;
assign micromatrizz[9][439] = 9'b111111111;
assign micromatrizz[9][440] = 9'b111111111;
assign micromatrizz[9][441] = 9'b111111111;
assign micromatrizz[9][442] = 9'b111111111;
assign micromatrizz[9][443] = 9'b111111111;
assign micromatrizz[9][444] = 9'b111111111;
assign micromatrizz[9][445] = 9'b111111111;
assign micromatrizz[9][446] = 9'b111111111;
assign micromatrizz[9][447] = 9'b111111111;
assign micromatrizz[9][448] = 9'b111111111;
assign micromatrizz[9][449] = 9'b111111111;
assign micromatrizz[9][450] = 9'b111111111;
assign micromatrizz[9][451] = 9'b111111111;
assign micromatrizz[9][452] = 9'b111111111;
assign micromatrizz[9][453] = 9'b111111111;
assign micromatrizz[9][454] = 9'b111111111;
assign micromatrizz[9][455] = 9'b111111111;
assign micromatrizz[9][456] = 9'b111111111;
assign micromatrizz[9][457] = 9'b111111111;
assign micromatrizz[9][458] = 9'b111111111;
assign micromatrizz[9][459] = 9'b111111111;
assign micromatrizz[9][460] = 9'b111111111;
assign micromatrizz[9][461] = 9'b111111111;
assign micromatrizz[9][462] = 9'b111111111;
assign micromatrizz[9][463] = 9'b111111111;
assign micromatrizz[9][464] = 9'b111111111;
assign micromatrizz[9][465] = 9'b111111111;
assign micromatrizz[9][466] = 9'b111111111;
assign micromatrizz[9][467] = 9'b111111111;
assign micromatrizz[9][468] = 9'b111111111;
assign micromatrizz[9][469] = 9'b111111111;
assign micromatrizz[9][470] = 9'b111111111;
assign micromatrizz[9][471] = 9'b111111111;
assign micromatrizz[9][472] = 9'b111111111;
assign micromatrizz[9][473] = 9'b111111111;
assign micromatrizz[9][474] = 9'b111111111;
assign micromatrizz[9][475] = 9'b111111111;
assign micromatrizz[9][476] = 9'b111111111;
assign micromatrizz[9][477] = 9'b111111111;
assign micromatrizz[9][478] = 9'b111111111;
assign micromatrizz[9][479] = 9'b111111111;
assign micromatrizz[9][480] = 9'b111111111;
assign micromatrizz[9][481] = 9'b111111111;
assign micromatrizz[9][482] = 9'b111111111;
assign micromatrizz[9][483] = 9'b111111111;
assign micromatrizz[9][484] = 9'b111111111;
assign micromatrizz[9][485] = 9'b111111111;
assign micromatrizz[9][486] = 9'b111111111;
assign micromatrizz[9][487] = 9'b111111111;
assign micromatrizz[9][488] = 9'b111111111;
assign micromatrizz[9][489] = 9'b111111111;
assign micromatrizz[9][490] = 9'b111111111;
assign micromatrizz[9][491] = 9'b111111111;
assign micromatrizz[9][492] = 9'b111111111;
assign micromatrizz[9][493] = 9'b111111111;
assign micromatrizz[9][494] = 9'b111111111;
assign micromatrizz[9][495] = 9'b111111111;
assign micromatrizz[9][496] = 9'b111111111;
assign micromatrizz[9][497] = 9'b111111111;
assign micromatrizz[9][498] = 9'b111111111;
assign micromatrizz[9][499] = 9'b111111111;
assign micromatrizz[9][500] = 9'b111111111;
assign micromatrizz[9][501] = 9'b111111111;
assign micromatrizz[9][502] = 9'b111111111;
assign micromatrizz[9][503] = 9'b111111111;
assign micromatrizz[9][504] = 9'b111111111;
assign micromatrizz[9][505] = 9'b111111111;
assign micromatrizz[9][506] = 9'b111111111;
assign micromatrizz[9][507] = 9'b111111111;
assign micromatrizz[9][508] = 9'b111111111;
assign micromatrizz[9][509] = 9'b111111111;
assign micromatrizz[9][510] = 9'b111111111;
assign micromatrizz[9][511] = 9'b111111111;
assign micromatrizz[9][512] = 9'b111111111;
assign micromatrizz[9][513] = 9'b111111111;
assign micromatrizz[9][514] = 9'b111111111;
assign micromatrizz[9][515] = 9'b111111111;
assign micromatrizz[9][516] = 9'b111111111;
assign micromatrizz[9][517] = 9'b111111111;
assign micromatrizz[9][518] = 9'b111111111;
assign micromatrizz[9][519] = 9'b111111111;
assign micromatrizz[9][520] = 9'b111111111;
assign micromatrizz[9][521] = 9'b111111111;
assign micromatrizz[9][522] = 9'b111111111;
assign micromatrizz[9][523] = 9'b111111111;
assign micromatrizz[9][524] = 9'b111111111;
assign micromatrizz[9][525] = 9'b111111111;
assign micromatrizz[9][526] = 9'b111111111;
assign micromatrizz[9][527] = 9'b111111111;
assign micromatrizz[9][528] = 9'b111111111;
assign micromatrizz[9][529] = 9'b111111111;
assign micromatrizz[9][530] = 9'b111111111;
assign micromatrizz[9][531] = 9'b111111111;
assign micromatrizz[9][532] = 9'b111111111;
assign micromatrizz[9][533] = 9'b111111111;
assign micromatrizz[9][534] = 9'b111111111;
assign micromatrizz[9][535] = 9'b111111111;
assign micromatrizz[9][536] = 9'b111111111;
assign micromatrizz[9][537] = 9'b111111111;
assign micromatrizz[9][538] = 9'b111111111;
assign micromatrizz[9][539] = 9'b111111111;
assign micromatrizz[9][540] = 9'b111111111;
assign micromatrizz[9][541] = 9'b111111111;
assign micromatrizz[9][542] = 9'b111111111;
assign micromatrizz[9][543] = 9'b111111111;
assign micromatrizz[9][544] = 9'b111111111;
assign micromatrizz[9][545] = 9'b111111111;
assign micromatrizz[9][546] = 9'b111111111;
assign micromatrizz[9][547] = 9'b111111111;
assign micromatrizz[9][548] = 9'b111111111;
assign micromatrizz[9][549] = 9'b111111111;
assign micromatrizz[9][550] = 9'b111111111;
assign micromatrizz[9][551] = 9'b111111111;
assign micromatrizz[9][552] = 9'b111111111;
assign micromatrizz[9][553] = 9'b111111111;
assign micromatrizz[9][554] = 9'b111111111;
assign micromatrizz[9][555] = 9'b111111111;
assign micromatrizz[9][556] = 9'b111111111;
assign micromatrizz[9][557] = 9'b111111111;
assign micromatrizz[9][558] = 9'b111111111;
assign micromatrizz[9][559] = 9'b111111111;
assign micromatrizz[9][560] = 9'b111111111;
assign micromatrizz[9][561] = 9'b111111111;
assign micromatrizz[9][562] = 9'b111111111;
assign micromatrizz[9][563] = 9'b111111111;
assign micromatrizz[9][564] = 9'b111111111;
assign micromatrizz[9][565] = 9'b111111111;
assign micromatrizz[9][566] = 9'b111111111;
assign micromatrizz[9][567] = 9'b111111111;
assign micromatrizz[9][568] = 9'b111111111;
assign micromatrizz[9][569] = 9'b111111111;
assign micromatrizz[9][570] = 9'b111111111;
assign micromatrizz[9][571] = 9'b111111111;
assign micromatrizz[9][572] = 9'b111111111;
assign micromatrizz[9][573] = 9'b111111111;
assign micromatrizz[9][574] = 9'b111111111;
assign micromatrizz[9][575] = 9'b111111111;
assign micromatrizz[9][576] = 9'b111111111;
assign micromatrizz[9][577] = 9'b111111111;
assign micromatrizz[9][578] = 9'b111111111;
assign micromatrizz[9][579] = 9'b111111111;
assign micromatrizz[9][580] = 9'b111111111;
assign micromatrizz[9][581] = 9'b111111111;
assign micromatrizz[9][582] = 9'b111111111;
assign micromatrizz[9][583] = 9'b111111111;
assign micromatrizz[9][584] = 9'b111111111;
assign micromatrizz[9][585] = 9'b111111111;
assign micromatrizz[9][586] = 9'b111111111;
assign micromatrizz[9][587] = 9'b111111111;
assign micromatrizz[9][588] = 9'b111111111;
assign micromatrizz[9][589] = 9'b111111111;
assign micromatrizz[9][590] = 9'b111111111;
assign micromatrizz[9][591] = 9'b111111111;
assign micromatrizz[9][592] = 9'b111111111;
assign micromatrizz[9][593] = 9'b111111111;
assign micromatrizz[9][594] = 9'b111111111;
assign micromatrizz[9][595] = 9'b111111111;
assign micromatrizz[9][596] = 9'b111111111;
assign micromatrizz[9][597] = 9'b111111111;
assign micromatrizz[9][598] = 9'b111111111;
assign micromatrizz[9][599] = 9'b111111111;
assign micromatrizz[9][600] = 9'b111111111;
assign micromatrizz[9][601] = 9'b111111111;
assign micromatrizz[9][602] = 9'b111111111;
assign micromatrizz[9][603] = 9'b111111111;
assign micromatrizz[9][604] = 9'b111111111;
assign micromatrizz[9][605] = 9'b111111111;
assign micromatrizz[9][606] = 9'b111111111;
assign micromatrizz[9][607] = 9'b111111111;
assign micromatrizz[9][608] = 9'b111111111;
assign micromatrizz[9][609] = 9'b111111111;
assign micromatrizz[9][610] = 9'b111111111;
assign micromatrizz[9][611] = 9'b111111111;
assign micromatrizz[9][612] = 9'b111111111;
assign micromatrizz[9][613] = 9'b111111111;
assign micromatrizz[9][614] = 9'b111111111;
assign micromatrizz[9][615] = 9'b111111111;
assign micromatrizz[9][616] = 9'b111111111;
assign micromatrizz[9][617] = 9'b111111111;
assign micromatrizz[9][618] = 9'b111111111;
assign micromatrizz[9][619] = 9'b111111111;
assign micromatrizz[9][620] = 9'b111111111;
assign micromatrizz[9][621] = 9'b111111111;
assign micromatrizz[9][622] = 9'b111111111;
assign micromatrizz[9][623] = 9'b111111111;
assign micromatrizz[9][624] = 9'b111111111;
assign micromatrizz[9][625] = 9'b111111111;
assign micromatrizz[9][626] = 9'b111111111;
assign micromatrizz[9][627] = 9'b111111111;
assign micromatrizz[9][628] = 9'b111111111;
assign micromatrizz[9][629] = 9'b111111111;
assign micromatrizz[9][630] = 9'b111111111;
assign micromatrizz[9][631] = 9'b111111111;
assign micromatrizz[9][632] = 9'b111111111;
assign micromatrizz[9][633] = 9'b111111111;
assign micromatrizz[9][634] = 9'b111111111;
assign micromatrizz[9][635] = 9'b111111111;
assign micromatrizz[9][636] = 9'b111111111;
assign micromatrizz[9][637] = 9'b111111111;
assign micromatrizz[9][638] = 9'b111111111;
assign micromatrizz[9][639] = 9'b111111111;
assign micromatrizz[10][0] = 9'b111111111;
assign micromatrizz[10][1] = 9'b111111111;
assign micromatrizz[10][2] = 9'b111111111;
assign micromatrizz[10][3] = 9'b111111111;
assign micromatrizz[10][4] = 9'b111111111;
assign micromatrizz[10][5] = 9'b111111111;
assign micromatrizz[10][6] = 9'b111111111;
assign micromatrizz[10][7] = 9'b111111111;
assign micromatrizz[10][8] = 9'b111111111;
assign micromatrizz[10][9] = 9'b111111111;
assign micromatrizz[10][10] = 9'b111111111;
assign micromatrizz[10][11] = 9'b111111111;
assign micromatrizz[10][12] = 9'b111111111;
assign micromatrizz[10][13] = 9'b111111111;
assign micromatrizz[10][14] = 9'b111111111;
assign micromatrizz[10][15] = 9'b111111111;
assign micromatrizz[10][16] = 9'b111111111;
assign micromatrizz[10][17] = 9'b111111111;
assign micromatrizz[10][18] = 9'b111111111;
assign micromatrizz[10][19] = 9'b111111111;
assign micromatrizz[10][20] = 9'b111111111;
assign micromatrizz[10][21] = 9'b111111111;
assign micromatrizz[10][22] = 9'b111111111;
assign micromatrizz[10][23] = 9'b111111111;
assign micromatrizz[10][24] = 9'b111111111;
assign micromatrizz[10][25] = 9'b111111111;
assign micromatrizz[10][26] = 9'b111111111;
assign micromatrizz[10][27] = 9'b111111111;
assign micromatrizz[10][28] = 9'b111111111;
assign micromatrizz[10][29] = 9'b111111111;
assign micromatrizz[10][30] = 9'b111111111;
assign micromatrizz[10][31] = 9'b111111111;
assign micromatrizz[10][32] = 9'b111111111;
assign micromatrizz[10][33] = 9'b111111111;
assign micromatrizz[10][34] = 9'b111111111;
assign micromatrizz[10][35] = 9'b111111111;
assign micromatrizz[10][36] = 9'b111111111;
assign micromatrizz[10][37] = 9'b111111111;
assign micromatrizz[10][38] = 9'b111111111;
assign micromatrizz[10][39] = 9'b111111111;
assign micromatrizz[10][40] = 9'b111111111;
assign micromatrizz[10][41] = 9'b111111111;
assign micromatrizz[10][42] = 9'b111111111;
assign micromatrizz[10][43] = 9'b111111111;
assign micromatrizz[10][44] = 9'b111111111;
assign micromatrizz[10][45] = 9'b111111111;
assign micromatrizz[10][46] = 9'b111111111;
assign micromatrizz[10][47] = 9'b111111111;
assign micromatrizz[10][48] = 9'b111111111;
assign micromatrizz[10][49] = 9'b111111111;
assign micromatrizz[10][50] = 9'b111111111;
assign micromatrizz[10][51] = 9'b111111111;
assign micromatrizz[10][52] = 9'b111111111;
assign micromatrizz[10][53] = 9'b111111111;
assign micromatrizz[10][54] = 9'b111111111;
assign micromatrizz[10][55] = 9'b111111111;
assign micromatrizz[10][56] = 9'b111111111;
assign micromatrizz[10][57] = 9'b111111111;
assign micromatrizz[10][58] = 9'b111111111;
assign micromatrizz[10][59] = 9'b111111111;
assign micromatrizz[10][60] = 9'b111111111;
assign micromatrizz[10][61] = 9'b111111111;
assign micromatrizz[10][62] = 9'b111111111;
assign micromatrizz[10][63] = 9'b111111111;
assign micromatrizz[10][64] = 9'b111111111;
assign micromatrizz[10][65] = 9'b111111111;
assign micromatrizz[10][66] = 9'b111111111;
assign micromatrizz[10][67] = 9'b111111111;
assign micromatrizz[10][68] = 9'b111111111;
assign micromatrizz[10][69] = 9'b111111111;
assign micromatrizz[10][70] = 9'b111111111;
assign micromatrizz[10][71] = 9'b111111111;
assign micromatrizz[10][72] = 9'b111111111;
assign micromatrizz[10][73] = 9'b111111111;
assign micromatrizz[10][74] = 9'b111111111;
assign micromatrizz[10][75] = 9'b111111111;
assign micromatrizz[10][76] = 9'b111111111;
assign micromatrizz[10][77] = 9'b111111111;
assign micromatrizz[10][78] = 9'b111111111;
assign micromatrizz[10][79] = 9'b111111111;
assign micromatrizz[10][80] = 9'b111111111;
assign micromatrizz[10][81] = 9'b111111111;
assign micromatrizz[10][82] = 9'b111111111;
assign micromatrizz[10][83] = 9'b111111111;
assign micromatrizz[10][84] = 9'b111111111;
assign micromatrizz[10][85] = 9'b111111111;
assign micromatrizz[10][86] = 9'b111111111;
assign micromatrizz[10][87] = 9'b111111111;
assign micromatrizz[10][88] = 9'b111111111;
assign micromatrizz[10][89] = 9'b111111111;
assign micromatrizz[10][90] = 9'b111111111;
assign micromatrizz[10][91] = 9'b111111111;
assign micromatrizz[10][92] = 9'b111111111;
assign micromatrizz[10][93] = 9'b111111111;
assign micromatrizz[10][94] = 9'b111111111;
assign micromatrizz[10][95] = 9'b111111111;
assign micromatrizz[10][96] = 9'b111111111;
assign micromatrizz[10][97] = 9'b111111111;
assign micromatrizz[10][98] = 9'b111111111;
assign micromatrizz[10][99] = 9'b111111111;
assign micromatrizz[10][100] = 9'b111111111;
assign micromatrizz[10][101] = 9'b111111111;
assign micromatrizz[10][102] = 9'b111111111;
assign micromatrizz[10][103] = 9'b111111111;
assign micromatrizz[10][104] = 9'b111111111;
assign micromatrizz[10][105] = 9'b111111111;
assign micromatrizz[10][106] = 9'b111111111;
assign micromatrizz[10][107] = 9'b111111111;
assign micromatrizz[10][108] = 9'b111111111;
assign micromatrizz[10][109] = 9'b111111111;
assign micromatrizz[10][110] = 9'b111111111;
assign micromatrizz[10][111] = 9'b111111111;
assign micromatrizz[10][112] = 9'b111111111;
assign micromatrizz[10][113] = 9'b111111111;
assign micromatrizz[10][114] = 9'b111111111;
assign micromatrizz[10][115] = 9'b111111111;
assign micromatrizz[10][116] = 9'b111111111;
assign micromatrizz[10][117] = 9'b111111111;
assign micromatrizz[10][118] = 9'b111111111;
assign micromatrizz[10][119] = 9'b111111111;
assign micromatrizz[10][120] = 9'b111111111;
assign micromatrizz[10][121] = 9'b111111111;
assign micromatrizz[10][122] = 9'b111111111;
assign micromatrizz[10][123] = 9'b111111111;
assign micromatrizz[10][124] = 9'b111111111;
assign micromatrizz[10][125] = 9'b111111111;
assign micromatrizz[10][126] = 9'b111111111;
assign micromatrizz[10][127] = 9'b111111111;
assign micromatrizz[10][128] = 9'b111111111;
assign micromatrizz[10][129] = 9'b111111111;
assign micromatrizz[10][130] = 9'b111111111;
assign micromatrizz[10][131] = 9'b111111111;
assign micromatrizz[10][132] = 9'b111111111;
assign micromatrizz[10][133] = 9'b111111111;
assign micromatrizz[10][134] = 9'b111111111;
assign micromatrizz[10][135] = 9'b111111111;
assign micromatrizz[10][136] = 9'b111111111;
assign micromatrizz[10][137] = 9'b111111111;
assign micromatrizz[10][138] = 9'b111111111;
assign micromatrizz[10][139] = 9'b111111111;
assign micromatrizz[10][140] = 9'b111111111;
assign micromatrizz[10][141] = 9'b111111111;
assign micromatrizz[10][142] = 9'b111111111;
assign micromatrizz[10][143] = 9'b111111111;
assign micromatrizz[10][144] = 9'b111111111;
assign micromatrizz[10][145] = 9'b111111111;
assign micromatrizz[10][146] = 9'b111111111;
assign micromatrizz[10][147] = 9'b111111111;
assign micromatrizz[10][148] = 9'b111111111;
assign micromatrizz[10][149] = 9'b111111111;
assign micromatrizz[10][150] = 9'b111111111;
assign micromatrizz[10][151] = 9'b111111111;
assign micromatrizz[10][152] = 9'b111111111;
assign micromatrizz[10][153] = 9'b111111111;
assign micromatrizz[10][154] = 9'b111111111;
assign micromatrizz[10][155] = 9'b111111111;
assign micromatrizz[10][156] = 9'b111111111;
assign micromatrizz[10][157] = 9'b111111111;
assign micromatrizz[10][158] = 9'b111111111;
assign micromatrizz[10][159] = 9'b111111111;
assign micromatrizz[10][160] = 9'b111111111;
assign micromatrizz[10][161] = 9'b111111111;
assign micromatrizz[10][162] = 9'b111111111;
assign micromatrizz[10][163] = 9'b111111111;
assign micromatrizz[10][164] = 9'b111111111;
assign micromatrizz[10][165] = 9'b111111111;
assign micromatrizz[10][166] = 9'b111111111;
assign micromatrizz[10][167] = 9'b111111111;
assign micromatrizz[10][168] = 9'b111111111;
assign micromatrizz[10][169] = 9'b111111111;
assign micromatrizz[10][170] = 9'b111111111;
assign micromatrizz[10][171] = 9'b111111111;
assign micromatrizz[10][172] = 9'b111111111;
assign micromatrizz[10][173] = 9'b111111111;
assign micromatrizz[10][174] = 9'b111111111;
assign micromatrizz[10][175] = 9'b111111111;
assign micromatrizz[10][176] = 9'b111111111;
assign micromatrizz[10][177] = 9'b111111111;
assign micromatrizz[10][178] = 9'b111111111;
assign micromatrizz[10][179] = 9'b111111111;
assign micromatrizz[10][180] = 9'b111111111;
assign micromatrizz[10][181] = 9'b111111111;
assign micromatrizz[10][182] = 9'b111111111;
assign micromatrizz[10][183] = 9'b111111111;
assign micromatrizz[10][184] = 9'b111111111;
assign micromatrizz[10][185] = 9'b111111111;
assign micromatrizz[10][186] = 9'b111111111;
assign micromatrizz[10][187] = 9'b111111111;
assign micromatrizz[10][188] = 9'b111111111;
assign micromatrizz[10][189] = 9'b111111111;
assign micromatrizz[10][190] = 9'b111111111;
assign micromatrizz[10][191] = 9'b111111111;
assign micromatrizz[10][192] = 9'b111111111;
assign micromatrizz[10][193] = 9'b111111111;
assign micromatrizz[10][194] = 9'b111111111;
assign micromatrizz[10][195] = 9'b111111111;
assign micromatrizz[10][196] = 9'b111111111;
assign micromatrizz[10][197] = 9'b111111111;
assign micromatrizz[10][198] = 9'b111111111;
assign micromatrizz[10][199] = 9'b111111111;
assign micromatrizz[10][200] = 9'b111111111;
assign micromatrizz[10][201] = 9'b111111111;
assign micromatrizz[10][202] = 9'b111111111;
assign micromatrizz[10][203] = 9'b111111111;
assign micromatrizz[10][204] = 9'b111111111;
assign micromatrizz[10][205] = 9'b111111111;
assign micromatrizz[10][206] = 9'b111111111;
assign micromatrizz[10][207] = 9'b111111111;
assign micromatrizz[10][208] = 9'b111111111;
assign micromatrizz[10][209] = 9'b111111111;
assign micromatrizz[10][210] = 9'b111111111;
assign micromatrizz[10][211] = 9'b111111111;
assign micromatrizz[10][212] = 9'b111111111;
assign micromatrizz[10][213] = 9'b111111111;
assign micromatrizz[10][214] = 9'b111111111;
assign micromatrizz[10][215] = 9'b111111111;
assign micromatrizz[10][216] = 9'b111111111;
assign micromatrizz[10][217] = 9'b111111111;
assign micromatrizz[10][218] = 9'b111111111;
assign micromatrizz[10][219] = 9'b111111111;
assign micromatrizz[10][220] = 9'b111111111;
assign micromatrizz[10][221] = 9'b111111111;
assign micromatrizz[10][222] = 9'b111111111;
assign micromatrizz[10][223] = 9'b111111111;
assign micromatrizz[10][224] = 9'b111111111;
assign micromatrizz[10][225] = 9'b111111111;
assign micromatrizz[10][226] = 9'b111111111;
assign micromatrizz[10][227] = 9'b111111111;
assign micromatrizz[10][228] = 9'b111111111;
assign micromatrizz[10][229] = 9'b111111111;
assign micromatrizz[10][230] = 9'b111111111;
assign micromatrizz[10][231] = 9'b111111111;
assign micromatrizz[10][232] = 9'b111111111;
assign micromatrizz[10][233] = 9'b111111111;
assign micromatrizz[10][234] = 9'b111111111;
assign micromatrizz[10][235] = 9'b111111111;
assign micromatrizz[10][236] = 9'b111111111;
assign micromatrizz[10][237] = 9'b111111111;
assign micromatrizz[10][238] = 9'b111111111;
assign micromatrizz[10][239] = 9'b111111111;
assign micromatrizz[10][240] = 9'b111111111;
assign micromatrizz[10][241] = 9'b111111111;
assign micromatrizz[10][242] = 9'b111111111;
assign micromatrizz[10][243] = 9'b111111111;
assign micromatrizz[10][244] = 9'b111111111;
assign micromatrizz[10][245] = 9'b111111111;
assign micromatrizz[10][246] = 9'b111111111;
assign micromatrizz[10][247] = 9'b111111111;
assign micromatrizz[10][248] = 9'b111111111;
assign micromatrizz[10][249] = 9'b111111111;
assign micromatrizz[10][250] = 9'b111111111;
assign micromatrizz[10][251] = 9'b111111111;
assign micromatrizz[10][252] = 9'b111111111;
assign micromatrizz[10][253] = 9'b111111111;
assign micromatrizz[10][254] = 9'b111111111;
assign micromatrizz[10][255] = 9'b111111111;
assign micromatrizz[10][256] = 9'b111111111;
assign micromatrizz[10][257] = 9'b111111111;
assign micromatrizz[10][258] = 9'b111111111;
assign micromatrizz[10][259] = 9'b111111111;
assign micromatrizz[10][260] = 9'b111111111;
assign micromatrizz[10][261] = 9'b111111111;
assign micromatrizz[10][262] = 9'b111111111;
assign micromatrizz[10][263] = 9'b111111111;
assign micromatrizz[10][264] = 9'b111111111;
assign micromatrizz[10][265] = 9'b111111111;
assign micromatrizz[10][266] = 9'b111111111;
assign micromatrizz[10][267] = 9'b111111111;
assign micromatrizz[10][268] = 9'b111111111;
assign micromatrizz[10][269] = 9'b111111111;
assign micromatrizz[10][270] = 9'b111111111;
assign micromatrizz[10][271] = 9'b111111111;
assign micromatrizz[10][272] = 9'b111111111;
assign micromatrizz[10][273] = 9'b111111111;
assign micromatrizz[10][274] = 9'b111111111;
assign micromatrizz[10][275] = 9'b111111111;
assign micromatrizz[10][276] = 9'b111111111;
assign micromatrizz[10][277] = 9'b111111111;
assign micromatrizz[10][278] = 9'b111111111;
assign micromatrizz[10][279] = 9'b111111111;
assign micromatrizz[10][280] = 9'b111111111;
assign micromatrizz[10][281] = 9'b111111111;
assign micromatrizz[10][282] = 9'b111111111;
assign micromatrizz[10][283] = 9'b111111111;
assign micromatrizz[10][284] = 9'b111111111;
assign micromatrizz[10][285] = 9'b111111111;
assign micromatrizz[10][286] = 9'b111111111;
assign micromatrizz[10][287] = 9'b111111111;
assign micromatrizz[10][288] = 9'b111111111;
assign micromatrizz[10][289] = 9'b111111111;
assign micromatrizz[10][290] = 9'b111111111;
assign micromatrizz[10][291] = 9'b111111111;
assign micromatrizz[10][292] = 9'b111111111;
assign micromatrizz[10][293] = 9'b111111111;
assign micromatrizz[10][294] = 9'b111111111;
assign micromatrizz[10][295] = 9'b111111111;
assign micromatrizz[10][296] = 9'b111111111;
assign micromatrizz[10][297] = 9'b111111111;
assign micromatrizz[10][298] = 9'b111111111;
assign micromatrizz[10][299] = 9'b111111111;
assign micromatrizz[10][300] = 9'b111111111;
assign micromatrizz[10][301] = 9'b111111111;
assign micromatrizz[10][302] = 9'b111111111;
assign micromatrizz[10][303] = 9'b111111111;
assign micromatrizz[10][304] = 9'b111111111;
assign micromatrizz[10][305] = 9'b111111111;
assign micromatrizz[10][306] = 9'b111111111;
assign micromatrizz[10][307] = 9'b111111111;
assign micromatrizz[10][308] = 9'b111111111;
assign micromatrizz[10][309] = 9'b111111111;
assign micromatrizz[10][310] = 9'b111111111;
assign micromatrizz[10][311] = 9'b111111111;
assign micromatrizz[10][312] = 9'b111111111;
assign micromatrizz[10][313] = 9'b111111111;
assign micromatrizz[10][314] = 9'b111111111;
assign micromatrizz[10][315] = 9'b111111111;
assign micromatrizz[10][316] = 9'b111111111;
assign micromatrizz[10][317] = 9'b111111111;
assign micromatrizz[10][318] = 9'b111111111;
assign micromatrizz[10][319] = 9'b111111111;
assign micromatrizz[10][320] = 9'b111111111;
assign micromatrizz[10][321] = 9'b111111111;
assign micromatrizz[10][322] = 9'b111111111;
assign micromatrizz[10][323] = 9'b111111111;
assign micromatrizz[10][324] = 9'b111111111;
assign micromatrizz[10][325] = 9'b111111111;
assign micromatrizz[10][326] = 9'b111111111;
assign micromatrizz[10][327] = 9'b111111111;
assign micromatrizz[10][328] = 9'b111111111;
assign micromatrizz[10][329] = 9'b111111111;
assign micromatrizz[10][330] = 9'b111111111;
assign micromatrizz[10][331] = 9'b111111111;
assign micromatrizz[10][332] = 9'b111111111;
assign micromatrizz[10][333] = 9'b111111111;
assign micromatrizz[10][334] = 9'b111111111;
assign micromatrizz[10][335] = 9'b111111111;
assign micromatrizz[10][336] = 9'b111111111;
assign micromatrizz[10][337] = 9'b111111111;
assign micromatrizz[10][338] = 9'b111111111;
assign micromatrizz[10][339] = 9'b111111111;
assign micromatrizz[10][340] = 9'b111111111;
assign micromatrizz[10][341] = 9'b111111111;
assign micromatrizz[10][342] = 9'b111111111;
assign micromatrizz[10][343] = 9'b111111111;
assign micromatrizz[10][344] = 9'b111111111;
assign micromatrizz[10][345] = 9'b111111111;
assign micromatrizz[10][346] = 9'b111111111;
assign micromatrizz[10][347] = 9'b111111111;
assign micromatrizz[10][348] = 9'b111111111;
assign micromatrizz[10][349] = 9'b111111111;
assign micromatrizz[10][350] = 9'b111111111;
assign micromatrizz[10][351] = 9'b111111111;
assign micromatrizz[10][352] = 9'b111111111;
assign micromatrizz[10][353] = 9'b111111111;
assign micromatrizz[10][354] = 9'b111111111;
assign micromatrizz[10][355] = 9'b111111111;
assign micromatrizz[10][356] = 9'b111111111;
assign micromatrizz[10][357] = 9'b111111111;
assign micromatrizz[10][358] = 9'b111111111;
assign micromatrizz[10][359] = 9'b111111111;
assign micromatrizz[10][360] = 9'b111111111;
assign micromatrizz[10][361] = 9'b111111111;
assign micromatrizz[10][362] = 9'b111111111;
assign micromatrizz[10][363] = 9'b111111111;
assign micromatrizz[10][364] = 9'b111111111;
assign micromatrizz[10][365] = 9'b111111111;
assign micromatrizz[10][366] = 9'b111111111;
assign micromatrizz[10][367] = 9'b111111111;
assign micromatrizz[10][368] = 9'b111111111;
assign micromatrizz[10][369] = 9'b111111111;
assign micromatrizz[10][370] = 9'b111111111;
assign micromatrizz[10][371] = 9'b111111111;
assign micromatrizz[10][372] = 9'b111111111;
assign micromatrizz[10][373] = 9'b111111111;
assign micromatrizz[10][374] = 9'b111111111;
assign micromatrizz[10][375] = 9'b111111111;
assign micromatrizz[10][376] = 9'b111111111;
assign micromatrizz[10][377] = 9'b111111111;
assign micromatrizz[10][378] = 9'b111111111;
assign micromatrizz[10][379] = 9'b111111111;
assign micromatrizz[10][380] = 9'b111111111;
assign micromatrizz[10][381] = 9'b111111111;
assign micromatrizz[10][382] = 9'b111111111;
assign micromatrizz[10][383] = 9'b111111111;
assign micromatrizz[10][384] = 9'b111111111;
assign micromatrizz[10][385] = 9'b111111111;
assign micromatrizz[10][386] = 9'b111111111;
assign micromatrizz[10][387] = 9'b111111111;
assign micromatrizz[10][388] = 9'b111111111;
assign micromatrizz[10][389] = 9'b111111111;
assign micromatrizz[10][390] = 9'b111111111;
assign micromatrizz[10][391] = 9'b111111111;
assign micromatrizz[10][392] = 9'b111111111;
assign micromatrizz[10][393] = 9'b111111111;
assign micromatrizz[10][394] = 9'b111111111;
assign micromatrizz[10][395] = 9'b111111111;
assign micromatrizz[10][396] = 9'b111111111;
assign micromatrizz[10][397] = 9'b111111111;
assign micromatrizz[10][398] = 9'b111111111;
assign micromatrizz[10][399] = 9'b111111111;
assign micromatrizz[10][400] = 9'b111111111;
assign micromatrizz[10][401] = 9'b111111111;
assign micromatrizz[10][402] = 9'b111111111;
assign micromatrizz[10][403] = 9'b111111111;
assign micromatrizz[10][404] = 9'b111111111;
assign micromatrizz[10][405] = 9'b111111111;
assign micromatrizz[10][406] = 9'b111111111;
assign micromatrizz[10][407] = 9'b111111111;
assign micromatrizz[10][408] = 9'b111111111;
assign micromatrizz[10][409] = 9'b111111111;
assign micromatrizz[10][410] = 9'b111111111;
assign micromatrizz[10][411] = 9'b111111111;
assign micromatrizz[10][412] = 9'b111111111;
assign micromatrizz[10][413] = 9'b111111111;
assign micromatrizz[10][414] = 9'b111111111;
assign micromatrizz[10][415] = 9'b111111111;
assign micromatrizz[10][416] = 9'b111111111;
assign micromatrizz[10][417] = 9'b111111111;
assign micromatrizz[10][418] = 9'b111111111;
assign micromatrizz[10][419] = 9'b111111111;
assign micromatrizz[10][420] = 9'b111111111;
assign micromatrizz[10][421] = 9'b111111111;
assign micromatrizz[10][422] = 9'b111111111;
assign micromatrizz[10][423] = 9'b111111111;
assign micromatrizz[10][424] = 9'b111111111;
assign micromatrizz[10][425] = 9'b111111111;
assign micromatrizz[10][426] = 9'b111111111;
assign micromatrizz[10][427] = 9'b111111111;
assign micromatrizz[10][428] = 9'b111111111;
assign micromatrizz[10][429] = 9'b111111111;
assign micromatrizz[10][430] = 9'b111111111;
assign micromatrizz[10][431] = 9'b111111111;
assign micromatrizz[10][432] = 9'b111111111;
assign micromatrizz[10][433] = 9'b111111111;
assign micromatrizz[10][434] = 9'b111111111;
assign micromatrizz[10][435] = 9'b111111111;
assign micromatrizz[10][436] = 9'b111111111;
assign micromatrizz[10][437] = 9'b111111111;
assign micromatrizz[10][438] = 9'b111111111;
assign micromatrizz[10][439] = 9'b111111111;
assign micromatrizz[10][440] = 9'b111111111;
assign micromatrizz[10][441] = 9'b111111111;
assign micromatrizz[10][442] = 9'b111111111;
assign micromatrizz[10][443] = 9'b111111111;
assign micromatrizz[10][444] = 9'b111111111;
assign micromatrizz[10][445] = 9'b111111111;
assign micromatrizz[10][446] = 9'b111111111;
assign micromatrizz[10][447] = 9'b111111111;
assign micromatrizz[10][448] = 9'b111111111;
assign micromatrizz[10][449] = 9'b111111111;
assign micromatrizz[10][450] = 9'b111111111;
assign micromatrizz[10][451] = 9'b111111111;
assign micromatrizz[10][452] = 9'b111111111;
assign micromatrizz[10][453] = 9'b111111111;
assign micromatrizz[10][454] = 9'b111111111;
assign micromatrizz[10][455] = 9'b111111111;
assign micromatrizz[10][456] = 9'b111111111;
assign micromatrizz[10][457] = 9'b111111111;
assign micromatrizz[10][458] = 9'b111111111;
assign micromatrizz[10][459] = 9'b111111111;
assign micromatrizz[10][460] = 9'b111111111;
assign micromatrizz[10][461] = 9'b111111111;
assign micromatrizz[10][462] = 9'b111111111;
assign micromatrizz[10][463] = 9'b111111111;
assign micromatrizz[10][464] = 9'b111111111;
assign micromatrizz[10][465] = 9'b111111111;
assign micromatrizz[10][466] = 9'b111111111;
assign micromatrizz[10][467] = 9'b111111111;
assign micromatrizz[10][468] = 9'b111111111;
assign micromatrizz[10][469] = 9'b111111111;
assign micromatrizz[10][470] = 9'b111111111;
assign micromatrizz[10][471] = 9'b111111111;
assign micromatrizz[10][472] = 9'b111111111;
assign micromatrizz[10][473] = 9'b111111111;
assign micromatrizz[10][474] = 9'b111111111;
assign micromatrizz[10][475] = 9'b111111111;
assign micromatrizz[10][476] = 9'b111111111;
assign micromatrizz[10][477] = 9'b111111111;
assign micromatrizz[10][478] = 9'b111111111;
assign micromatrizz[10][479] = 9'b111111111;
assign micromatrizz[10][480] = 9'b111111111;
assign micromatrizz[10][481] = 9'b111111111;
assign micromatrizz[10][482] = 9'b111111111;
assign micromatrizz[10][483] = 9'b111111111;
assign micromatrizz[10][484] = 9'b111111111;
assign micromatrizz[10][485] = 9'b111111111;
assign micromatrizz[10][486] = 9'b111111111;
assign micromatrizz[10][487] = 9'b111111111;
assign micromatrizz[10][488] = 9'b111111111;
assign micromatrizz[10][489] = 9'b111111111;
assign micromatrizz[10][490] = 9'b111111111;
assign micromatrizz[10][491] = 9'b111111111;
assign micromatrizz[10][492] = 9'b111111111;
assign micromatrizz[10][493] = 9'b111111111;
assign micromatrizz[10][494] = 9'b111111111;
assign micromatrizz[10][495] = 9'b111111111;
assign micromatrizz[10][496] = 9'b111111111;
assign micromatrizz[10][497] = 9'b111111111;
assign micromatrizz[10][498] = 9'b111111111;
assign micromatrizz[10][499] = 9'b111111111;
assign micromatrizz[10][500] = 9'b111111111;
assign micromatrizz[10][501] = 9'b111111111;
assign micromatrizz[10][502] = 9'b111111111;
assign micromatrizz[10][503] = 9'b111111111;
assign micromatrizz[10][504] = 9'b111111111;
assign micromatrizz[10][505] = 9'b111111111;
assign micromatrizz[10][506] = 9'b111111111;
assign micromatrizz[10][507] = 9'b111111111;
assign micromatrizz[10][508] = 9'b111111111;
assign micromatrizz[10][509] = 9'b111111111;
assign micromatrizz[10][510] = 9'b111111111;
assign micromatrizz[10][511] = 9'b111111111;
assign micromatrizz[10][512] = 9'b111111111;
assign micromatrizz[10][513] = 9'b111111111;
assign micromatrizz[10][514] = 9'b111111111;
assign micromatrizz[10][515] = 9'b111111111;
assign micromatrizz[10][516] = 9'b111111111;
assign micromatrizz[10][517] = 9'b111111111;
assign micromatrizz[10][518] = 9'b111111111;
assign micromatrizz[10][519] = 9'b111111111;
assign micromatrizz[10][520] = 9'b111111111;
assign micromatrizz[10][521] = 9'b111111111;
assign micromatrizz[10][522] = 9'b111111111;
assign micromatrizz[10][523] = 9'b111111111;
assign micromatrizz[10][524] = 9'b111111111;
assign micromatrizz[10][525] = 9'b111111111;
assign micromatrizz[10][526] = 9'b111111111;
assign micromatrizz[10][527] = 9'b111111111;
assign micromatrizz[10][528] = 9'b111111111;
assign micromatrizz[10][529] = 9'b111111111;
assign micromatrizz[10][530] = 9'b111111111;
assign micromatrizz[10][531] = 9'b111111111;
assign micromatrizz[10][532] = 9'b111111111;
assign micromatrizz[10][533] = 9'b111111111;
assign micromatrizz[10][534] = 9'b111111111;
assign micromatrizz[10][535] = 9'b111111111;
assign micromatrizz[10][536] = 9'b111111111;
assign micromatrizz[10][537] = 9'b111111111;
assign micromatrizz[10][538] = 9'b111111111;
assign micromatrizz[10][539] = 9'b111111111;
assign micromatrizz[10][540] = 9'b111111111;
assign micromatrizz[10][541] = 9'b111111111;
assign micromatrizz[10][542] = 9'b111111111;
assign micromatrizz[10][543] = 9'b111111111;
assign micromatrizz[10][544] = 9'b111111111;
assign micromatrizz[10][545] = 9'b111111111;
assign micromatrizz[10][546] = 9'b111111111;
assign micromatrizz[10][547] = 9'b111111111;
assign micromatrizz[10][548] = 9'b111111111;
assign micromatrizz[10][549] = 9'b111111111;
assign micromatrizz[10][550] = 9'b111111111;
assign micromatrizz[10][551] = 9'b111111111;
assign micromatrizz[10][552] = 9'b111111111;
assign micromatrizz[10][553] = 9'b111111111;
assign micromatrizz[10][554] = 9'b111111111;
assign micromatrizz[10][555] = 9'b111111111;
assign micromatrizz[10][556] = 9'b111111111;
assign micromatrizz[10][557] = 9'b111111111;
assign micromatrizz[10][558] = 9'b111111111;
assign micromatrizz[10][559] = 9'b111111111;
assign micromatrizz[10][560] = 9'b111111111;
assign micromatrizz[10][561] = 9'b111111111;
assign micromatrizz[10][562] = 9'b111111111;
assign micromatrizz[10][563] = 9'b111111111;
assign micromatrizz[10][564] = 9'b111111111;
assign micromatrizz[10][565] = 9'b111111111;
assign micromatrizz[10][566] = 9'b111111111;
assign micromatrizz[10][567] = 9'b111111111;
assign micromatrizz[10][568] = 9'b111111111;
assign micromatrizz[10][569] = 9'b111111111;
assign micromatrizz[10][570] = 9'b111111111;
assign micromatrizz[10][571] = 9'b111111111;
assign micromatrizz[10][572] = 9'b111111111;
assign micromatrizz[10][573] = 9'b111111111;
assign micromatrizz[10][574] = 9'b111111111;
assign micromatrizz[10][575] = 9'b111111111;
assign micromatrizz[10][576] = 9'b111111111;
assign micromatrizz[10][577] = 9'b111111111;
assign micromatrizz[10][578] = 9'b111111111;
assign micromatrizz[10][579] = 9'b111111111;
assign micromatrizz[10][580] = 9'b111111111;
assign micromatrizz[10][581] = 9'b111111111;
assign micromatrizz[10][582] = 9'b111111111;
assign micromatrizz[10][583] = 9'b111111111;
assign micromatrizz[10][584] = 9'b111111111;
assign micromatrizz[10][585] = 9'b111111111;
assign micromatrizz[10][586] = 9'b111111111;
assign micromatrizz[10][587] = 9'b111111111;
assign micromatrizz[10][588] = 9'b111111111;
assign micromatrizz[10][589] = 9'b111111111;
assign micromatrizz[10][590] = 9'b111111111;
assign micromatrizz[10][591] = 9'b111111111;
assign micromatrizz[10][592] = 9'b111111111;
assign micromatrizz[10][593] = 9'b111111111;
assign micromatrizz[10][594] = 9'b111111111;
assign micromatrizz[10][595] = 9'b111111111;
assign micromatrizz[10][596] = 9'b111111111;
assign micromatrizz[10][597] = 9'b111111111;
assign micromatrizz[10][598] = 9'b111111111;
assign micromatrizz[10][599] = 9'b111111111;
assign micromatrizz[10][600] = 9'b111111111;
assign micromatrizz[10][601] = 9'b111111111;
assign micromatrizz[10][602] = 9'b111111111;
assign micromatrizz[10][603] = 9'b111111111;
assign micromatrizz[10][604] = 9'b111111111;
assign micromatrizz[10][605] = 9'b111111111;
assign micromatrizz[10][606] = 9'b111111111;
assign micromatrizz[10][607] = 9'b111111111;
assign micromatrizz[10][608] = 9'b111111111;
assign micromatrizz[10][609] = 9'b111111111;
assign micromatrizz[10][610] = 9'b111111111;
assign micromatrizz[10][611] = 9'b111111111;
assign micromatrizz[10][612] = 9'b111111111;
assign micromatrizz[10][613] = 9'b111111111;
assign micromatrizz[10][614] = 9'b111111111;
assign micromatrizz[10][615] = 9'b111111111;
assign micromatrizz[10][616] = 9'b111111111;
assign micromatrizz[10][617] = 9'b111111111;
assign micromatrizz[10][618] = 9'b111111111;
assign micromatrizz[10][619] = 9'b111111111;
assign micromatrizz[10][620] = 9'b111111111;
assign micromatrizz[10][621] = 9'b111111111;
assign micromatrizz[10][622] = 9'b111111111;
assign micromatrizz[10][623] = 9'b111111111;
assign micromatrizz[10][624] = 9'b111111111;
assign micromatrizz[10][625] = 9'b111111111;
assign micromatrizz[10][626] = 9'b111111111;
assign micromatrizz[10][627] = 9'b111111111;
assign micromatrizz[10][628] = 9'b111111111;
assign micromatrizz[10][629] = 9'b111111111;
assign micromatrizz[10][630] = 9'b111111111;
assign micromatrizz[10][631] = 9'b111111111;
assign micromatrizz[10][632] = 9'b111111111;
assign micromatrizz[10][633] = 9'b111111111;
assign micromatrizz[10][634] = 9'b111111111;
assign micromatrizz[10][635] = 9'b111111111;
assign micromatrizz[10][636] = 9'b111111111;
assign micromatrizz[10][637] = 9'b111111111;
assign micromatrizz[10][638] = 9'b111111111;
assign micromatrizz[10][639] = 9'b111111111;
assign micromatrizz[11][0] = 9'b111111111;
assign micromatrizz[11][1] = 9'b111111111;
assign micromatrizz[11][2] = 9'b111111111;
assign micromatrizz[11][3] = 9'b111111111;
assign micromatrizz[11][4] = 9'b111111111;
assign micromatrizz[11][5] = 9'b111111111;
assign micromatrizz[11][6] = 9'b111111111;
assign micromatrizz[11][7] = 9'b111111111;
assign micromatrizz[11][8] = 9'b111111111;
assign micromatrizz[11][9] = 9'b111111111;
assign micromatrizz[11][10] = 9'b111111111;
assign micromatrizz[11][11] = 9'b111111111;
assign micromatrizz[11][12] = 9'b111111111;
assign micromatrizz[11][13] = 9'b111111111;
assign micromatrizz[11][14] = 9'b111111111;
assign micromatrizz[11][15] = 9'b111111111;
assign micromatrizz[11][16] = 9'b111111111;
assign micromatrizz[11][17] = 9'b111111111;
assign micromatrizz[11][18] = 9'b111111111;
assign micromatrizz[11][19] = 9'b111111111;
assign micromatrizz[11][20] = 9'b111111111;
assign micromatrizz[11][21] = 9'b111111111;
assign micromatrizz[11][22] = 9'b111111111;
assign micromatrizz[11][23] = 9'b111111111;
assign micromatrizz[11][24] = 9'b111111111;
assign micromatrizz[11][25] = 9'b111111111;
assign micromatrizz[11][26] = 9'b111111111;
assign micromatrizz[11][27] = 9'b111111111;
assign micromatrizz[11][28] = 9'b111111111;
assign micromatrizz[11][29] = 9'b111111111;
assign micromatrizz[11][30] = 9'b111111111;
assign micromatrizz[11][31] = 9'b111111111;
assign micromatrizz[11][32] = 9'b111111111;
assign micromatrizz[11][33] = 9'b111111111;
assign micromatrizz[11][34] = 9'b111111111;
assign micromatrizz[11][35] = 9'b111111111;
assign micromatrizz[11][36] = 9'b111111111;
assign micromatrizz[11][37] = 9'b111111111;
assign micromatrizz[11][38] = 9'b111111111;
assign micromatrizz[11][39] = 9'b111111111;
assign micromatrizz[11][40] = 9'b111111111;
assign micromatrizz[11][41] = 9'b111111111;
assign micromatrizz[11][42] = 9'b111111111;
assign micromatrizz[11][43] = 9'b111111111;
assign micromatrizz[11][44] = 9'b111111111;
assign micromatrizz[11][45] = 9'b111111111;
assign micromatrizz[11][46] = 9'b111111111;
assign micromatrizz[11][47] = 9'b111111111;
assign micromatrizz[11][48] = 9'b111111111;
assign micromatrizz[11][49] = 9'b111111111;
assign micromatrizz[11][50] = 9'b111111111;
assign micromatrizz[11][51] = 9'b111111111;
assign micromatrizz[11][52] = 9'b111111111;
assign micromatrizz[11][53] = 9'b111111111;
assign micromatrizz[11][54] = 9'b111111111;
assign micromatrizz[11][55] = 9'b111111111;
assign micromatrizz[11][56] = 9'b111111111;
assign micromatrizz[11][57] = 9'b111111111;
assign micromatrizz[11][58] = 9'b111111111;
assign micromatrizz[11][59] = 9'b111111111;
assign micromatrizz[11][60] = 9'b111111111;
assign micromatrizz[11][61] = 9'b111111111;
assign micromatrizz[11][62] = 9'b111111111;
assign micromatrizz[11][63] = 9'b111111111;
assign micromatrizz[11][64] = 9'b111111111;
assign micromatrizz[11][65] = 9'b111111111;
assign micromatrizz[11][66] = 9'b111111111;
assign micromatrizz[11][67] = 9'b111111111;
assign micromatrizz[11][68] = 9'b111111111;
assign micromatrizz[11][69] = 9'b111111111;
assign micromatrizz[11][70] = 9'b111111111;
assign micromatrizz[11][71] = 9'b111111111;
assign micromatrizz[11][72] = 9'b111111111;
assign micromatrizz[11][73] = 9'b111111111;
assign micromatrizz[11][74] = 9'b111111111;
assign micromatrizz[11][75] = 9'b111111111;
assign micromatrizz[11][76] = 9'b111111111;
assign micromatrizz[11][77] = 9'b111111111;
assign micromatrizz[11][78] = 9'b111111111;
assign micromatrizz[11][79] = 9'b111111111;
assign micromatrizz[11][80] = 9'b111111111;
assign micromatrizz[11][81] = 9'b111111111;
assign micromatrizz[11][82] = 9'b111111111;
assign micromatrizz[11][83] = 9'b111111111;
assign micromatrizz[11][84] = 9'b111111111;
assign micromatrizz[11][85] = 9'b111111111;
assign micromatrizz[11][86] = 9'b111111111;
assign micromatrizz[11][87] = 9'b111111111;
assign micromatrizz[11][88] = 9'b111111111;
assign micromatrizz[11][89] = 9'b111111111;
assign micromatrizz[11][90] = 9'b111111111;
assign micromatrizz[11][91] = 9'b111111111;
assign micromatrizz[11][92] = 9'b111111111;
assign micromatrizz[11][93] = 9'b111111111;
assign micromatrizz[11][94] = 9'b111111111;
assign micromatrizz[11][95] = 9'b111111111;
assign micromatrizz[11][96] = 9'b111111111;
assign micromatrizz[11][97] = 9'b111111111;
assign micromatrizz[11][98] = 9'b111111111;
assign micromatrizz[11][99] = 9'b111111111;
assign micromatrizz[11][100] = 9'b111111111;
assign micromatrizz[11][101] = 9'b111111111;
assign micromatrizz[11][102] = 9'b111111111;
assign micromatrizz[11][103] = 9'b111111111;
assign micromatrizz[11][104] = 9'b111111111;
assign micromatrizz[11][105] = 9'b111111111;
assign micromatrizz[11][106] = 9'b111111111;
assign micromatrizz[11][107] = 9'b111111111;
assign micromatrizz[11][108] = 9'b111111111;
assign micromatrizz[11][109] = 9'b111111111;
assign micromatrizz[11][110] = 9'b111111111;
assign micromatrizz[11][111] = 9'b111111111;
assign micromatrizz[11][112] = 9'b111111111;
assign micromatrizz[11][113] = 9'b111111111;
assign micromatrizz[11][114] = 9'b111111111;
assign micromatrizz[11][115] = 9'b111111111;
assign micromatrizz[11][116] = 9'b111111111;
assign micromatrizz[11][117] = 9'b111111111;
assign micromatrizz[11][118] = 9'b111111111;
assign micromatrizz[11][119] = 9'b111111111;
assign micromatrizz[11][120] = 9'b111111111;
assign micromatrizz[11][121] = 9'b111111111;
assign micromatrizz[11][122] = 9'b111111111;
assign micromatrizz[11][123] = 9'b111111111;
assign micromatrizz[11][124] = 9'b111111111;
assign micromatrizz[11][125] = 9'b111111111;
assign micromatrizz[11][126] = 9'b111111111;
assign micromatrizz[11][127] = 9'b111111111;
assign micromatrizz[11][128] = 9'b111111111;
assign micromatrizz[11][129] = 9'b111111111;
assign micromatrizz[11][130] = 9'b111111111;
assign micromatrizz[11][131] = 9'b111111111;
assign micromatrizz[11][132] = 9'b111111111;
assign micromatrizz[11][133] = 9'b111111111;
assign micromatrizz[11][134] = 9'b111111111;
assign micromatrizz[11][135] = 9'b111111111;
assign micromatrizz[11][136] = 9'b111111111;
assign micromatrizz[11][137] = 9'b111111111;
assign micromatrizz[11][138] = 9'b111111111;
assign micromatrizz[11][139] = 9'b111111111;
assign micromatrizz[11][140] = 9'b111111111;
assign micromatrizz[11][141] = 9'b111111111;
assign micromatrizz[11][142] = 9'b111111111;
assign micromatrizz[11][143] = 9'b111111111;
assign micromatrizz[11][144] = 9'b111111111;
assign micromatrizz[11][145] = 9'b111111111;
assign micromatrizz[11][146] = 9'b111111111;
assign micromatrizz[11][147] = 9'b111111111;
assign micromatrizz[11][148] = 9'b111111111;
assign micromatrizz[11][149] = 9'b111111111;
assign micromatrizz[11][150] = 9'b111111111;
assign micromatrizz[11][151] = 9'b111111111;
assign micromatrizz[11][152] = 9'b111111111;
assign micromatrizz[11][153] = 9'b111111111;
assign micromatrizz[11][154] = 9'b111111111;
assign micromatrizz[11][155] = 9'b111111111;
assign micromatrizz[11][156] = 9'b111111111;
assign micromatrizz[11][157] = 9'b111111111;
assign micromatrizz[11][158] = 9'b111111111;
assign micromatrizz[11][159] = 9'b111111111;
assign micromatrizz[11][160] = 9'b111111111;
assign micromatrizz[11][161] = 9'b111111111;
assign micromatrizz[11][162] = 9'b111111111;
assign micromatrizz[11][163] = 9'b111111111;
assign micromatrizz[11][164] = 9'b111111111;
assign micromatrizz[11][165] = 9'b111111111;
assign micromatrizz[11][166] = 9'b111111111;
assign micromatrizz[11][167] = 9'b111111111;
assign micromatrizz[11][168] = 9'b111111111;
assign micromatrizz[11][169] = 9'b111111111;
assign micromatrizz[11][170] = 9'b111111111;
assign micromatrizz[11][171] = 9'b111111111;
assign micromatrizz[11][172] = 9'b111111111;
assign micromatrizz[11][173] = 9'b111111111;
assign micromatrizz[11][174] = 9'b111111111;
assign micromatrizz[11][175] = 9'b111111111;
assign micromatrizz[11][176] = 9'b111111111;
assign micromatrizz[11][177] = 9'b111111111;
assign micromatrizz[11][178] = 9'b111111111;
assign micromatrizz[11][179] = 9'b111111111;
assign micromatrizz[11][180] = 9'b111111111;
assign micromatrizz[11][181] = 9'b111111111;
assign micromatrizz[11][182] = 9'b111111111;
assign micromatrizz[11][183] = 9'b111111111;
assign micromatrizz[11][184] = 9'b111111111;
assign micromatrizz[11][185] = 9'b111111111;
assign micromatrizz[11][186] = 9'b111111111;
assign micromatrizz[11][187] = 9'b111111111;
assign micromatrizz[11][188] = 9'b111111111;
assign micromatrizz[11][189] = 9'b111111111;
assign micromatrizz[11][190] = 9'b111111111;
assign micromatrizz[11][191] = 9'b111111111;
assign micromatrizz[11][192] = 9'b111111111;
assign micromatrizz[11][193] = 9'b111111111;
assign micromatrizz[11][194] = 9'b111111111;
assign micromatrizz[11][195] = 9'b111111111;
assign micromatrizz[11][196] = 9'b111111111;
assign micromatrizz[11][197] = 9'b111111111;
assign micromatrizz[11][198] = 9'b111111111;
assign micromatrizz[11][199] = 9'b111111111;
assign micromatrizz[11][200] = 9'b111111111;
assign micromatrizz[11][201] = 9'b111111111;
assign micromatrizz[11][202] = 9'b111111111;
assign micromatrizz[11][203] = 9'b111111111;
assign micromatrizz[11][204] = 9'b111111111;
assign micromatrizz[11][205] = 9'b111111111;
assign micromatrizz[11][206] = 9'b111111111;
assign micromatrizz[11][207] = 9'b111111111;
assign micromatrizz[11][208] = 9'b111111111;
assign micromatrizz[11][209] = 9'b111111111;
assign micromatrizz[11][210] = 9'b111111111;
assign micromatrizz[11][211] = 9'b111111111;
assign micromatrizz[11][212] = 9'b111111111;
assign micromatrizz[11][213] = 9'b111111111;
assign micromatrizz[11][214] = 9'b111111111;
assign micromatrizz[11][215] = 9'b111111111;
assign micromatrizz[11][216] = 9'b111111111;
assign micromatrizz[11][217] = 9'b111111111;
assign micromatrizz[11][218] = 9'b111111111;
assign micromatrizz[11][219] = 9'b111111111;
assign micromatrizz[11][220] = 9'b111111111;
assign micromatrizz[11][221] = 9'b111111111;
assign micromatrizz[11][222] = 9'b111111111;
assign micromatrizz[11][223] = 9'b111111111;
assign micromatrizz[11][224] = 9'b111111111;
assign micromatrizz[11][225] = 9'b111111111;
assign micromatrizz[11][226] = 9'b111111111;
assign micromatrizz[11][227] = 9'b111111111;
assign micromatrizz[11][228] = 9'b111111111;
assign micromatrizz[11][229] = 9'b111111111;
assign micromatrizz[11][230] = 9'b111111111;
assign micromatrizz[11][231] = 9'b111111111;
assign micromatrizz[11][232] = 9'b111111111;
assign micromatrizz[11][233] = 9'b111111111;
assign micromatrizz[11][234] = 9'b111111111;
assign micromatrizz[11][235] = 9'b111111111;
assign micromatrizz[11][236] = 9'b111111111;
assign micromatrizz[11][237] = 9'b111111111;
assign micromatrizz[11][238] = 9'b111111111;
assign micromatrizz[11][239] = 9'b111111111;
assign micromatrizz[11][240] = 9'b111111111;
assign micromatrizz[11][241] = 9'b111111111;
assign micromatrizz[11][242] = 9'b111111111;
assign micromatrizz[11][243] = 9'b111111111;
assign micromatrizz[11][244] = 9'b111111111;
assign micromatrizz[11][245] = 9'b111111111;
assign micromatrizz[11][246] = 9'b111111111;
assign micromatrizz[11][247] = 9'b111111111;
assign micromatrizz[11][248] = 9'b111111111;
assign micromatrizz[11][249] = 9'b111111111;
assign micromatrizz[11][250] = 9'b111111111;
assign micromatrizz[11][251] = 9'b111111111;
assign micromatrizz[11][252] = 9'b111111111;
assign micromatrizz[11][253] = 9'b111111111;
assign micromatrizz[11][254] = 9'b111111111;
assign micromatrizz[11][255] = 9'b111111111;
assign micromatrizz[11][256] = 9'b111111111;
assign micromatrizz[11][257] = 9'b111111111;
assign micromatrizz[11][258] = 9'b111111111;
assign micromatrizz[11][259] = 9'b111111111;
assign micromatrizz[11][260] = 9'b111111111;
assign micromatrizz[11][261] = 9'b111111111;
assign micromatrizz[11][262] = 9'b111111111;
assign micromatrizz[11][263] = 9'b111111111;
assign micromatrizz[11][264] = 9'b111111111;
assign micromatrizz[11][265] = 9'b111111111;
assign micromatrizz[11][266] = 9'b111111111;
assign micromatrizz[11][267] = 9'b111111111;
assign micromatrizz[11][268] = 9'b111111111;
assign micromatrizz[11][269] = 9'b111111111;
assign micromatrizz[11][270] = 9'b111111111;
assign micromatrizz[11][271] = 9'b111111111;
assign micromatrizz[11][272] = 9'b111111111;
assign micromatrizz[11][273] = 9'b111111111;
assign micromatrizz[11][274] = 9'b111111111;
assign micromatrizz[11][275] = 9'b111111111;
assign micromatrizz[11][276] = 9'b111111111;
assign micromatrizz[11][277] = 9'b111111111;
assign micromatrizz[11][278] = 9'b111111111;
assign micromatrizz[11][279] = 9'b111111111;
assign micromatrizz[11][280] = 9'b111111111;
assign micromatrizz[11][281] = 9'b111111111;
assign micromatrizz[11][282] = 9'b111111111;
assign micromatrizz[11][283] = 9'b111111111;
assign micromatrizz[11][284] = 9'b111111111;
assign micromatrizz[11][285] = 9'b111111111;
assign micromatrizz[11][286] = 9'b111111111;
assign micromatrizz[11][287] = 9'b111111111;
assign micromatrizz[11][288] = 9'b111111111;
assign micromatrizz[11][289] = 9'b111111111;
assign micromatrizz[11][290] = 9'b111111111;
assign micromatrizz[11][291] = 9'b111111111;
assign micromatrizz[11][292] = 9'b111111111;
assign micromatrizz[11][293] = 9'b111111111;
assign micromatrizz[11][294] = 9'b111111111;
assign micromatrizz[11][295] = 9'b111111111;
assign micromatrizz[11][296] = 9'b111111111;
assign micromatrizz[11][297] = 9'b111111111;
assign micromatrizz[11][298] = 9'b111111111;
assign micromatrizz[11][299] = 9'b111111111;
assign micromatrizz[11][300] = 9'b111111111;
assign micromatrizz[11][301] = 9'b111111111;
assign micromatrizz[11][302] = 9'b111111111;
assign micromatrizz[11][303] = 9'b111111111;
assign micromatrizz[11][304] = 9'b111111111;
assign micromatrizz[11][305] = 9'b111111111;
assign micromatrizz[11][306] = 9'b111111111;
assign micromatrizz[11][307] = 9'b111111111;
assign micromatrizz[11][308] = 9'b111111111;
assign micromatrizz[11][309] = 9'b111111111;
assign micromatrizz[11][310] = 9'b111111111;
assign micromatrizz[11][311] = 9'b111111111;
assign micromatrizz[11][312] = 9'b111111111;
assign micromatrizz[11][313] = 9'b111111111;
assign micromatrizz[11][314] = 9'b111111111;
assign micromatrizz[11][315] = 9'b111111111;
assign micromatrizz[11][316] = 9'b111111111;
assign micromatrizz[11][317] = 9'b111111111;
assign micromatrizz[11][318] = 9'b111111111;
assign micromatrizz[11][319] = 9'b111111111;
assign micromatrizz[11][320] = 9'b111111111;
assign micromatrizz[11][321] = 9'b111111111;
assign micromatrizz[11][322] = 9'b111111111;
assign micromatrizz[11][323] = 9'b111111111;
assign micromatrizz[11][324] = 9'b111111111;
assign micromatrizz[11][325] = 9'b111111111;
assign micromatrizz[11][326] = 9'b111111111;
assign micromatrizz[11][327] = 9'b111111111;
assign micromatrizz[11][328] = 9'b111111111;
assign micromatrizz[11][329] = 9'b111111111;
assign micromatrizz[11][330] = 9'b111111111;
assign micromatrizz[11][331] = 9'b111111111;
assign micromatrizz[11][332] = 9'b111111111;
assign micromatrizz[11][333] = 9'b111111111;
assign micromatrizz[11][334] = 9'b111111111;
assign micromatrizz[11][335] = 9'b111111111;
assign micromatrizz[11][336] = 9'b111111111;
assign micromatrizz[11][337] = 9'b111111111;
assign micromatrizz[11][338] = 9'b111111111;
assign micromatrizz[11][339] = 9'b111111111;
assign micromatrizz[11][340] = 9'b111111111;
assign micromatrizz[11][341] = 9'b111111111;
assign micromatrizz[11][342] = 9'b111111111;
assign micromatrizz[11][343] = 9'b111111111;
assign micromatrizz[11][344] = 9'b111111111;
assign micromatrizz[11][345] = 9'b111111111;
assign micromatrizz[11][346] = 9'b111111111;
assign micromatrizz[11][347] = 9'b111111111;
assign micromatrizz[11][348] = 9'b111111111;
assign micromatrizz[11][349] = 9'b111111111;
assign micromatrizz[11][350] = 9'b111111111;
assign micromatrizz[11][351] = 9'b111111111;
assign micromatrizz[11][352] = 9'b111111111;
assign micromatrizz[11][353] = 9'b111111111;
assign micromatrizz[11][354] = 9'b111111111;
assign micromatrizz[11][355] = 9'b111111111;
assign micromatrizz[11][356] = 9'b111111111;
assign micromatrizz[11][357] = 9'b111111111;
assign micromatrizz[11][358] = 9'b111111111;
assign micromatrizz[11][359] = 9'b111111111;
assign micromatrizz[11][360] = 9'b111111111;
assign micromatrizz[11][361] = 9'b111111111;
assign micromatrizz[11][362] = 9'b111111111;
assign micromatrizz[11][363] = 9'b111111111;
assign micromatrizz[11][364] = 9'b111111111;
assign micromatrizz[11][365] = 9'b111111111;
assign micromatrizz[11][366] = 9'b111111111;
assign micromatrizz[11][367] = 9'b111111111;
assign micromatrizz[11][368] = 9'b111111111;
assign micromatrizz[11][369] = 9'b111111111;
assign micromatrizz[11][370] = 9'b111111111;
assign micromatrizz[11][371] = 9'b111111111;
assign micromatrizz[11][372] = 9'b111111111;
assign micromatrizz[11][373] = 9'b111111111;
assign micromatrizz[11][374] = 9'b111111111;
assign micromatrizz[11][375] = 9'b111111111;
assign micromatrizz[11][376] = 9'b111111111;
assign micromatrizz[11][377] = 9'b111111111;
assign micromatrizz[11][378] = 9'b111111111;
assign micromatrizz[11][379] = 9'b111111111;
assign micromatrizz[11][380] = 9'b111111111;
assign micromatrizz[11][381] = 9'b111111111;
assign micromatrizz[11][382] = 9'b111111111;
assign micromatrizz[11][383] = 9'b111111111;
assign micromatrizz[11][384] = 9'b111111111;
assign micromatrizz[11][385] = 9'b111111111;
assign micromatrizz[11][386] = 9'b111111111;
assign micromatrizz[11][387] = 9'b111111111;
assign micromatrizz[11][388] = 9'b111111111;
assign micromatrizz[11][389] = 9'b111111111;
assign micromatrizz[11][390] = 9'b111111111;
assign micromatrizz[11][391] = 9'b111111111;
assign micromatrizz[11][392] = 9'b111111111;
assign micromatrizz[11][393] = 9'b111111111;
assign micromatrizz[11][394] = 9'b111111111;
assign micromatrizz[11][395] = 9'b111111111;
assign micromatrizz[11][396] = 9'b111111111;
assign micromatrizz[11][397] = 9'b111111111;
assign micromatrizz[11][398] = 9'b111111111;
assign micromatrizz[11][399] = 9'b111111111;
assign micromatrizz[11][400] = 9'b111111111;
assign micromatrizz[11][401] = 9'b111111111;
assign micromatrizz[11][402] = 9'b111111111;
assign micromatrizz[11][403] = 9'b111111111;
assign micromatrizz[11][404] = 9'b111111111;
assign micromatrizz[11][405] = 9'b111111111;
assign micromatrizz[11][406] = 9'b111111111;
assign micromatrizz[11][407] = 9'b111111111;
assign micromatrizz[11][408] = 9'b111111111;
assign micromatrizz[11][409] = 9'b111111111;
assign micromatrizz[11][410] = 9'b111111111;
assign micromatrizz[11][411] = 9'b111111111;
assign micromatrizz[11][412] = 9'b111111111;
assign micromatrizz[11][413] = 9'b111111111;
assign micromatrizz[11][414] = 9'b111111111;
assign micromatrizz[11][415] = 9'b111111111;
assign micromatrizz[11][416] = 9'b111111111;
assign micromatrizz[11][417] = 9'b111111111;
assign micromatrizz[11][418] = 9'b111111111;
assign micromatrizz[11][419] = 9'b111111111;
assign micromatrizz[11][420] = 9'b111111111;
assign micromatrizz[11][421] = 9'b111111111;
assign micromatrizz[11][422] = 9'b111111111;
assign micromatrizz[11][423] = 9'b111111111;
assign micromatrizz[11][424] = 9'b111111111;
assign micromatrizz[11][425] = 9'b111111111;
assign micromatrizz[11][426] = 9'b111111111;
assign micromatrizz[11][427] = 9'b111111111;
assign micromatrizz[11][428] = 9'b111111111;
assign micromatrizz[11][429] = 9'b111111111;
assign micromatrizz[11][430] = 9'b111111111;
assign micromatrizz[11][431] = 9'b111111111;
assign micromatrizz[11][432] = 9'b111111111;
assign micromatrizz[11][433] = 9'b111111111;
assign micromatrizz[11][434] = 9'b111111111;
assign micromatrizz[11][435] = 9'b111111111;
assign micromatrizz[11][436] = 9'b111111111;
assign micromatrizz[11][437] = 9'b111111111;
assign micromatrizz[11][438] = 9'b111111111;
assign micromatrizz[11][439] = 9'b111111111;
assign micromatrizz[11][440] = 9'b111111111;
assign micromatrizz[11][441] = 9'b111111111;
assign micromatrizz[11][442] = 9'b111111111;
assign micromatrizz[11][443] = 9'b111111111;
assign micromatrizz[11][444] = 9'b111111111;
assign micromatrizz[11][445] = 9'b111111111;
assign micromatrizz[11][446] = 9'b111111111;
assign micromatrizz[11][447] = 9'b111111111;
assign micromatrizz[11][448] = 9'b111111111;
assign micromatrizz[11][449] = 9'b111111111;
assign micromatrizz[11][450] = 9'b111111111;
assign micromatrizz[11][451] = 9'b111111111;
assign micromatrizz[11][452] = 9'b111111111;
assign micromatrizz[11][453] = 9'b111111111;
assign micromatrizz[11][454] = 9'b111111111;
assign micromatrizz[11][455] = 9'b111111111;
assign micromatrizz[11][456] = 9'b111111111;
assign micromatrizz[11][457] = 9'b111111111;
assign micromatrizz[11][458] = 9'b111111111;
assign micromatrizz[11][459] = 9'b111111111;
assign micromatrizz[11][460] = 9'b111111111;
assign micromatrizz[11][461] = 9'b111111111;
assign micromatrizz[11][462] = 9'b111111111;
assign micromatrizz[11][463] = 9'b111111111;
assign micromatrizz[11][464] = 9'b111111111;
assign micromatrizz[11][465] = 9'b111111111;
assign micromatrizz[11][466] = 9'b111111111;
assign micromatrizz[11][467] = 9'b111111111;
assign micromatrizz[11][468] = 9'b111111111;
assign micromatrizz[11][469] = 9'b111111111;
assign micromatrizz[11][470] = 9'b111111111;
assign micromatrizz[11][471] = 9'b111111111;
assign micromatrizz[11][472] = 9'b111111111;
assign micromatrizz[11][473] = 9'b111111111;
assign micromatrizz[11][474] = 9'b111111111;
assign micromatrizz[11][475] = 9'b111111111;
assign micromatrizz[11][476] = 9'b111111111;
assign micromatrizz[11][477] = 9'b111111111;
assign micromatrizz[11][478] = 9'b111111111;
assign micromatrizz[11][479] = 9'b111111111;
assign micromatrizz[11][480] = 9'b111111111;
assign micromatrizz[11][481] = 9'b111111111;
assign micromatrizz[11][482] = 9'b111111111;
assign micromatrizz[11][483] = 9'b111111111;
assign micromatrizz[11][484] = 9'b111111111;
assign micromatrizz[11][485] = 9'b111111111;
assign micromatrizz[11][486] = 9'b111111111;
assign micromatrizz[11][487] = 9'b111111111;
assign micromatrizz[11][488] = 9'b111111111;
assign micromatrizz[11][489] = 9'b111111111;
assign micromatrizz[11][490] = 9'b111111111;
assign micromatrizz[11][491] = 9'b111111111;
assign micromatrizz[11][492] = 9'b111111111;
assign micromatrizz[11][493] = 9'b111111111;
assign micromatrizz[11][494] = 9'b111111111;
assign micromatrizz[11][495] = 9'b111111111;
assign micromatrizz[11][496] = 9'b111111111;
assign micromatrizz[11][497] = 9'b111111111;
assign micromatrizz[11][498] = 9'b111111111;
assign micromatrizz[11][499] = 9'b111111111;
assign micromatrizz[11][500] = 9'b111111111;
assign micromatrizz[11][501] = 9'b111111111;
assign micromatrizz[11][502] = 9'b111111111;
assign micromatrizz[11][503] = 9'b111111111;
assign micromatrizz[11][504] = 9'b111111111;
assign micromatrizz[11][505] = 9'b111111111;
assign micromatrizz[11][506] = 9'b111111111;
assign micromatrizz[11][507] = 9'b111111111;
assign micromatrizz[11][508] = 9'b111111111;
assign micromatrizz[11][509] = 9'b111111111;
assign micromatrizz[11][510] = 9'b111111111;
assign micromatrizz[11][511] = 9'b111111111;
assign micromatrizz[11][512] = 9'b111111111;
assign micromatrizz[11][513] = 9'b111111111;
assign micromatrizz[11][514] = 9'b111111111;
assign micromatrizz[11][515] = 9'b111111111;
assign micromatrizz[11][516] = 9'b111111111;
assign micromatrizz[11][517] = 9'b111111111;
assign micromatrizz[11][518] = 9'b111111111;
assign micromatrizz[11][519] = 9'b111111111;
assign micromatrizz[11][520] = 9'b111111111;
assign micromatrizz[11][521] = 9'b111111111;
assign micromatrizz[11][522] = 9'b111111111;
assign micromatrizz[11][523] = 9'b111111111;
assign micromatrizz[11][524] = 9'b111111111;
assign micromatrizz[11][525] = 9'b111111111;
assign micromatrizz[11][526] = 9'b111111111;
assign micromatrizz[11][527] = 9'b111111111;
assign micromatrizz[11][528] = 9'b111111111;
assign micromatrizz[11][529] = 9'b111111111;
assign micromatrizz[11][530] = 9'b111111111;
assign micromatrizz[11][531] = 9'b111111111;
assign micromatrizz[11][532] = 9'b111111111;
assign micromatrizz[11][533] = 9'b111111111;
assign micromatrizz[11][534] = 9'b111111111;
assign micromatrizz[11][535] = 9'b111111111;
assign micromatrizz[11][536] = 9'b111111111;
assign micromatrizz[11][537] = 9'b111111111;
assign micromatrizz[11][538] = 9'b111111111;
assign micromatrizz[11][539] = 9'b111111111;
assign micromatrizz[11][540] = 9'b111111111;
assign micromatrizz[11][541] = 9'b111111111;
assign micromatrizz[11][542] = 9'b111111111;
assign micromatrizz[11][543] = 9'b111111111;
assign micromatrizz[11][544] = 9'b111111111;
assign micromatrizz[11][545] = 9'b111111111;
assign micromatrizz[11][546] = 9'b111111111;
assign micromatrizz[11][547] = 9'b111111111;
assign micromatrizz[11][548] = 9'b111111111;
assign micromatrizz[11][549] = 9'b111111111;
assign micromatrizz[11][550] = 9'b111111111;
assign micromatrizz[11][551] = 9'b111111111;
assign micromatrizz[11][552] = 9'b111111111;
assign micromatrizz[11][553] = 9'b111111111;
assign micromatrizz[11][554] = 9'b111111111;
assign micromatrizz[11][555] = 9'b111111111;
assign micromatrizz[11][556] = 9'b111111111;
assign micromatrizz[11][557] = 9'b111111111;
assign micromatrizz[11][558] = 9'b111111111;
assign micromatrizz[11][559] = 9'b111111111;
assign micromatrizz[11][560] = 9'b111111111;
assign micromatrizz[11][561] = 9'b111111111;
assign micromatrizz[11][562] = 9'b111111111;
assign micromatrizz[11][563] = 9'b111111111;
assign micromatrizz[11][564] = 9'b111111111;
assign micromatrizz[11][565] = 9'b111111111;
assign micromatrizz[11][566] = 9'b111111111;
assign micromatrizz[11][567] = 9'b111111111;
assign micromatrizz[11][568] = 9'b111111111;
assign micromatrizz[11][569] = 9'b111111111;
assign micromatrizz[11][570] = 9'b111111111;
assign micromatrizz[11][571] = 9'b111111111;
assign micromatrizz[11][572] = 9'b111111111;
assign micromatrizz[11][573] = 9'b111111111;
assign micromatrizz[11][574] = 9'b111111111;
assign micromatrizz[11][575] = 9'b111111111;
assign micromatrizz[11][576] = 9'b111111111;
assign micromatrizz[11][577] = 9'b111111111;
assign micromatrizz[11][578] = 9'b111111111;
assign micromatrizz[11][579] = 9'b111111111;
assign micromatrizz[11][580] = 9'b111111111;
assign micromatrizz[11][581] = 9'b111111111;
assign micromatrizz[11][582] = 9'b111111111;
assign micromatrizz[11][583] = 9'b111111111;
assign micromatrizz[11][584] = 9'b111111111;
assign micromatrizz[11][585] = 9'b111111111;
assign micromatrizz[11][586] = 9'b111111111;
assign micromatrizz[11][587] = 9'b111111111;
assign micromatrizz[11][588] = 9'b111111111;
assign micromatrizz[11][589] = 9'b111111111;
assign micromatrizz[11][590] = 9'b111111111;
assign micromatrizz[11][591] = 9'b111111111;
assign micromatrizz[11][592] = 9'b111111111;
assign micromatrizz[11][593] = 9'b111111111;
assign micromatrizz[11][594] = 9'b111111111;
assign micromatrizz[11][595] = 9'b111111111;
assign micromatrizz[11][596] = 9'b111111111;
assign micromatrizz[11][597] = 9'b111111111;
assign micromatrizz[11][598] = 9'b111111111;
assign micromatrizz[11][599] = 9'b111111111;
assign micromatrizz[11][600] = 9'b111111111;
assign micromatrizz[11][601] = 9'b111111111;
assign micromatrizz[11][602] = 9'b111111111;
assign micromatrizz[11][603] = 9'b111111111;
assign micromatrizz[11][604] = 9'b111111111;
assign micromatrizz[11][605] = 9'b111111111;
assign micromatrizz[11][606] = 9'b111111111;
assign micromatrizz[11][607] = 9'b111111111;
assign micromatrizz[11][608] = 9'b111111111;
assign micromatrizz[11][609] = 9'b111111111;
assign micromatrizz[11][610] = 9'b111111111;
assign micromatrizz[11][611] = 9'b111111111;
assign micromatrizz[11][612] = 9'b111111111;
assign micromatrizz[11][613] = 9'b111111111;
assign micromatrizz[11][614] = 9'b111111111;
assign micromatrizz[11][615] = 9'b111111111;
assign micromatrizz[11][616] = 9'b111111111;
assign micromatrizz[11][617] = 9'b111111111;
assign micromatrizz[11][618] = 9'b111111111;
assign micromatrizz[11][619] = 9'b111111111;
assign micromatrizz[11][620] = 9'b111111111;
assign micromatrizz[11][621] = 9'b111111111;
assign micromatrizz[11][622] = 9'b111111111;
assign micromatrizz[11][623] = 9'b111111111;
assign micromatrizz[11][624] = 9'b111111111;
assign micromatrizz[11][625] = 9'b111111111;
assign micromatrizz[11][626] = 9'b111111111;
assign micromatrizz[11][627] = 9'b111111111;
assign micromatrizz[11][628] = 9'b111111111;
assign micromatrizz[11][629] = 9'b111111111;
assign micromatrizz[11][630] = 9'b111111111;
assign micromatrizz[11][631] = 9'b111111111;
assign micromatrizz[11][632] = 9'b111111111;
assign micromatrizz[11][633] = 9'b111111111;
assign micromatrizz[11][634] = 9'b111111111;
assign micromatrizz[11][635] = 9'b111111111;
assign micromatrizz[11][636] = 9'b111111111;
assign micromatrizz[11][637] = 9'b111111111;
assign micromatrizz[11][638] = 9'b111111111;
assign micromatrizz[11][639] = 9'b111111111;
assign micromatrizz[12][0] = 9'b111111111;
assign micromatrizz[12][1] = 9'b111111111;
assign micromatrizz[12][2] = 9'b111111111;
assign micromatrizz[12][3] = 9'b111111111;
assign micromatrizz[12][4] = 9'b111111111;
assign micromatrizz[12][5] = 9'b111111111;
assign micromatrizz[12][6] = 9'b111111111;
assign micromatrizz[12][7] = 9'b111111111;
assign micromatrizz[12][8] = 9'b111111111;
assign micromatrizz[12][9] = 9'b111111111;
assign micromatrizz[12][10] = 9'b111111111;
assign micromatrizz[12][11] = 9'b111111111;
assign micromatrizz[12][12] = 9'b111111111;
assign micromatrizz[12][13] = 9'b111111111;
assign micromatrizz[12][14] = 9'b111111111;
assign micromatrizz[12][15] = 9'b111111111;
assign micromatrizz[12][16] = 9'b111111111;
assign micromatrizz[12][17] = 9'b111111111;
assign micromatrizz[12][18] = 9'b111111111;
assign micromatrizz[12][19] = 9'b111111111;
assign micromatrizz[12][20] = 9'b111111111;
assign micromatrizz[12][21] = 9'b111111111;
assign micromatrizz[12][22] = 9'b111111111;
assign micromatrizz[12][23] = 9'b111111111;
assign micromatrizz[12][24] = 9'b111111111;
assign micromatrizz[12][25] = 9'b111111111;
assign micromatrizz[12][26] = 9'b111111111;
assign micromatrizz[12][27] = 9'b111111111;
assign micromatrizz[12][28] = 9'b111111111;
assign micromatrizz[12][29] = 9'b111111111;
assign micromatrizz[12][30] = 9'b111111111;
assign micromatrizz[12][31] = 9'b111111111;
assign micromatrizz[12][32] = 9'b111111111;
assign micromatrizz[12][33] = 9'b111111111;
assign micromatrizz[12][34] = 9'b111111111;
assign micromatrizz[12][35] = 9'b111111111;
assign micromatrizz[12][36] = 9'b111111111;
assign micromatrizz[12][37] = 9'b111111111;
assign micromatrizz[12][38] = 9'b111111111;
assign micromatrizz[12][39] = 9'b111111111;
assign micromatrizz[12][40] = 9'b111111111;
assign micromatrizz[12][41] = 9'b111111111;
assign micromatrizz[12][42] = 9'b111111111;
assign micromatrizz[12][43] = 9'b111111111;
assign micromatrizz[12][44] = 9'b111111111;
assign micromatrizz[12][45] = 9'b111111111;
assign micromatrizz[12][46] = 9'b111111111;
assign micromatrizz[12][47] = 9'b111111111;
assign micromatrizz[12][48] = 9'b111111111;
assign micromatrizz[12][49] = 9'b111111111;
assign micromatrizz[12][50] = 9'b111111111;
assign micromatrizz[12][51] = 9'b111111111;
assign micromatrizz[12][52] = 9'b111111111;
assign micromatrizz[12][53] = 9'b111111111;
assign micromatrizz[12][54] = 9'b111111111;
assign micromatrizz[12][55] = 9'b111111111;
assign micromatrizz[12][56] = 9'b111111111;
assign micromatrizz[12][57] = 9'b111111111;
assign micromatrizz[12][58] = 9'b111111111;
assign micromatrizz[12][59] = 9'b111111111;
assign micromatrizz[12][60] = 9'b111111111;
assign micromatrizz[12][61] = 9'b111111111;
assign micromatrizz[12][62] = 9'b111111111;
assign micromatrizz[12][63] = 9'b111111111;
assign micromatrizz[12][64] = 9'b111111111;
assign micromatrizz[12][65] = 9'b111111111;
assign micromatrizz[12][66] = 9'b111111111;
assign micromatrizz[12][67] = 9'b111111111;
assign micromatrizz[12][68] = 9'b111111111;
assign micromatrizz[12][69] = 9'b111111111;
assign micromatrizz[12][70] = 9'b111111111;
assign micromatrizz[12][71] = 9'b111111111;
assign micromatrizz[12][72] = 9'b111111111;
assign micromatrizz[12][73] = 9'b111111111;
assign micromatrizz[12][74] = 9'b111111111;
assign micromatrizz[12][75] = 9'b111111111;
assign micromatrizz[12][76] = 9'b111111111;
assign micromatrizz[12][77] = 9'b111111111;
assign micromatrizz[12][78] = 9'b111111111;
assign micromatrizz[12][79] = 9'b111111111;
assign micromatrizz[12][80] = 9'b111111111;
assign micromatrizz[12][81] = 9'b111111111;
assign micromatrizz[12][82] = 9'b111111111;
assign micromatrizz[12][83] = 9'b111111111;
assign micromatrizz[12][84] = 9'b111111111;
assign micromatrizz[12][85] = 9'b111111111;
assign micromatrizz[12][86] = 9'b111111111;
assign micromatrizz[12][87] = 9'b111111111;
assign micromatrizz[12][88] = 9'b111111111;
assign micromatrizz[12][89] = 9'b111111111;
assign micromatrizz[12][90] = 9'b111111111;
assign micromatrizz[12][91] = 9'b111111111;
assign micromatrizz[12][92] = 9'b111111111;
assign micromatrizz[12][93] = 9'b111111111;
assign micromatrizz[12][94] = 9'b111111111;
assign micromatrizz[12][95] = 9'b111111111;
assign micromatrizz[12][96] = 9'b111111111;
assign micromatrizz[12][97] = 9'b111111111;
assign micromatrizz[12][98] = 9'b111111111;
assign micromatrizz[12][99] = 9'b111111111;
assign micromatrizz[12][100] = 9'b111111111;
assign micromatrizz[12][101] = 9'b111111111;
assign micromatrizz[12][102] = 9'b111111111;
assign micromatrizz[12][103] = 9'b111111111;
assign micromatrizz[12][104] = 9'b111111111;
assign micromatrizz[12][105] = 9'b111111111;
assign micromatrizz[12][106] = 9'b111111111;
assign micromatrizz[12][107] = 9'b111111111;
assign micromatrizz[12][108] = 9'b111111111;
assign micromatrizz[12][109] = 9'b111111111;
assign micromatrizz[12][110] = 9'b111111111;
assign micromatrizz[12][111] = 9'b111111111;
assign micromatrizz[12][112] = 9'b111111111;
assign micromatrizz[12][113] = 9'b111111111;
assign micromatrizz[12][114] = 9'b111111111;
assign micromatrizz[12][115] = 9'b111111111;
assign micromatrizz[12][116] = 9'b111111111;
assign micromatrizz[12][117] = 9'b111111111;
assign micromatrizz[12][118] = 9'b111111111;
assign micromatrizz[12][119] = 9'b111111111;
assign micromatrizz[12][120] = 9'b111111111;
assign micromatrizz[12][121] = 9'b111111111;
assign micromatrizz[12][122] = 9'b111111111;
assign micromatrizz[12][123] = 9'b111111111;
assign micromatrizz[12][124] = 9'b111111111;
assign micromatrizz[12][125] = 9'b111111111;
assign micromatrizz[12][126] = 9'b111111111;
assign micromatrizz[12][127] = 9'b111111111;
assign micromatrizz[12][128] = 9'b111111111;
assign micromatrizz[12][129] = 9'b111111111;
assign micromatrizz[12][130] = 9'b111111111;
assign micromatrizz[12][131] = 9'b111111111;
assign micromatrizz[12][132] = 9'b111111111;
assign micromatrizz[12][133] = 9'b111111111;
assign micromatrizz[12][134] = 9'b111111111;
assign micromatrizz[12][135] = 9'b111111111;
assign micromatrizz[12][136] = 9'b111111111;
assign micromatrizz[12][137] = 9'b111111111;
assign micromatrizz[12][138] = 9'b111111111;
assign micromatrizz[12][139] = 9'b111111111;
assign micromatrizz[12][140] = 9'b111111111;
assign micromatrizz[12][141] = 9'b111111111;
assign micromatrizz[12][142] = 9'b111111111;
assign micromatrizz[12][143] = 9'b111111111;
assign micromatrizz[12][144] = 9'b111111111;
assign micromatrizz[12][145] = 9'b111111111;
assign micromatrizz[12][146] = 9'b111111111;
assign micromatrizz[12][147] = 9'b111111111;
assign micromatrizz[12][148] = 9'b111111111;
assign micromatrizz[12][149] = 9'b111111111;
assign micromatrizz[12][150] = 9'b111111111;
assign micromatrizz[12][151] = 9'b111111111;
assign micromatrizz[12][152] = 9'b111111111;
assign micromatrizz[12][153] = 9'b111111111;
assign micromatrizz[12][154] = 9'b111111111;
assign micromatrizz[12][155] = 9'b111111111;
assign micromatrizz[12][156] = 9'b111111111;
assign micromatrizz[12][157] = 9'b111111111;
assign micromatrizz[12][158] = 9'b111111111;
assign micromatrizz[12][159] = 9'b111111111;
assign micromatrizz[12][160] = 9'b111111111;
assign micromatrizz[12][161] = 9'b111111111;
assign micromatrizz[12][162] = 9'b111111111;
assign micromatrizz[12][163] = 9'b111111111;
assign micromatrizz[12][164] = 9'b111111111;
assign micromatrizz[12][165] = 9'b111111111;
assign micromatrizz[12][166] = 9'b111111111;
assign micromatrizz[12][167] = 9'b111111111;
assign micromatrizz[12][168] = 9'b111111111;
assign micromatrizz[12][169] = 9'b111111111;
assign micromatrizz[12][170] = 9'b111111111;
assign micromatrizz[12][171] = 9'b111111111;
assign micromatrizz[12][172] = 9'b111111111;
assign micromatrizz[12][173] = 9'b111111111;
assign micromatrizz[12][174] = 9'b111111111;
assign micromatrizz[12][175] = 9'b111111111;
assign micromatrizz[12][176] = 9'b111111111;
assign micromatrizz[12][177] = 9'b111111111;
assign micromatrizz[12][178] = 9'b111111111;
assign micromatrizz[12][179] = 9'b111111111;
assign micromatrizz[12][180] = 9'b111111111;
assign micromatrizz[12][181] = 9'b111111111;
assign micromatrizz[12][182] = 9'b111111111;
assign micromatrizz[12][183] = 9'b111111111;
assign micromatrizz[12][184] = 9'b111111111;
assign micromatrizz[12][185] = 9'b111111111;
assign micromatrizz[12][186] = 9'b111111111;
assign micromatrizz[12][187] = 9'b111111111;
assign micromatrizz[12][188] = 9'b111111111;
assign micromatrizz[12][189] = 9'b111111111;
assign micromatrizz[12][190] = 9'b111111111;
assign micromatrizz[12][191] = 9'b111111111;
assign micromatrizz[12][192] = 9'b111111111;
assign micromatrizz[12][193] = 9'b111111111;
assign micromatrizz[12][194] = 9'b111111111;
assign micromatrizz[12][195] = 9'b111111111;
assign micromatrizz[12][196] = 9'b111111111;
assign micromatrizz[12][197] = 9'b111111111;
assign micromatrizz[12][198] = 9'b111111111;
assign micromatrizz[12][199] = 9'b111111111;
assign micromatrizz[12][200] = 9'b111111111;
assign micromatrizz[12][201] = 9'b111111111;
assign micromatrizz[12][202] = 9'b111111111;
assign micromatrizz[12][203] = 9'b111111111;
assign micromatrizz[12][204] = 9'b111111111;
assign micromatrizz[12][205] = 9'b111111111;
assign micromatrizz[12][206] = 9'b111111111;
assign micromatrizz[12][207] = 9'b111111111;
assign micromatrizz[12][208] = 9'b111111111;
assign micromatrizz[12][209] = 9'b111111111;
assign micromatrizz[12][210] = 9'b111111111;
assign micromatrizz[12][211] = 9'b111111111;
assign micromatrizz[12][212] = 9'b111111111;
assign micromatrizz[12][213] = 9'b111111111;
assign micromatrizz[12][214] = 9'b111111111;
assign micromatrizz[12][215] = 9'b111111111;
assign micromatrizz[12][216] = 9'b111111111;
assign micromatrizz[12][217] = 9'b111111111;
assign micromatrizz[12][218] = 9'b111111111;
assign micromatrizz[12][219] = 9'b111111111;
assign micromatrizz[12][220] = 9'b111111111;
assign micromatrizz[12][221] = 9'b111111111;
assign micromatrizz[12][222] = 9'b111111111;
assign micromatrizz[12][223] = 9'b111111111;
assign micromatrizz[12][224] = 9'b111111111;
assign micromatrizz[12][225] = 9'b111111111;
assign micromatrizz[12][226] = 9'b111111111;
assign micromatrizz[12][227] = 9'b111111111;
assign micromatrizz[12][228] = 9'b111111111;
assign micromatrizz[12][229] = 9'b111111111;
assign micromatrizz[12][230] = 9'b111111111;
assign micromatrizz[12][231] = 9'b111111111;
assign micromatrizz[12][232] = 9'b111111111;
assign micromatrizz[12][233] = 9'b111111111;
assign micromatrizz[12][234] = 9'b111111111;
assign micromatrizz[12][235] = 9'b111111111;
assign micromatrizz[12][236] = 9'b111111111;
assign micromatrizz[12][237] = 9'b111111111;
assign micromatrizz[12][238] = 9'b111111111;
assign micromatrizz[12][239] = 9'b111111111;
assign micromatrizz[12][240] = 9'b111111111;
assign micromatrizz[12][241] = 9'b111111111;
assign micromatrizz[12][242] = 9'b111111111;
assign micromatrizz[12][243] = 9'b111111111;
assign micromatrizz[12][244] = 9'b111111111;
assign micromatrizz[12][245] = 9'b111111111;
assign micromatrizz[12][246] = 9'b111111111;
assign micromatrizz[12][247] = 9'b111111111;
assign micromatrizz[12][248] = 9'b111111111;
assign micromatrizz[12][249] = 9'b111111111;
assign micromatrizz[12][250] = 9'b111111111;
assign micromatrizz[12][251] = 9'b111111111;
assign micromatrizz[12][252] = 9'b111111111;
assign micromatrizz[12][253] = 9'b111111111;
assign micromatrizz[12][254] = 9'b111111111;
assign micromatrizz[12][255] = 9'b111111111;
assign micromatrizz[12][256] = 9'b111111111;
assign micromatrizz[12][257] = 9'b111111111;
assign micromatrizz[12][258] = 9'b111111111;
assign micromatrizz[12][259] = 9'b111111111;
assign micromatrizz[12][260] = 9'b111111111;
assign micromatrizz[12][261] = 9'b111111111;
assign micromatrizz[12][262] = 9'b111111111;
assign micromatrizz[12][263] = 9'b111111111;
assign micromatrizz[12][264] = 9'b111111111;
assign micromatrizz[12][265] = 9'b111111111;
assign micromatrizz[12][266] = 9'b111111111;
assign micromatrizz[12][267] = 9'b111111111;
assign micromatrizz[12][268] = 9'b111111111;
assign micromatrizz[12][269] = 9'b111111111;
assign micromatrizz[12][270] = 9'b111111111;
assign micromatrizz[12][271] = 9'b111111111;
assign micromatrizz[12][272] = 9'b111111111;
assign micromatrizz[12][273] = 9'b111111111;
assign micromatrizz[12][274] = 9'b111111111;
assign micromatrizz[12][275] = 9'b111111111;
assign micromatrizz[12][276] = 9'b111111111;
assign micromatrizz[12][277] = 9'b111111111;
assign micromatrizz[12][278] = 9'b111111111;
assign micromatrizz[12][279] = 9'b111111111;
assign micromatrizz[12][280] = 9'b111111111;
assign micromatrizz[12][281] = 9'b111111111;
assign micromatrizz[12][282] = 9'b111111111;
assign micromatrizz[12][283] = 9'b111111111;
assign micromatrizz[12][284] = 9'b111111111;
assign micromatrizz[12][285] = 9'b111111111;
assign micromatrizz[12][286] = 9'b111111111;
assign micromatrizz[12][287] = 9'b111111111;
assign micromatrizz[12][288] = 9'b111111111;
assign micromatrizz[12][289] = 9'b111111111;
assign micromatrizz[12][290] = 9'b111111111;
assign micromatrizz[12][291] = 9'b111111111;
assign micromatrizz[12][292] = 9'b111111111;
assign micromatrizz[12][293] = 9'b111111111;
assign micromatrizz[12][294] = 9'b111111111;
assign micromatrizz[12][295] = 9'b111111111;
assign micromatrizz[12][296] = 9'b111111111;
assign micromatrizz[12][297] = 9'b111111111;
assign micromatrizz[12][298] = 9'b111111111;
assign micromatrizz[12][299] = 9'b111111111;
assign micromatrizz[12][300] = 9'b111111111;
assign micromatrizz[12][301] = 9'b111111111;
assign micromatrizz[12][302] = 9'b111111111;
assign micromatrizz[12][303] = 9'b111111111;
assign micromatrizz[12][304] = 9'b111111111;
assign micromatrizz[12][305] = 9'b111111111;
assign micromatrizz[12][306] = 9'b111111111;
assign micromatrizz[12][307] = 9'b111111111;
assign micromatrizz[12][308] = 9'b111111111;
assign micromatrizz[12][309] = 9'b111111111;
assign micromatrizz[12][310] = 9'b111111111;
assign micromatrizz[12][311] = 9'b111111111;
assign micromatrizz[12][312] = 9'b111111111;
assign micromatrizz[12][313] = 9'b111111111;
assign micromatrizz[12][314] = 9'b111111111;
assign micromatrizz[12][315] = 9'b111111111;
assign micromatrizz[12][316] = 9'b111111111;
assign micromatrizz[12][317] = 9'b111111111;
assign micromatrizz[12][318] = 9'b111111111;
assign micromatrizz[12][319] = 9'b111111111;
assign micromatrizz[12][320] = 9'b111111111;
assign micromatrizz[12][321] = 9'b111111111;
assign micromatrizz[12][322] = 9'b111111111;
assign micromatrizz[12][323] = 9'b111111111;
assign micromatrizz[12][324] = 9'b111111111;
assign micromatrizz[12][325] = 9'b111111111;
assign micromatrizz[12][326] = 9'b111111111;
assign micromatrizz[12][327] = 9'b111111111;
assign micromatrizz[12][328] = 9'b111111111;
assign micromatrizz[12][329] = 9'b111111111;
assign micromatrizz[12][330] = 9'b111111111;
assign micromatrizz[12][331] = 9'b111111111;
assign micromatrizz[12][332] = 9'b111111111;
assign micromatrizz[12][333] = 9'b111111111;
assign micromatrizz[12][334] = 9'b111111111;
assign micromatrizz[12][335] = 9'b111111111;
assign micromatrizz[12][336] = 9'b111111111;
assign micromatrizz[12][337] = 9'b111111111;
assign micromatrizz[12][338] = 9'b111111111;
assign micromatrizz[12][339] = 9'b111111111;
assign micromatrizz[12][340] = 9'b111111111;
assign micromatrizz[12][341] = 9'b111111111;
assign micromatrizz[12][342] = 9'b111111111;
assign micromatrizz[12][343] = 9'b111111111;
assign micromatrizz[12][344] = 9'b111111111;
assign micromatrizz[12][345] = 9'b111111111;
assign micromatrizz[12][346] = 9'b111111111;
assign micromatrizz[12][347] = 9'b111111111;
assign micromatrizz[12][348] = 9'b111111111;
assign micromatrizz[12][349] = 9'b111111111;
assign micromatrizz[12][350] = 9'b111111111;
assign micromatrizz[12][351] = 9'b111111111;
assign micromatrizz[12][352] = 9'b111111111;
assign micromatrizz[12][353] = 9'b111111111;
assign micromatrizz[12][354] = 9'b111111111;
assign micromatrizz[12][355] = 9'b111111111;
assign micromatrizz[12][356] = 9'b111111111;
assign micromatrizz[12][357] = 9'b111111111;
assign micromatrizz[12][358] = 9'b111111111;
assign micromatrizz[12][359] = 9'b111111111;
assign micromatrizz[12][360] = 9'b111111111;
assign micromatrizz[12][361] = 9'b111111111;
assign micromatrizz[12][362] = 9'b111111111;
assign micromatrizz[12][363] = 9'b111111111;
assign micromatrizz[12][364] = 9'b111111111;
assign micromatrizz[12][365] = 9'b111111111;
assign micromatrizz[12][366] = 9'b111111111;
assign micromatrizz[12][367] = 9'b111111111;
assign micromatrizz[12][368] = 9'b111111111;
assign micromatrizz[12][369] = 9'b111111111;
assign micromatrizz[12][370] = 9'b111111111;
assign micromatrizz[12][371] = 9'b111111111;
assign micromatrizz[12][372] = 9'b111111111;
assign micromatrizz[12][373] = 9'b111111111;
assign micromatrizz[12][374] = 9'b111111111;
assign micromatrizz[12][375] = 9'b111111111;
assign micromatrizz[12][376] = 9'b111111111;
assign micromatrizz[12][377] = 9'b111111111;
assign micromatrizz[12][378] = 9'b111111111;
assign micromatrizz[12][379] = 9'b111111111;
assign micromatrizz[12][380] = 9'b111111111;
assign micromatrizz[12][381] = 9'b111111111;
assign micromatrizz[12][382] = 9'b111111111;
assign micromatrizz[12][383] = 9'b111111111;
assign micromatrizz[12][384] = 9'b111111111;
assign micromatrizz[12][385] = 9'b111111111;
assign micromatrizz[12][386] = 9'b111111111;
assign micromatrizz[12][387] = 9'b111111111;
assign micromatrizz[12][388] = 9'b111111111;
assign micromatrizz[12][389] = 9'b111111111;
assign micromatrizz[12][390] = 9'b111111111;
assign micromatrizz[12][391] = 9'b111111111;
assign micromatrizz[12][392] = 9'b111111111;
assign micromatrizz[12][393] = 9'b111111111;
assign micromatrizz[12][394] = 9'b111111111;
assign micromatrizz[12][395] = 9'b111111111;
assign micromatrizz[12][396] = 9'b111111111;
assign micromatrizz[12][397] = 9'b111111111;
assign micromatrizz[12][398] = 9'b111111111;
assign micromatrizz[12][399] = 9'b111111111;
assign micromatrizz[12][400] = 9'b111111111;
assign micromatrizz[12][401] = 9'b111111111;
assign micromatrizz[12][402] = 9'b111111111;
assign micromatrizz[12][403] = 9'b111111111;
assign micromatrizz[12][404] = 9'b111111111;
assign micromatrizz[12][405] = 9'b111111111;
assign micromatrizz[12][406] = 9'b111111111;
assign micromatrizz[12][407] = 9'b111111111;
assign micromatrizz[12][408] = 9'b111111111;
assign micromatrizz[12][409] = 9'b111111111;
assign micromatrizz[12][410] = 9'b111111111;
assign micromatrizz[12][411] = 9'b111111111;
assign micromatrizz[12][412] = 9'b111111111;
assign micromatrizz[12][413] = 9'b111111111;
assign micromatrizz[12][414] = 9'b111111111;
assign micromatrizz[12][415] = 9'b111111111;
assign micromatrizz[12][416] = 9'b111111111;
assign micromatrizz[12][417] = 9'b111111111;
assign micromatrizz[12][418] = 9'b111111111;
assign micromatrizz[12][419] = 9'b111111111;
assign micromatrizz[12][420] = 9'b111111111;
assign micromatrizz[12][421] = 9'b111111111;
assign micromatrizz[12][422] = 9'b111111111;
assign micromatrizz[12][423] = 9'b111111111;
assign micromatrizz[12][424] = 9'b111111111;
assign micromatrizz[12][425] = 9'b111111111;
assign micromatrizz[12][426] = 9'b111111111;
assign micromatrizz[12][427] = 9'b111111111;
assign micromatrizz[12][428] = 9'b111111111;
assign micromatrizz[12][429] = 9'b111111111;
assign micromatrizz[12][430] = 9'b111111111;
assign micromatrizz[12][431] = 9'b111111111;
assign micromatrizz[12][432] = 9'b111111111;
assign micromatrizz[12][433] = 9'b111111111;
assign micromatrizz[12][434] = 9'b111111111;
assign micromatrizz[12][435] = 9'b111111111;
assign micromatrizz[12][436] = 9'b111111111;
assign micromatrizz[12][437] = 9'b111111111;
assign micromatrizz[12][438] = 9'b111111111;
assign micromatrizz[12][439] = 9'b111111111;
assign micromatrizz[12][440] = 9'b111111111;
assign micromatrizz[12][441] = 9'b111111111;
assign micromatrizz[12][442] = 9'b111111111;
assign micromatrizz[12][443] = 9'b111111111;
assign micromatrizz[12][444] = 9'b111111111;
assign micromatrizz[12][445] = 9'b111111111;
assign micromatrizz[12][446] = 9'b111111111;
assign micromatrizz[12][447] = 9'b111111111;
assign micromatrizz[12][448] = 9'b111111111;
assign micromatrizz[12][449] = 9'b111111111;
assign micromatrizz[12][450] = 9'b111111111;
assign micromatrizz[12][451] = 9'b111111111;
assign micromatrizz[12][452] = 9'b111111111;
assign micromatrizz[12][453] = 9'b111111111;
assign micromatrizz[12][454] = 9'b111111111;
assign micromatrizz[12][455] = 9'b111111111;
assign micromatrizz[12][456] = 9'b111111111;
assign micromatrizz[12][457] = 9'b111111111;
assign micromatrizz[12][458] = 9'b111111111;
assign micromatrizz[12][459] = 9'b111111111;
assign micromatrizz[12][460] = 9'b111111111;
assign micromatrizz[12][461] = 9'b111111111;
assign micromatrizz[12][462] = 9'b111111111;
assign micromatrizz[12][463] = 9'b111111111;
assign micromatrizz[12][464] = 9'b111111111;
assign micromatrizz[12][465] = 9'b111111111;
assign micromatrizz[12][466] = 9'b111111111;
assign micromatrizz[12][467] = 9'b111111111;
assign micromatrizz[12][468] = 9'b111111111;
assign micromatrizz[12][469] = 9'b111111111;
assign micromatrizz[12][470] = 9'b111111111;
assign micromatrizz[12][471] = 9'b111111111;
assign micromatrizz[12][472] = 9'b111111111;
assign micromatrizz[12][473] = 9'b111111111;
assign micromatrizz[12][474] = 9'b111111111;
assign micromatrizz[12][475] = 9'b111111111;
assign micromatrizz[12][476] = 9'b111111111;
assign micromatrizz[12][477] = 9'b111111111;
assign micromatrizz[12][478] = 9'b111111111;
assign micromatrizz[12][479] = 9'b111111111;
assign micromatrizz[12][480] = 9'b111111111;
assign micromatrizz[12][481] = 9'b111111111;
assign micromatrizz[12][482] = 9'b111111111;
assign micromatrizz[12][483] = 9'b111111111;
assign micromatrizz[12][484] = 9'b111111111;
assign micromatrizz[12][485] = 9'b111111111;
assign micromatrizz[12][486] = 9'b111111111;
assign micromatrizz[12][487] = 9'b111111111;
assign micromatrizz[12][488] = 9'b111111111;
assign micromatrizz[12][489] = 9'b111111111;
assign micromatrizz[12][490] = 9'b111111111;
assign micromatrizz[12][491] = 9'b111111111;
assign micromatrizz[12][492] = 9'b111111111;
assign micromatrizz[12][493] = 9'b111111111;
assign micromatrizz[12][494] = 9'b111111111;
assign micromatrizz[12][495] = 9'b111111111;
assign micromatrizz[12][496] = 9'b111111111;
assign micromatrizz[12][497] = 9'b111111111;
assign micromatrizz[12][498] = 9'b111111111;
assign micromatrizz[12][499] = 9'b111111111;
assign micromatrizz[12][500] = 9'b111111111;
assign micromatrizz[12][501] = 9'b111111111;
assign micromatrizz[12][502] = 9'b111111111;
assign micromatrizz[12][503] = 9'b111111111;
assign micromatrizz[12][504] = 9'b111111111;
assign micromatrizz[12][505] = 9'b111111111;
assign micromatrizz[12][506] = 9'b111111111;
assign micromatrizz[12][507] = 9'b111111111;
assign micromatrizz[12][508] = 9'b111111111;
assign micromatrizz[12][509] = 9'b111111111;
assign micromatrizz[12][510] = 9'b111111111;
assign micromatrizz[12][511] = 9'b111111111;
assign micromatrizz[12][512] = 9'b111111111;
assign micromatrizz[12][513] = 9'b111111111;
assign micromatrizz[12][514] = 9'b111111111;
assign micromatrizz[12][515] = 9'b111111111;
assign micromatrizz[12][516] = 9'b111111111;
assign micromatrizz[12][517] = 9'b111111111;
assign micromatrizz[12][518] = 9'b111111111;
assign micromatrizz[12][519] = 9'b111111111;
assign micromatrizz[12][520] = 9'b111111111;
assign micromatrizz[12][521] = 9'b111111111;
assign micromatrizz[12][522] = 9'b111111111;
assign micromatrizz[12][523] = 9'b111111111;
assign micromatrizz[12][524] = 9'b111111111;
assign micromatrizz[12][525] = 9'b111111111;
assign micromatrizz[12][526] = 9'b111111111;
assign micromatrizz[12][527] = 9'b111111111;
assign micromatrizz[12][528] = 9'b111111111;
assign micromatrizz[12][529] = 9'b111111111;
assign micromatrizz[12][530] = 9'b111111111;
assign micromatrizz[12][531] = 9'b111111111;
assign micromatrizz[12][532] = 9'b111111111;
assign micromatrizz[12][533] = 9'b111111111;
assign micromatrizz[12][534] = 9'b111111111;
assign micromatrizz[12][535] = 9'b111111111;
assign micromatrizz[12][536] = 9'b111111111;
assign micromatrizz[12][537] = 9'b111111111;
assign micromatrizz[12][538] = 9'b111111111;
assign micromatrizz[12][539] = 9'b111111111;
assign micromatrizz[12][540] = 9'b111111111;
assign micromatrizz[12][541] = 9'b111111111;
assign micromatrizz[12][542] = 9'b111111111;
assign micromatrizz[12][543] = 9'b111111111;
assign micromatrizz[12][544] = 9'b111111111;
assign micromatrizz[12][545] = 9'b111111111;
assign micromatrizz[12][546] = 9'b111111111;
assign micromatrizz[12][547] = 9'b111111111;
assign micromatrizz[12][548] = 9'b111111111;
assign micromatrizz[12][549] = 9'b111111111;
assign micromatrizz[12][550] = 9'b111111111;
assign micromatrizz[12][551] = 9'b111111111;
assign micromatrizz[12][552] = 9'b111111111;
assign micromatrizz[12][553] = 9'b111111111;
assign micromatrizz[12][554] = 9'b111111111;
assign micromatrizz[12][555] = 9'b111111111;
assign micromatrizz[12][556] = 9'b111111111;
assign micromatrizz[12][557] = 9'b111111111;
assign micromatrizz[12][558] = 9'b111111111;
assign micromatrizz[12][559] = 9'b111111111;
assign micromatrizz[12][560] = 9'b111111111;
assign micromatrizz[12][561] = 9'b111111111;
assign micromatrizz[12][562] = 9'b111111111;
assign micromatrizz[12][563] = 9'b111111111;
assign micromatrizz[12][564] = 9'b111111111;
assign micromatrizz[12][565] = 9'b111111111;
assign micromatrizz[12][566] = 9'b111111111;
assign micromatrizz[12][567] = 9'b111111111;
assign micromatrizz[12][568] = 9'b111111111;
assign micromatrizz[12][569] = 9'b111111111;
assign micromatrizz[12][570] = 9'b111111111;
assign micromatrizz[12][571] = 9'b111111111;
assign micromatrizz[12][572] = 9'b111111111;
assign micromatrizz[12][573] = 9'b111111111;
assign micromatrizz[12][574] = 9'b111111111;
assign micromatrizz[12][575] = 9'b111111111;
assign micromatrizz[12][576] = 9'b111111111;
assign micromatrizz[12][577] = 9'b111111111;
assign micromatrizz[12][578] = 9'b111111111;
assign micromatrizz[12][579] = 9'b111111111;
assign micromatrizz[12][580] = 9'b111111111;
assign micromatrizz[12][581] = 9'b111111111;
assign micromatrizz[12][582] = 9'b111111111;
assign micromatrizz[12][583] = 9'b111111111;
assign micromatrizz[12][584] = 9'b111111111;
assign micromatrizz[12][585] = 9'b111111111;
assign micromatrizz[12][586] = 9'b111111111;
assign micromatrizz[12][587] = 9'b111111111;
assign micromatrizz[12][588] = 9'b111111111;
assign micromatrizz[12][589] = 9'b111111111;
assign micromatrizz[12][590] = 9'b111111111;
assign micromatrizz[12][591] = 9'b111111111;
assign micromatrizz[12][592] = 9'b111111111;
assign micromatrizz[12][593] = 9'b111111111;
assign micromatrizz[12][594] = 9'b111111111;
assign micromatrizz[12][595] = 9'b111111111;
assign micromatrizz[12][596] = 9'b111111111;
assign micromatrizz[12][597] = 9'b111111111;
assign micromatrizz[12][598] = 9'b111111111;
assign micromatrizz[12][599] = 9'b111111111;
assign micromatrizz[12][600] = 9'b111111111;
assign micromatrizz[12][601] = 9'b111111111;
assign micromatrizz[12][602] = 9'b111111111;
assign micromatrizz[12][603] = 9'b111111111;
assign micromatrizz[12][604] = 9'b111111111;
assign micromatrizz[12][605] = 9'b111111111;
assign micromatrizz[12][606] = 9'b111111111;
assign micromatrizz[12][607] = 9'b111111111;
assign micromatrizz[12][608] = 9'b111111111;
assign micromatrizz[12][609] = 9'b111111111;
assign micromatrizz[12][610] = 9'b111111111;
assign micromatrizz[12][611] = 9'b111111111;
assign micromatrizz[12][612] = 9'b111111111;
assign micromatrizz[12][613] = 9'b111111111;
assign micromatrizz[12][614] = 9'b111111111;
assign micromatrizz[12][615] = 9'b111111111;
assign micromatrizz[12][616] = 9'b111111111;
assign micromatrizz[12][617] = 9'b111111111;
assign micromatrizz[12][618] = 9'b111111111;
assign micromatrizz[12][619] = 9'b111111111;
assign micromatrizz[12][620] = 9'b111111111;
assign micromatrizz[12][621] = 9'b111111111;
assign micromatrizz[12][622] = 9'b111111111;
assign micromatrizz[12][623] = 9'b111111111;
assign micromatrizz[12][624] = 9'b111111111;
assign micromatrizz[12][625] = 9'b111111111;
assign micromatrizz[12][626] = 9'b111111111;
assign micromatrizz[12][627] = 9'b111111111;
assign micromatrizz[12][628] = 9'b111111111;
assign micromatrizz[12][629] = 9'b111111111;
assign micromatrizz[12][630] = 9'b111111111;
assign micromatrizz[12][631] = 9'b111111111;
assign micromatrizz[12][632] = 9'b111111111;
assign micromatrizz[12][633] = 9'b111111111;
assign micromatrizz[12][634] = 9'b111111111;
assign micromatrizz[12][635] = 9'b111111111;
assign micromatrizz[12][636] = 9'b111111111;
assign micromatrizz[12][637] = 9'b111111111;
assign micromatrizz[12][638] = 9'b111111111;
assign micromatrizz[12][639] = 9'b111111111;
assign micromatrizz[13][0] = 9'b111111111;
assign micromatrizz[13][1] = 9'b111111111;
assign micromatrizz[13][2] = 9'b111111111;
assign micromatrizz[13][3] = 9'b111111111;
assign micromatrizz[13][4] = 9'b111111111;
assign micromatrizz[13][5] = 9'b111111111;
assign micromatrizz[13][6] = 9'b111111111;
assign micromatrizz[13][7] = 9'b111111111;
assign micromatrizz[13][8] = 9'b111111111;
assign micromatrizz[13][9] = 9'b111111111;
assign micromatrizz[13][10] = 9'b111111111;
assign micromatrizz[13][11] = 9'b111111111;
assign micromatrizz[13][12] = 9'b111111111;
assign micromatrizz[13][13] = 9'b111111111;
assign micromatrizz[13][14] = 9'b111111111;
assign micromatrizz[13][15] = 9'b111111111;
assign micromatrizz[13][16] = 9'b111111111;
assign micromatrizz[13][17] = 9'b111111111;
assign micromatrizz[13][18] = 9'b111111111;
assign micromatrizz[13][19] = 9'b111111111;
assign micromatrizz[13][20] = 9'b111111111;
assign micromatrizz[13][21] = 9'b111111111;
assign micromatrizz[13][22] = 9'b111111111;
assign micromatrizz[13][23] = 9'b111111111;
assign micromatrizz[13][24] = 9'b111111111;
assign micromatrizz[13][25] = 9'b111111111;
assign micromatrizz[13][26] = 9'b111111111;
assign micromatrizz[13][27] = 9'b111111111;
assign micromatrizz[13][28] = 9'b111111111;
assign micromatrizz[13][29] = 9'b111111111;
assign micromatrizz[13][30] = 9'b111111111;
assign micromatrizz[13][31] = 9'b111111111;
assign micromatrizz[13][32] = 9'b111111111;
assign micromatrizz[13][33] = 9'b111111111;
assign micromatrizz[13][34] = 9'b111111111;
assign micromatrizz[13][35] = 9'b111111111;
assign micromatrizz[13][36] = 9'b111111111;
assign micromatrizz[13][37] = 9'b111111111;
assign micromatrizz[13][38] = 9'b111111111;
assign micromatrizz[13][39] = 9'b111111111;
assign micromatrizz[13][40] = 9'b111111111;
assign micromatrizz[13][41] = 9'b111111111;
assign micromatrizz[13][42] = 9'b111111111;
assign micromatrizz[13][43] = 9'b111111111;
assign micromatrizz[13][44] = 9'b111111111;
assign micromatrizz[13][45] = 9'b111111111;
assign micromatrizz[13][46] = 9'b111111111;
assign micromatrizz[13][47] = 9'b111111111;
assign micromatrizz[13][48] = 9'b111111111;
assign micromatrizz[13][49] = 9'b111111111;
assign micromatrizz[13][50] = 9'b111111111;
assign micromatrizz[13][51] = 9'b111111111;
assign micromatrizz[13][52] = 9'b111111111;
assign micromatrizz[13][53] = 9'b111111111;
assign micromatrizz[13][54] = 9'b111111111;
assign micromatrizz[13][55] = 9'b111111111;
assign micromatrizz[13][56] = 9'b111111111;
assign micromatrizz[13][57] = 9'b111111111;
assign micromatrizz[13][58] = 9'b111111111;
assign micromatrizz[13][59] = 9'b111111111;
assign micromatrizz[13][60] = 9'b111111111;
assign micromatrizz[13][61] = 9'b111111111;
assign micromatrizz[13][62] = 9'b111111111;
assign micromatrizz[13][63] = 9'b111111111;
assign micromatrizz[13][64] = 9'b111111111;
assign micromatrizz[13][65] = 9'b111111111;
assign micromatrizz[13][66] = 9'b111111111;
assign micromatrizz[13][67] = 9'b111111111;
assign micromatrizz[13][68] = 9'b111111111;
assign micromatrizz[13][69] = 9'b111111111;
assign micromatrizz[13][70] = 9'b111111111;
assign micromatrizz[13][71] = 9'b111111111;
assign micromatrizz[13][72] = 9'b111111111;
assign micromatrizz[13][73] = 9'b111111111;
assign micromatrizz[13][74] = 9'b111111111;
assign micromatrizz[13][75] = 9'b111111111;
assign micromatrizz[13][76] = 9'b111111111;
assign micromatrizz[13][77] = 9'b111111111;
assign micromatrizz[13][78] = 9'b111111111;
assign micromatrizz[13][79] = 9'b111111111;
assign micromatrizz[13][80] = 9'b111111111;
assign micromatrizz[13][81] = 9'b111111111;
assign micromatrizz[13][82] = 9'b111111111;
assign micromatrizz[13][83] = 9'b111111111;
assign micromatrizz[13][84] = 9'b111111111;
assign micromatrizz[13][85] = 9'b111111111;
assign micromatrizz[13][86] = 9'b111111111;
assign micromatrizz[13][87] = 9'b111111111;
assign micromatrizz[13][88] = 9'b111111111;
assign micromatrizz[13][89] = 9'b111111111;
assign micromatrizz[13][90] = 9'b111111111;
assign micromatrizz[13][91] = 9'b111111111;
assign micromatrizz[13][92] = 9'b111111111;
assign micromatrizz[13][93] = 9'b111111111;
assign micromatrizz[13][94] = 9'b111111111;
assign micromatrizz[13][95] = 9'b111111111;
assign micromatrizz[13][96] = 9'b111111111;
assign micromatrizz[13][97] = 9'b111111111;
assign micromatrizz[13][98] = 9'b111111111;
assign micromatrizz[13][99] = 9'b111111111;
assign micromatrizz[13][100] = 9'b111111111;
assign micromatrizz[13][101] = 9'b111111111;
assign micromatrizz[13][102] = 9'b111111111;
assign micromatrizz[13][103] = 9'b111111111;
assign micromatrizz[13][104] = 9'b111111111;
assign micromatrizz[13][105] = 9'b111111111;
assign micromatrizz[13][106] = 9'b111111111;
assign micromatrizz[13][107] = 9'b111111111;
assign micromatrizz[13][108] = 9'b111111111;
assign micromatrizz[13][109] = 9'b111111111;
assign micromatrizz[13][110] = 9'b111111111;
assign micromatrizz[13][111] = 9'b111111111;
assign micromatrizz[13][112] = 9'b111111111;
assign micromatrizz[13][113] = 9'b111111111;
assign micromatrizz[13][114] = 9'b111111111;
assign micromatrizz[13][115] = 9'b111111111;
assign micromatrizz[13][116] = 9'b111111111;
assign micromatrizz[13][117] = 9'b111111111;
assign micromatrizz[13][118] = 9'b111111111;
assign micromatrizz[13][119] = 9'b111111111;
assign micromatrizz[13][120] = 9'b111111111;
assign micromatrizz[13][121] = 9'b111111111;
assign micromatrizz[13][122] = 9'b111111111;
assign micromatrizz[13][123] = 9'b111111111;
assign micromatrizz[13][124] = 9'b111111111;
assign micromatrizz[13][125] = 9'b111111111;
assign micromatrizz[13][126] = 9'b111111111;
assign micromatrizz[13][127] = 9'b111111111;
assign micromatrizz[13][128] = 9'b111111111;
assign micromatrizz[13][129] = 9'b111111111;
assign micromatrizz[13][130] = 9'b111111111;
assign micromatrizz[13][131] = 9'b111111111;
assign micromatrizz[13][132] = 9'b111111111;
assign micromatrizz[13][133] = 9'b111111111;
assign micromatrizz[13][134] = 9'b111111111;
assign micromatrizz[13][135] = 9'b111111111;
assign micromatrizz[13][136] = 9'b111111111;
assign micromatrizz[13][137] = 9'b111111111;
assign micromatrizz[13][138] = 9'b111111111;
assign micromatrizz[13][139] = 9'b111111111;
assign micromatrizz[13][140] = 9'b111111111;
assign micromatrizz[13][141] = 9'b111111111;
assign micromatrizz[13][142] = 9'b111111111;
assign micromatrizz[13][143] = 9'b111111111;
assign micromatrizz[13][144] = 9'b111111111;
assign micromatrizz[13][145] = 9'b111111111;
assign micromatrizz[13][146] = 9'b111111111;
assign micromatrizz[13][147] = 9'b111111111;
assign micromatrizz[13][148] = 9'b111111111;
assign micromatrizz[13][149] = 9'b111111111;
assign micromatrizz[13][150] = 9'b111111111;
assign micromatrizz[13][151] = 9'b111111111;
assign micromatrizz[13][152] = 9'b111111111;
assign micromatrizz[13][153] = 9'b111111111;
assign micromatrizz[13][154] = 9'b111111111;
assign micromatrizz[13][155] = 9'b111111111;
assign micromatrizz[13][156] = 9'b111111111;
assign micromatrizz[13][157] = 9'b111111111;
assign micromatrizz[13][158] = 9'b111111111;
assign micromatrizz[13][159] = 9'b111111111;
assign micromatrizz[13][160] = 9'b111111111;
assign micromatrizz[13][161] = 9'b111111111;
assign micromatrizz[13][162] = 9'b111111111;
assign micromatrizz[13][163] = 9'b111111111;
assign micromatrizz[13][164] = 9'b111111111;
assign micromatrizz[13][165] = 9'b111111111;
assign micromatrizz[13][166] = 9'b111111111;
assign micromatrizz[13][167] = 9'b111111111;
assign micromatrizz[13][168] = 9'b111111111;
assign micromatrizz[13][169] = 9'b111111111;
assign micromatrizz[13][170] = 9'b111111111;
assign micromatrizz[13][171] = 9'b111111111;
assign micromatrizz[13][172] = 9'b111111111;
assign micromatrizz[13][173] = 9'b111111111;
assign micromatrizz[13][174] = 9'b111111111;
assign micromatrizz[13][175] = 9'b111111111;
assign micromatrizz[13][176] = 9'b111111111;
assign micromatrizz[13][177] = 9'b111111111;
assign micromatrizz[13][178] = 9'b111111111;
assign micromatrizz[13][179] = 9'b111111111;
assign micromatrizz[13][180] = 9'b111111111;
assign micromatrizz[13][181] = 9'b111111111;
assign micromatrizz[13][182] = 9'b111111111;
assign micromatrizz[13][183] = 9'b111111111;
assign micromatrizz[13][184] = 9'b111111111;
assign micromatrizz[13][185] = 9'b111111111;
assign micromatrizz[13][186] = 9'b111111111;
assign micromatrizz[13][187] = 9'b111111111;
assign micromatrizz[13][188] = 9'b111111111;
assign micromatrizz[13][189] = 9'b111111111;
assign micromatrizz[13][190] = 9'b111111111;
assign micromatrizz[13][191] = 9'b111111111;
assign micromatrizz[13][192] = 9'b111111111;
assign micromatrizz[13][193] = 9'b111111111;
assign micromatrizz[13][194] = 9'b111111111;
assign micromatrizz[13][195] = 9'b111111111;
assign micromatrizz[13][196] = 9'b111111111;
assign micromatrizz[13][197] = 9'b111111111;
assign micromatrizz[13][198] = 9'b111111111;
assign micromatrizz[13][199] = 9'b111111111;
assign micromatrizz[13][200] = 9'b111111111;
assign micromatrizz[13][201] = 9'b111111111;
assign micromatrizz[13][202] = 9'b111111111;
assign micromatrizz[13][203] = 9'b111111111;
assign micromatrizz[13][204] = 9'b111111111;
assign micromatrizz[13][205] = 9'b111111111;
assign micromatrizz[13][206] = 9'b111111111;
assign micromatrizz[13][207] = 9'b111111111;
assign micromatrizz[13][208] = 9'b111111111;
assign micromatrizz[13][209] = 9'b111111111;
assign micromatrizz[13][210] = 9'b111111111;
assign micromatrizz[13][211] = 9'b111111111;
assign micromatrizz[13][212] = 9'b111111111;
assign micromatrizz[13][213] = 9'b111111111;
assign micromatrizz[13][214] = 9'b111111111;
assign micromatrizz[13][215] = 9'b111111111;
assign micromatrizz[13][216] = 9'b111111111;
assign micromatrizz[13][217] = 9'b111111111;
assign micromatrizz[13][218] = 9'b111111111;
assign micromatrizz[13][219] = 9'b111111111;
assign micromatrizz[13][220] = 9'b111111111;
assign micromatrizz[13][221] = 9'b111111111;
assign micromatrizz[13][222] = 9'b111111111;
assign micromatrizz[13][223] = 9'b111111111;
assign micromatrizz[13][224] = 9'b111111111;
assign micromatrizz[13][225] = 9'b111111111;
assign micromatrizz[13][226] = 9'b111111111;
assign micromatrizz[13][227] = 9'b111111111;
assign micromatrizz[13][228] = 9'b111111111;
assign micromatrizz[13][229] = 9'b111111111;
assign micromatrizz[13][230] = 9'b111111111;
assign micromatrizz[13][231] = 9'b111111111;
assign micromatrizz[13][232] = 9'b111111111;
assign micromatrizz[13][233] = 9'b111111111;
assign micromatrizz[13][234] = 9'b111111111;
assign micromatrizz[13][235] = 9'b111111111;
assign micromatrizz[13][236] = 9'b111111111;
assign micromatrizz[13][237] = 9'b111111111;
assign micromatrizz[13][238] = 9'b111111111;
assign micromatrizz[13][239] = 9'b111111111;
assign micromatrizz[13][240] = 9'b111111111;
assign micromatrizz[13][241] = 9'b111111111;
assign micromatrizz[13][242] = 9'b111111111;
assign micromatrizz[13][243] = 9'b111111111;
assign micromatrizz[13][244] = 9'b111111111;
assign micromatrizz[13][245] = 9'b111111111;
assign micromatrizz[13][246] = 9'b111111111;
assign micromatrizz[13][247] = 9'b111111111;
assign micromatrizz[13][248] = 9'b111111111;
assign micromatrizz[13][249] = 9'b111111111;
assign micromatrizz[13][250] = 9'b111111111;
assign micromatrizz[13][251] = 9'b111111111;
assign micromatrizz[13][252] = 9'b111111111;
assign micromatrizz[13][253] = 9'b111111111;
assign micromatrizz[13][254] = 9'b111111111;
assign micromatrizz[13][255] = 9'b111111111;
assign micromatrizz[13][256] = 9'b111111111;
assign micromatrizz[13][257] = 9'b111111111;
assign micromatrizz[13][258] = 9'b111111111;
assign micromatrizz[13][259] = 9'b111111111;
assign micromatrizz[13][260] = 9'b111111111;
assign micromatrizz[13][261] = 9'b111111111;
assign micromatrizz[13][262] = 9'b111111111;
assign micromatrizz[13][263] = 9'b111111111;
assign micromatrizz[13][264] = 9'b111111111;
assign micromatrizz[13][265] = 9'b111111111;
assign micromatrizz[13][266] = 9'b111111111;
assign micromatrizz[13][267] = 9'b111111111;
assign micromatrizz[13][268] = 9'b111111111;
assign micromatrizz[13][269] = 9'b111111111;
assign micromatrizz[13][270] = 9'b111111111;
assign micromatrizz[13][271] = 9'b111111111;
assign micromatrizz[13][272] = 9'b111111111;
assign micromatrizz[13][273] = 9'b111111111;
assign micromatrizz[13][274] = 9'b111111111;
assign micromatrizz[13][275] = 9'b111111111;
assign micromatrizz[13][276] = 9'b111111111;
assign micromatrizz[13][277] = 9'b111111111;
assign micromatrizz[13][278] = 9'b111111111;
assign micromatrizz[13][279] = 9'b111111111;
assign micromatrizz[13][280] = 9'b111111111;
assign micromatrizz[13][281] = 9'b111111111;
assign micromatrizz[13][282] = 9'b111111111;
assign micromatrizz[13][283] = 9'b111111111;
assign micromatrizz[13][284] = 9'b111111111;
assign micromatrizz[13][285] = 9'b111111111;
assign micromatrizz[13][286] = 9'b111111111;
assign micromatrizz[13][287] = 9'b111111111;
assign micromatrizz[13][288] = 9'b111111111;
assign micromatrizz[13][289] = 9'b111111111;
assign micromatrizz[13][290] = 9'b111111111;
assign micromatrizz[13][291] = 9'b111111111;
assign micromatrizz[13][292] = 9'b111111111;
assign micromatrizz[13][293] = 9'b111111111;
assign micromatrizz[13][294] = 9'b111111111;
assign micromatrizz[13][295] = 9'b111111111;
assign micromatrizz[13][296] = 9'b111111111;
assign micromatrizz[13][297] = 9'b111111111;
assign micromatrizz[13][298] = 9'b111111111;
assign micromatrizz[13][299] = 9'b111111111;
assign micromatrizz[13][300] = 9'b111111111;
assign micromatrizz[13][301] = 9'b111111111;
assign micromatrizz[13][302] = 9'b111111111;
assign micromatrizz[13][303] = 9'b111111111;
assign micromatrizz[13][304] = 9'b111111111;
assign micromatrizz[13][305] = 9'b111111111;
assign micromatrizz[13][306] = 9'b111111111;
assign micromatrizz[13][307] = 9'b111111111;
assign micromatrizz[13][308] = 9'b111111111;
assign micromatrizz[13][309] = 9'b111111111;
assign micromatrizz[13][310] = 9'b111111111;
assign micromatrizz[13][311] = 9'b111111111;
assign micromatrizz[13][312] = 9'b111111111;
assign micromatrizz[13][313] = 9'b111111111;
assign micromatrizz[13][314] = 9'b111111111;
assign micromatrizz[13][315] = 9'b111111111;
assign micromatrizz[13][316] = 9'b111111111;
assign micromatrizz[13][317] = 9'b111111111;
assign micromatrizz[13][318] = 9'b111111111;
assign micromatrizz[13][319] = 9'b111111111;
assign micromatrizz[13][320] = 9'b111111111;
assign micromatrizz[13][321] = 9'b111111111;
assign micromatrizz[13][322] = 9'b111111111;
assign micromatrizz[13][323] = 9'b111111111;
assign micromatrizz[13][324] = 9'b111111111;
assign micromatrizz[13][325] = 9'b111111111;
assign micromatrizz[13][326] = 9'b111111111;
assign micromatrizz[13][327] = 9'b111111111;
assign micromatrizz[13][328] = 9'b111111111;
assign micromatrizz[13][329] = 9'b111111111;
assign micromatrizz[13][330] = 9'b111111111;
assign micromatrizz[13][331] = 9'b111111111;
assign micromatrizz[13][332] = 9'b111111111;
assign micromatrizz[13][333] = 9'b111111111;
assign micromatrizz[13][334] = 9'b111111111;
assign micromatrizz[13][335] = 9'b111111111;
assign micromatrizz[13][336] = 9'b111111111;
assign micromatrizz[13][337] = 9'b111111111;
assign micromatrizz[13][338] = 9'b111111111;
assign micromatrizz[13][339] = 9'b111111111;
assign micromatrizz[13][340] = 9'b111111111;
assign micromatrizz[13][341] = 9'b111111111;
assign micromatrizz[13][342] = 9'b111111111;
assign micromatrizz[13][343] = 9'b111111111;
assign micromatrizz[13][344] = 9'b111111111;
assign micromatrizz[13][345] = 9'b111111111;
assign micromatrizz[13][346] = 9'b111111111;
assign micromatrizz[13][347] = 9'b111111111;
assign micromatrizz[13][348] = 9'b111111111;
assign micromatrizz[13][349] = 9'b111111111;
assign micromatrizz[13][350] = 9'b111111111;
assign micromatrizz[13][351] = 9'b111111111;
assign micromatrizz[13][352] = 9'b111111111;
assign micromatrizz[13][353] = 9'b111111111;
assign micromatrizz[13][354] = 9'b111111111;
assign micromatrizz[13][355] = 9'b111111111;
assign micromatrizz[13][356] = 9'b111111111;
assign micromatrizz[13][357] = 9'b111111111;
assign micromatrizz[13][358] = 9'b111111111;
assign micromatrizz[13][359] = 9'b111111111;
assign micromatrizz[13][360] = 9'b111111111;
assign micromatrizz[13][361] = 9'b111111111;
assign micromatrizz[13][362] = 9'b111111111;
assign micromatrizz[13][363] = 9'b111111111;
assign micromatrizz[13][364] = 9'b111111111;
assign micromatrizz[13][365] = 9'b111111111;
assign micromatrizz[13][366] = 9'b111111111;
assign micromatrizz[13][367] = 9'b111111111;
assign micromatrizz[13][368] = 9'b111111111;
assign micromatrizz[13][369] = 9'b111111111;
assign micromatrizz[13][370] = 9'b111111111;
assign micromatrizz[13][371] = 9'b111111111;
assign micromatrizz[13][372] = 9'b111111111;
assign micromatrizz[13][373] = 9'b111111111;
assign micromatrizz[13][374] = 9'b111111111;
assign micromatrizz[13][375] = 9'b111111111;
assign micromatrizz[13][376] = 9'b111111111;
assign micromatrizz[13][377] = 9'b111111111;
assign micromatrizz[13][378] = 9'b111111111;
assign micromatrizz[13][379] = 9'b111111111;
assign micromatrizz[13][380] = 9'b111111111;
assign micromatrizz[13][381] = 9'b111111111;
assign micromatrizz[13][382] = 9'b111111111;
assign micromatrizz[13][383] = 9'b111111111;
assign micromatrizz[13][384] = 9'b111111111;
assign micromatrizz[13][385] = 9'b111111111;
assign micromatrizz[13][386] = 9'b111111111;
assign micromatrizz[13][387] = 9'b111111111;
assign micromatrizz[13][388] = 9'b111111111;
assign micromatrizz[13][389] = 9'b111111111;
assign micromatrizz[13][390] = 9'b111111111;
assign micromatrizz[13][391] = 9'b111111111;
assign micromatrizz[13][392] = 9'b111111111;
assign micromatrizz[13][393] = 9'b111111111;
assign micromatrizz[13][394] = 9'b111111111;
assign micromatrizz[13][395] = 9'b111111111;
assign micromatrizz[13][396] = 9'b111111111;
assign micromatrizz[13][397] = 9'b111111111;
assign micromatrizz[13][398] = 9'b111111111;
assign micromatrizz[13][399] = 9'b111111111;
assign micromatrizz[13][400] = 9'b111111111;
assign micromatrizz[13][401] = 9'b111111111;
assign micromatrizz[13][402] = 9'b111111111;
assign micromatrizz[13][403] = 9'b111111111;
assign micromatrizz[13][404] = 9'b111111111;
assign micromatrizz[13][405] = 9'b111111111;
assign micromatrizz[13][406] = 9'b111111111;
assign micromatrizz[13][407] = 9'b111111111;
assign micromatrizz[13][408] = 9'b111111111;
assign micromatrizz[13][409] = 9'b111111111;
assign micromatrizz[13][410] = 9'b111111111;
assign micromatrizz[13][411] = 9'b111111111;
assign micromatrizz[13][412] = 9'b111111111;
assign micromatrizz[13][413] = 9'b111111111;
assign micromatrizz[13][414] = 9'b111111111;
assign micromatrizz[13][415] = 9'b111111111;
assign micromatrizz[13][416] = 9'b111111111;
assign micromatrizz[13][417] = 9'b111111111;
assign micromatrizz[13][418] = 9'b111111111;
assign micromatrizz[13][419] = 9'b111111111;
assign micromatrizz[13][420] = 9'b111111111;
assign micromatrizz[13][421] = 9'b111111111;
assign micromatrizz[13][422] = 9'b111111111;
assign micromatrizz[13][423] = 9'b111111111;
assign micromatrizz[13][424] = 9'b111111111;
assign micromatrizz[13][425] = 9'b111111111;
assign micromatrizz[13][426] = 9'b111111111;
assign micromatrizz[13][427] = 9'b111111111;
assign micromatrizz[13][428] = 9'b111111111;
assign micromatrizz[13][429] = 9'b111111111;
assign micromatrizz[13][430] = 9'b111111111;
assign micromatrizz[13][431] = 9'b111111111;
assign micromatrizz[13][432] = 9'b111111111;
assign micromatrizz[13][433] = 9'b111111111;
assign micromatrizz[13][434] = 9'b111111111;
assign micromatrizz[13][435] = 9'b111111111;
assign micromatrizz[13][436] = 9'b111111111;
assign micromatrizz[13][437] = 9'b111111111;
assign micromatrizz[13][438] = 9'b111111111;
assign micromatrizz[13][439] = 9'b111111111;
assign micromatrizz[13][440] = 9'b111111111;
assign micromatrizz[13][441] = 9'b111111111;
assign micromatrizz[13][442] = 9'b111111111;
assign micromatrizz[13][443] = 9'b111111111;
assign micromatrizz[13][444] = 9'b111111111;
assign micromatrizz[13][445] = 9'b111111111;
assign micromatrizz[13][446] = 9'b111111111;
assign micromatrizz[13][447] = 9'b111111111;
assign micromatrizz[13][448] = 9'b111111111;
assign micromatrizz[13][449] = 9'b111111111;
assign micromatrizz[13][450] = 9'b111111111;
assign micromatrizz[13][451] = 9'b111111111;
assign micromatrizz[13][452] = 9'b111111111;
assign micromatrizz[13][453] = 9'b111111111;
assign micromatrizz[13][454] = 9'b111111111;
assign micromatrizz[13][455] = 9'b111111111;
assign micromatrizz[13][456] = 9'b111111111;
assign micromatrizz[13][457] = 9'b111111111;
assign micromatrizz[13][458] = 9'b111111111;
assign micromatrizz[13][459] = 9'b111111111;
assign micromatrizz[13][460] = 9'b111111111;
assign micromatrizz[13][461] = 9'b111111111;
assign micromatrizz[13][462] = 9'b111111111;
assign micromatrizz[13][463] = 9'b111111111;
assign micromatrizz[13][464] = 9'b111111111;
assign micromatrizz[13][465] = 9'b111111111;
assign micromatrizz[13][466] = 9'b111111111;
assign micromatrizz[13][467] = 9'b111111111;
assign micromatrizz[13][468] = 9'b111111111;
assign micromatrizz[13][469] = 9'b111111111;
assign micromatrizz[13][470] = 9'b111111111;
assign micromatrizz[13][471] = 9'b111111111;
assign micromatrizz[13][472] = 9'b111111111;
assign micromatrizz[13][473] = 9'b111111111;
assign micromatrizz[13][474] = 9'b111111111;
assign micromatrizz[13][475] = 9'b111111111;
assign micromatrizz[13][476] = 9'b111111111;
assign micromatrizz[13][477] = 9'b111111111;
assign micromatrizz[13][478] = 9'b111111111;
assign micromatrizz[13][479] = 9'b111111111;
assign micromatrizz[13][480] = 9'b111111111;
assign micromatrizz[13][481] = 9'b111111111;
assign micromatrizz[13][482] = 9'b111111111;
assign micromatrizz[13][483] = 9'b111111111;
assign micromatrizz[13][484] = 9'b111111111;
assign micromatrizz[13][485] = 9'b111111111;
assign micromatrizz[13][486] = 9'b111111111;
assign micromatrizz[13][487] = 9'b111111111;
assign micromatrizz[13][488] = 9'b111111111;
assign micromatrizz[13][489] = 9'b111111111;
assign micromatrizz[13][490] = 9'b111111111;
assign micromatrizz[13][491] = 9'b111111111;
assign micromatrizz[13][492] = 9'b111111111;
assign micromatrizz[13][493] = 9'b111111111;
assign micromatrizz[13][494] = 9'b111111111;
assign micromatrizz[13][495] = 9'b111111111;
assign micromatrizz[13][496] = 9'b111111111;
assign micromatrizz[13][497] = 9'b111111111;
assign micromatrizz[13][498] = 9'b111111111;
assign micromatrizz[13][499] = 9'b111111111;
assign micromatrizz[13][500] = 9'b111111111;
assign micromatrizz[13][501] = 9'b111111111;
assign micromatrizz[13][502] = 9'b111111111;
assign micromatrizz[13][503] = 9'b111111111;
assign micromatrizz[13][504] = 9'b111111111;
assign micromatrizz[13][505] = 9'b111111111;
assign micromatrizz[13][506] = 9'b111111111;
assign micromatrizz[13][507] = 9'b111111111;
assign micromatrizz[13][508] = 9'b111111111;
assign micromatrizz[13][509] = 9'b111111111;
assign micromatrizz[13][510] = 9'b111111111;
assign micromatrizz[13][511] = 9'b111111111;
assign micromatrizz[13][512] = 9'b111111111;
assign micromatrizz[13][513] = 9'b111111111;
assign micromatrizz[13][514] = 9'b111111111;
assign micromatrizz[13][515] = 9'b111111111;
assign micromatrizz[13][516] = 9'b111111111;
assign micromatrizz[13][517] = 9'b111111111;
assign micromatrizz[13][518] = 9'b111111111;
assign micromatrizz[13][519] = 9'b111111111;
assign micromatrizz[13][520] = 9'b111111111;
assign micromatrizz[13][521] = 9'b111111111;
assign micromatrizz[13][522] = 9'b111111111;
assign micromatrizz[13][523] = 9'b111111111;
assign micromatrizz[13][524] = 9'b111111111;
assign micromatrizz[13][525] = 9'b111111111;
assign micromatrizz[13][526] = 9'b111111111;
assign micromatrizz[13][527] = 9'b111111111;
assign micromatrizz[13][528] = 9'b111111111;
assign micromatrizz[13][529] = 9'b111111111;
assign micromatrizz[13][530] = 9'b111111111;
assign micromatrizz[13][531] = 9'b111111111;
assign micromatrizz[13][532] = 9'b111111111;
assign micromatrizz[13][533] = 9'b111111111;
assign micromatrizz[13][534] = 9'b111111111;
assign micromatrizz[13][535] = 9'b111111111;
assign micromatrizz[13][536] = 9'b111111111;
assign micromatrizz[13][537] = 9'b111111111;
assign micromatrizz[13][538] = 9'b111111111;
assign micromatrizz[13][539] = 9'b111111111;
assign micromatrizz[13][540] = 9'b111111111;
assign micromatrizz[13][541] = 9'b111111111;
assign micromatrizz[13][542] = 9'b111111111;
assign micromatrizz[13][543] = 9'b111111111;
assign micromatrizz[13][544] = 9'b111111111;
assign micromatrizz[13][545] = 9'b111111111;
assign micromatrizz[13][546] = 9'b111111111;
assign micromatrizz[13][547] = 9'b111111111;
assign micromatrizz[13][548] = 9'b111111111;
assign micromatrizz[13][549] = 9'b111111111;
assign micromatrizz[13][550] = 9'b111111111;
assign micromatrizz[13][551] = 9'b111111111;
assign micromatrizz[13][552] = 9'b111111111;
assign micromatrizz[13][553] = 9'b111111111;
assign micromatrizz[13][554] = 9'b111111111;
assign micromatrizz[13][555] = 9'b111111111;
assign micromatrizz[13][556] = 9'b111111111;
assign micromatrizz[13][557] = 9'b111111111;
assign micromatrizz[13][558] = 9'b111111111;
assign micromatrizz[13][559] = 9'b111111111;
assign micromatrizz[13][560] = 9'b111111111;
assign micromatrizz[13][561] = 9'b111111111;
assign micromatrizz[13][562] = 9'b111111111;
assign micromatrizz[13][563] = 9'b111111111;
assign micromatrizz[13][564] = 9'b111111111;
assign micromatrizz[13][565] = 9'b111111111;
assign micromatrizz[13][566] = 9'b111111111;
assign micromatrizz[13][567] = 9'b111111111;
assign micromatrizz[13][568] = 9'b111111111;
assign micromatrizz[13][569] = 9'b111111111;
assign micromatrizz[13][570] = 9'b111111111;
assign micromatrizz[13][571] = 9'b111111111;
assign micromatrizz[13][572] = 9'b111111111;
assign micromatrizz[13][573] = 9'b111111111;
assign micromatrizz[13][574] = 9'b111111111;
assign micromatrizz[13][575] = 9'b111111111;
assign micromatrizz[13][576] = 9'b111111111;
assign micromatrizz[13][577] = 9'b111111111;
assign micromatrizz[13][578] = 9'b111111111;
assign micromatrizz[13][579] = 9'b111111111;
assign micromatrizz[13][580] = 9'b111111111;
assign micromatrizz[13][581] = 9'b111111111;
assign micromatrizz[13][582] = 9'b111111111;
assign micromatrizz[13][583] = 9'b111111111;
assign micromatrizz[13][584] = 9'b111111111;
assign micromatrizz[13][585] = 9'b111111111;
assign micromatrizz[13][586] = 9'b111111111;
assign micromatrizz[13][587] = 9'b111111111;
assign micromatrizz[13][588] = 9'b111111111;
assign micromatrizz[13][589] = 9'b111111111;
assign micromatrizz[13][590] = 9'b111111111;
assign micromatrizz[13][591] = 9'b111111111;
assign micromatrizz[13][592] = 9'b111111111;
assign micromatrizz[13][593] = 9'b111111111;
assign micromatrizz[13][594] = 9'b111111111;
assign micromatrizz[13][595] = 9'b111111111;
assign micromatrizz[13][596] = 9'b111111111;
assign micromatrizz[13][597] = 9'b111111111;
assign micromatrizz[13][598] = 9'b111111111;
assign micromatrizz[13][599] = 9'b111111111;
assign micromatrizz[13][600] = 9'b111111111;
assign micromatrizz[13][601] = 9'b111111111;
assign micromatrizz[13][602] = 9'b111111111;
assign micromatrizz[13][603] = 9'b111111111;
assign micromatrizz[13][604] = 9'b111111111;
assign micromatrizz[13][605] = 9'b111111111;
assign micromatrizz[13][606] = 9'b111111111;
assign micromatrizz[13][607] = 9'b111111111;
assign micromatrizz[13][608] = 9'b111111111;
assign micromatrizz[13][609] = 9'b111111111;
assign micromatrizz[13][610] = 9'b111111111;
assign micromatrizz[13][611] = 9'b111111111;
assign micromatrizz[13][612] = 9'b111111111;
assign micromatrizz[13][613] = 9'b111111111;
assign micromatrizz[13][614] = 9'b111111111;
assign micromatrizz[13][615] = 9'b111111111;
assign micromatrizz[13][616] = 9'b111111111;
assign micromatrizz[13][617] = 9'b111111111;
assign micromatrizz[13][618] = 9'b111111111;
assign micromatrizz[13][619] = 9'b111111111;
assign micromatrizz[13][620] = 9'b111111111;
assign micromatrizz[13][621] = 9'b111111111;
assign micromatrizz[13][622] = 9'b111111111;
assign micromatrizz[13][623] = 9'b111111111;
assign micromatrizz[13][624] = 9'b111111111;
assign micromatrizz[13][625] = 9'b111111111;
assign micromatrizz[13][626] = 9'b111111111;
assign micromatrizz[13][627] = 9'b111111111;
assign micromatrizz[13][628] = 9'b111111111;
assign micromatrizz[13][629] = 9'b111111111;
assign micromatrizz[13][630] = 9'b111111111;
assign micromatrizz[13][631] = 9'b111111111;
assign micromatrizz[13][632] = 9'b111111111;
assign micromatrizz[13][633] = 9'b111111111;
assign micromatrizz[13][634] = 9'b111111111;
assign micromatrizz[13][635] = 9'b111111111;
assign micromatrizz[13][636] = 9'b111111111;
assign micromatrizz[13][637] = 9'b111111111;
assign micromatrizz[13][638] = 9'b111111111;
assign micromatrizz[13][639] = 9'b111111111;
assign micromatrizz[14][0] = 9'b111111111;
assign micromatrizz[14][1] = 9'b111111111;
assign micromatrizz[14][2] = 9'b111111111;
assign micromatrizz[14][3] = 9'b111111111;
assign micromatrizz[14][4] = 9'b111111111;
assign micromatrizz[14][5] = 9'b111111111;
assign micromatrizz[14][6] = 9'b111111111;
assign micromatrizz[14][7] = 9'b111111111;
assign micromatrizz[14][8] = 9'b111111111;
assign micromatrizz[14][9] = 9'b111111111;
assign micromatrizz[14][10] = 9'b111111111;
assign micromatrizz[14][11] = 9'b111111111;
assign micromatrizz[14][12] = 9'b111111111;
assign micromatrizz[14][13] = 9'b111111111;
assign micromatrizz[14][14] = 9'b111111111;
assign micromatrizz[14][15] = 9'b111111111;
assign micromatrizz[14][16] = 9'b111111111;
assign micromatrizz[14][17] = 9'b111111111;
assign micromatrizz[14][18] = 9'b111111111;
assign micromatrizz[14][19] = 9'b111111111;
assign micromatrizz[14][20] = 9'b111111111;
assign micromatrizz[14][21] = 9'b111111111;
assign micromatrizz[14][22] = 9'b111111111;
assign micromatrizz[14][23] = 9'b111111111;
assign micromatrizz[14][24] = 9'b111111111;
assign micromatrizz[14][25] = 9'b111111111;
assign micromatrizz[14][26] = 9'b111111111;
assign micromatrizz[14][27] = 9'b111111111;
assign micromatrizz[14][28] = 9'b111111111;
assign micromatrizz[14][29] = 9'b111111111;
assign micromatrizz[14][30] = 9'b111111111;
assign micromatrizz[14][31] = 9'b111111111;
assign micromatrizz[14][32] = 9'b111111111;
assign micromatrizz[14][33] = 9'b111111111;
assign micromatrizz[14][34] = 9'b111111111;
assign micromatrizz[14][35] = 9'b111111111;
assign micromatrizz[14][36] = 9'b111111111;
assign micromatrizz[14][37] = 9'b111111111;
assign micromatrizz[14][38] = 9'b111111111;
assign micromatrizz[14][39] = 9'b111111111;
assign micromatrizz[14][40] = 9'b111111111;
assign micromatrizz[14][41] = 9'b111111111;
assign micromatrizz[14][42] = 9'b111111111;
assign micromatrizz[14][43] = 9'b111111111;
assign micromatrizz[14][44] = 9'b111111111;
assign micromatrizz[14][45] = 9'b111111111;
assign micromatrizz[14][46] = 9'b111111111;
assign micromatrizz[14][47] = 9'b111111111;
assign micromatrizz[14][48] = 9'b111111111;
assign micromatrizz[14][49] = 9'b111111111;
assign micromatrizz[14][50] = 9'b111111111;
assign micromatrizz[14][51] = 9'b111111111;
assign micromatrizz[14][52] = 9'b111111111;
assign micromatrizz[14][53] = 9'b111111111;
assign micromatrizz[14][54] = 9'b111111111;
assign micromatrizz[14][55] = 9'b111111111;
assign micromatrizz[14][56] = 9'b111111111;
assign micromatrizz[14][57] = 9'b111111111;
assign micromatrizz[14][58] = 9'b111111111;
assign micromatrizz[14][59] = 9'b111111111;
assign micromatrizz[14][60] = 9'b111111111;
assign micromatrizz[14][61] = 9'b111111111;
assign micromatrizz[14][62] = 9'b111111111;
assign micromatrizz[14][63] = 9'b111111111;
assign micromatrizz[14][64] = 9'b111111111;
assign micromatrizz[14][65] = 9'b111111111;
assign micromatrizz[14][66] = 9'b111111111;
assign micromatrizz[14][67] = 9'b111111111;
assign micromatrizz[14][68] = 9'b111111111;
assign micromatrizz[14][69] = 9'b111111111;
assign micromatrizz[14][70] = 9'b111111111;
assign micromatrizz[14][71] = 9'b111111111;
assign micromatrizz[14][72] = 9'b111111111;
assign micromatrizz[14][73] = 9'b111111111;
assign micromatrizz[14][74] = 9'b111111111;
assign micromatrizz[14][75] = 9'b111111111;
assign micromatrizz[14][76] = 9'b111111111;
assign micromatrizz[14][77] = 9'b111111111;
assign micromatrizz[14][78] = 9'b111111111;
assign micromatrizz[14][79] = 9'b111111111;
assign micromatrizz[14][80] = 9'b111111111;
assign micromatrizz[14][81] = 9'b111111111;
assign micromatrizz[14][82] = 9'b111111111;
assign micromatrizz[14][83] = 9'b111111111;
assign micromatrizz[14][84] = 9'b111111111;
assign micromatrizz[14][85] = 9'b111111111;
assign micromatrizz[14][86] = 9'b111111111;
assign micromatrizz[14][87] = 9'b111111111;
assign micromatrizz[14][88] = 9'b111111111;
assign micromatrizz[14][89] = 9'b111111111;
assign micromatrizz[14][90] = 9'b111111111;
assign micromatrizz[14][91] = 9'b111111111;
assign micromatrizz[14][92] = 9'b111111111;
assign micromatrizz[14][93] = 9'b111111111;
assign micromatrizz[14][94] = 9'b111111111;
assign micromatrizz[14][95] = 9'b111111111;
assign micromatrizz[14][96] = 9'b111111111;
assign micromatrizz[14][97] = 9'b111111111;
assign micromatrizz[14][98] = 9'b111111111;
assign micromatrizz[14][99] = 9'b111111111;
assign micromatrizz[14][100] = 9'b111111111;
assign micromatrizz[14][101] = 9'b111111111;
assign micromatrizz[14][102] = 9'b111111111;
assign micromatrizz[14][103] = 9'b111111111;
assign micromatrizz[14][104] = 9'b111111111;
assign micromatrizz[14][105] = 9'b111111111;
assign micromatrizz[14][106] = 9'b111111111;
assign micromatrizz[14][107] = 9'b111111111;
assign micromatrizz[14][108] = 9'b111111111;
assign micromatrizz[14][109] = 9'b111111111;
assign micromatrizz[14][110] = 9'b111111111;
assign micromatrizz[14][111] = 9'b111111111;
assign micromatrizz[14][112] = 9'b111111111;
assign micromatrizz[14][113] = 9'b111111111;
assign micromatrizz[14][114] = 9'b111111111;
assign micromatrizz[14][115] = 9'b111111111;
assign micromatrizz[14][116] = 9'b111111111;
assign micromatrizz[14][117] = 9'b111111111;
assign micromatrizz[14][118] = 9'b111111111;
assign micromatrizz[14][119] = 9'b111111111;
assign micromatrizz[14][120] = 9'b111111111;
assign micromatrizz[14][121] = 9'b111111111;
assign micromatrizz[14][122] = 9'b111111111;
assign micromatrizz[14][123] = 9'b111111111;
assign micromatrizz[14][124] = 9'b111111111;
assign micromatrizz[14][125] = 9'b111111111;
assign micromatrizz[14][126] = 9'b111111111;
assign micromatrizz[14][127] = 9'b111111111;
assign micromatrizz[14][128] = 9'b111111111;
assign micromatrizz[14][129] = 9'b111111111;
assign micromatrizz[14][130] = 9'b111111111;
assign micromatrizz[14][131] = 9'b111111111;
assign micromatrizz[14][132] = 9'b111111111;
assign micromatrizz[14][133] = 9'b111111111;
assign micromatrizz[14][134] = 9'b111111111;
assign micromatrizz[14][135] = 9'b111111111;
assign micromatrizz[14][136] = 9'b111111111;
assign micromatrizz[14][137] = 9'b111111111;
assign micromatrizz[14][138] = 9'b111111111;
assign micromatrizz[14][139] = 9'b111111111;
assign micromatrizz[14][140] = 9'b111111111;
assign micromatrizz[14][141] = 9'b111111111;
assign micromatrizz[14][142] = 9'b111111111;
assign micromatrizz[14][143] = 9'b111111111;
assign micromatrizz[14][144] = 9'b111111111;
assign micromatrizz[14][145] = 9'b111111111;
assign micromatrizz[14][146] = 9'b111111111;
assign micromatrizz[14][147] = 9'b111111111;
assign micromatrizz[14][148] = 9'b111111111;
assign micromatrizz[14][149] = 9'b111111111;
assign micromatrizz[14][150] = 9'b111111111;
assign micromatrizz[14][151] = 9'b111111111;
assign micromatrizz[14][152] = 9'b111111111;
assign micromatrizz[14][153] = 9'b111111111;
assign micromatrizz[14][154] = 9'b111111111;
assign micromatrizz[14][155] = 9'b111111111;
assign micromatrizz[14][156] = 9'b111111111;
assign micromatrizz[14][157] = 9'b111111111;
assign micromatrizz[14][158] = 9'b111111111;
assign micromatrizz[14][159] = 9'b111111111;
assign micromatrizz[14][160] = 9'b111111111;
assign micromatrizz[14][161] = 9'b111111111;
assign micromatrizz[14][162] = 9'b111111111;
assign micromatrizz[14][163] = 9'b111111111;
assign micromatrizz[14][164] = 9'b111111111;
assign micromatrizz[14][165] = 9'b111111111;
assign micromatrizz[14][166] = 9'b111111111;
assign micromatrizz[14][167] = 9'b111111111;
assign micromatrizz[14][168] = 9'b111111111;
assign micromatrizz[14][169] = 9'b111111111;
assign micromatrizz[14][170] = 9'b111111111;
assign micromatrizz[14][171] = 9'b111111111;
assign micromatrizz[14][172] = 9'b111111111;
assign micromatrizz[14][173] = 9'b111111111;
assign micromatrizz[14][174] = 9'b111111111;
assign micromatrizz[14][175] = 9'b111111111;
assign micromatrizz[14][176] = 9'b111111111;
assign micromatrizz[14][177] = 9'b111111111;
assign micromatrizz[14][178] = 9'b111111111;
assign micromatrizz[14][179] = 9'b111111111;
assign micromatrizz[14][180] = 9'b111111111;
assign micromatrizz[14][181] = 9'b111111111;
assign micromatrizz[14][182] = 9'b111111111;
assign micromatrizz[14][183] = 9'b111111111;
assign micromatrizz[14][184] = 9'b111111111;
assign micromatrizz[14][185] = 9'b111111111;
assign micromatrizz[14][186] = 9'b111111111;
assign micromatrizz[14][187] = 9'b111111111;
assign micromatrizz[14][188] = 9'b111111111;
assign micromatrizz[14][189] = 9'b111111111;
assign micromatrizz[14][190] = 9'b111111111;
assign micromatrizz[14][191] = 9'b111111111;
assign micromatrizz[14][192] = 9'b111111111;
assign micromatrizz[14][193] = 9'b111111111;
assign micromatrizz[14][194] = 9'b111111111;
assign micromatrizz[14][195] = 9'b111111111;
assign micromatrizz[14][196] = 9'b111111111;
assign micromatrizz[14][197] = 9'b111111111;
assign micromatrizz[14][198] = 9'b111111111;
assign micromatrizz[14][199] = 9'b111111111;
assign micromatrizz[14][200] = 9'b111111111;
assign micromatrizz[14][201] = 9'b111111111;
assign micromatrizz[14][202] = 9'b111111111;
assign micromatrizz[14][203] = 9'b111111111;
assign micromatrizz[14][204] = 9'b111111111;
assign micromatrizz[14][205] = 9'b111111111;
assign micromatrizz[14][206] = 9'b111111111;
assign micromatrizz[14][207] = 9'b111111111;
assign micromatrizz[14][208] = 9'b111111111;
assign micromatrizz[14][209] = 9'b111111111;
assign micromatrizz[14][210] = 9'b111111111;
assign micromatrizz[14][211] = 9'b111111111;
assign micromatrizz[14][212] = 9'b111111111;
assign micromatrizz[14][213] = 9'b111111111;
assign micromatrizz[14][214] = 9'b111111111;
assign micromatrizz[14][215] = 9'b111111111;
assign micromatrizz[14][216] = 9'b111111111;
assign micromatrizz[14][217] = 9'b111111111;
assign micromatrizz[14][218] = 9'b111111111;
assign micromatrizz[14][219] = 9'b111111111;
assign micromatrizz[14][220] = 9'b111111111;
assign micromatrizz[14][221] = 9'b111111111;
assign micromatrizz[14][222] = 9'b111111111;
assign micromatrizz[14][223] = 9'b111111111;
assign micromatrizz[14][224] = 9'b111111111;
assign micromatrizz[14][225] = 9'b111111111;
assign micromatrizz[14][226] = 9'b111111111;
assign micromatrizz[14][227] = 9'b111111111;
assign micromatrizz[14][228] = 9'b111111111;
assign micromatrizz[14][229] = 9'b111111111;
assign micromatrizz[14][230] = 9'b111111111;
assign micromatrizz[14][231] = 9'b111111111;
assign micromatrizz[14][232] = 9'b111111111;
assign micromatrizz[14][233] = 9'b111111111;
assign micromatrizz[14][234] = 9'b111111111;
assign micromatrizz[14][235] = 9'b111111111;
assign micromatrizz[14][236] = 9'b111111111;
assign micromatrizz[14][237] = 9'b111111111;
assign micromatrizz[14][238] = 9'b111111111;
assign micromatrizz[14][239] = 9'b111111111;
assign micromatrizz[14][240] = 9'b111111111;
assign micromatrizz[14][241] = 9'b111111111;
assign micromatrizz[14][242] = 9'b111111111;
assign micromatrizz[14][243] = 9'b111111111;
assign micromatrizz[14][244] = 9'b111111111;
assign micromatrizz[14][245] = 9'b111111111;
assign micromatrizz[14][246] = 9'b111111111;
assign micromatrizz[14][247] = 9'b111111111;
assign micromatrizz[14][248] = 9'b111111111;
assign micromatrizz[14][249] = 9'b111111111;
assign micromatrizz[14][250] = 9'b111111111;
assign micromatrizz[14][251] = 9'b111111111;
assign micromatrizz[14][252] = 9'b111111111;
assign micromatrizz[14][253] = 9'b111111111;
assign micromatrizz[14][254] = 9'b111111111;
assign micromatrizz[14][255] = 9'b111111111;
assign micromatrizz[14][256] = 9'b111111111;
assign micromatrizz[14][257] = 9'b111111111;
assign micromatrizz[14][258] = 9'b111111111;
assign micromatrizz[14][259] = 9'b111111111;
assign micromatrizz[14][260] = 9'b111111111;
assign micromatrizz[14][261] = 9'b111111111;
assign micromatrizz[14][262] = 9'b111111111;
assign micromatrizz[14][263] = 9'b111111111;
assign micromatrizz[14][264] = 9'b111111111;
assign micromatrizz[14][265] = 9'b111111111;
assign micromatrizz[14][266] = 9'b111111111;
assign micromatrizz[14][267] = 9'b111111111;
assign micromatrizz[14][268] = 9'b111111111;
assign micromatrizz[14][269] = 9'b111111111;
assign micromatrizz[14][270] = 9'b111111111;
assign micromatrizz[14][271] = 9'b111111111;
assign micromatrizz[14][272] = 9'b111111111;
assign micromatrizz[14][273] = 9'b111111111;
assign micromatrizz[14][274] = 9'b111111111;
assign micromatrizz[14][275] = 9'b111111111;
assign micromatrizz[14][276] = 9'b111111111;
assign micromatrizz[14][277] = 9'b111111111;
assign micromatrizz[14][278] = 9'b111111111;
assign micromatrizz[14][279] = 9'b111111111;
assign micromatrizz[14][280] = 9'b111111111;
assign micromatrizz[14][281] = 9'b111111111;
assign micromatrizz[14][282] = 9'b111111111;
assign micromatrizz[14][283] = 9'b111111111;
assign micromatrizz[14][284] = 9'b111111111;
assign micromatrizz[14][285] = 9'b111111111;
assign micromatrizz[14][286] = 9'b111111111;
assign micromatrizz[14][287] = 9'b111111111;
assign micromatrizz[14][288] = 9'b111111111;
assign micromatrizz[14][289] = 9'b111111111;
assign micromatrizz[14][290] = 9'b111111111;
assign micromatrizz[14][291] = 9'b111111111;
assign micromatrizz[14][292] = 9'b111111111;
assign micromatrizz[14][293] = 9'b111111111;
assign micromatrizz[14][294] = 9'b111111111;
assign micromatrizz[14][295] = 9'b111111111;
assign micromatrizz[14][296] = 9'b111111111;
assign micromatrizz[14][297] = 9'b111111111;
assign micromatrizz[14][298] = 9'b111111111;
assign micromatrizz[14][299] = 9'b111111111;
assign micromatrizz[14][300] = 9'b111111111;
assign micromatrizz[14][301] = 9'b111111111;
assign micromatrizz[14][302] = 9'b111111111;
assign micromatrizz[14][303] = 9'b111111111;
assign micromatrizz[14][304] = 9'b111111111;
assign micromatrizz[14][305] = 9'b111111111;
assign micromatrizz[14][306] = 9'b111111111;
assign micromatrizz[14][307] = 9'b111111111;
assign micromatrizz[14][308] = 9'b111111111;
assign micromatrizz[14][309] = 9'b111111111;
assign micromatrizz[14][310] = 9'b111111111;
assign micromatrizz[14][311] = 9'b111111111;
assign micromatrizz[14][312] = 9'b111111111;
assign micromatrizz[14][313] = 9'b111111111;
assign micromatrizz[14][314] = 9'b111111111;
assign micromatrizz[14][315] = 9'b111111111;
assign micromatrizz[14][316] = 9'b111111111;
assign micromatrizz[14][317] = 9'b111111111;
assign micromatrizz[14][318] = 9'b111111111;
assign micromatrizz[14][319] = 9'b111111111;
assign micromatrizz[14][320] = 9'b111111111;
assign micromatrizz[14][321] = 9'b111111111;
assign micromatrizz[14][322] = 9'b111111111;
assign micromatrizz[14][323] = 9'b111111111;
assign micromatrizz[14][324] = 9'b111111111;
assign micromatrizz[14][325] = 9'b111111111;
assign micromatrizz[14][326] = 9'b111111111;
assign micromatrizz[14][327] = 9'b111111111;
assign micromatrizz[14][328] = 9'b111111111;
assign micromatrizz[14][329] = 9'b111111111;
assign micromatrizz[14][330] = 9'b111111111;
assign micromatrizz[14][331] = 9'b111111111;
assign micromatrizz[14][332] = 9'b111111111;
assign micromatrizz[14][333] = 9'b111111111;
assign micromatrizz[14][334] = 9'b111111111;
assign micromatrizz[14][335] = 9'b111111111;
assign micromatrizz[14][336] = 9'b111111111;
assign micromatrizz[14][337] = 9'b111111111;
assign micromatrizz[14][338] = 9'b111111111;
assign micromatrizz[14][339] = 9'b111111111;
assign micromatrizz[14][340] = 9'b111111111;
assign micromatrizz[14][341] = 9'b111111111;
assign micromatrizz[14][342] = 9'b111111111;
assign micromatrizz[14][343] = 9'b111111111;
assign micromatrizz[14][344] = 9'b111111111;
assign micromatrizz[14][345] = 9'b111111111;
assign micromatrizz[14][346] = 9'b111111111;
assign micromatrizz[14][347] = 9'b111111111;
assign micromatrizz[14][348] = 9'b111111111;
assign micromatrizz[14][349] = 9'b111111111;
assign micromatrizz[14][350] = 9'b111111111;
assign micromatrizz[14][351] = 9'b111111111;
assign micromatrizz[14][352] = 9'b111111111;
assign micromatrizz[14][353] = 9'b111111111;
assign micromatrizz[14][354] = 9'b111111111;
assign micromatrizz[14][355] = 9'b111111111;
assign micromatrizz[14][356] = 9'b111111111;
assign micromatrizz[14][357] = 9'b111111111;
assign micromatrizz[14][358] = 9'b111111111;
assign micromatrizz[14][359] = 9'b111111111;
assign micromatrizz[14][360] = 9'b111111111;
assign micromatrizz[14][361] = 9'b111111111;
assign micromatrizz[14][362] = 9'b111111111;
assign micromatrizz[14][363] = 9'b111111111;
assign micromatrizz[14][364] = 9'b111111111;
assign micromatrizz[14][365] = 9'b111111111;
assign micromatrizz[14][366] = 9'b111111111;
assign micromatrizz[14][367] = 9'b111111111;
assign micromatrizz[14][368] = 9'b111111111;
assign micromatrizz[14][369] = 9'b111111111;
assign micromatrizz[14][370] = 9'b111111111;
assign micromatrizz[14][371] = 9'b111111111;
assign micromatrizz[14][372] = 9'b111111111;
assign micromatrizz[14][373] = 9'b111111111;
assign micromatrizz[14][374] = 9'b111111111;
assign micromatrizz[14][375] = 9'b111111111;
assign micromatrizz[14][376] = 9'b111111111;
assign micromatrizz[14][377] = 9'b111111111;
assign micromatrizz[14][378] = 9'b111111111;
assign micromatrizz[14][379] = 9'b111111111;
assign micromatrizz[14][380] = 9'b111111111;
assign micromatrizz[14][381] = 9'b111111111;
assign micromatrizz[14][382] = 9'b111111111;
assign micromatrizz[14][383] = 9'b111111111;
assign micromatrizz[14][384] = 9'b111111111;
assign micromatrizz[14][385] = 9'b111111111;
assign micromatrizz[14][386] = 9'b111111111;
assign micromatrizz[14][387] = 9'b111111111;
assign micromatrizz[14][388] = 9'b111111111;
assign micromatrizz[14][389] = 9'b111111111;
assign micromatrizz[14][390] = 9'b111111111;
assign micromatrizz[14][391] = 9'b111111111;
assign micromatrizz[14][392] = 9'b111111111;
assign micromatrizz[14][393] = 9'b111111111;
assign micromatrizz[14][394] = 9'b111111111;
assign micromatrizz[14][395] = 9'b111111111;
assign micromatrizz[14][396] = 9'b111111111;
assign micromatrizz[14][397] = 9'b111111111;
assign micromatrizz[14][398] = 9'b111111111;
assign micromatrizz[14][399] = 9'b111111111;
assign micromatrizz[14][400] = 9'b111111111;
assign micromatrizz[14][401] = 9'b111111111;
assign micromatrizz[14][402] = 9'b111111111;
assign micromatrizz[14][403] = 9'b111111111;
assign micromatrizz[14][404] = 9'b111111111;
assign micromatrizz[14][405] = 9'b111111111;
assign micromatrizz[14][406] = 9'b111111111;
assign micromatrizz[14][407] = 9'b111111111;
assign micromatrizz[14][408] = 9'b111111111;
assign micromatrizz[14][409] = 9'b111111111;
assign micromatrizz[14][410] = 9'b111111111;
assign micromatrizz[14][411] = 9'b111111111;
assign micromatrizz[14][412] = 9'b111111111;
assign micromatrizz[14][413] = 9'b111111111;
assign micromatrizz[14][414] = 9'b111111111;
assign micromatrizz[14][415] = 9'b111111111;
assign micromatrizz[14][416] = 9'b111111111;
assign micromatrizz[14][417] = 9'b111111111;
assign micromatrizz[14][418] = 9'b111111111;
assign micromatrizz[14][419] = 9'b111111111;
assign micromatrizz[14][420] = 9'b111111111;
assign micromatrizz[14][421] = 9'b111111111;
assign micromatrizz[14][422] = 9'b111111111;
assign micromatrizz[14][423] = 9'b111111111;
assign micromatrizz[14][424] = 9'b111111111;
assign micromatrizz[14][425] = 9'b111111111;
assign micromatrizz[14][426] = 9'b111111111;
assign micromatrizz[14][427] = 9'b111111111;
assign micromatrizz[14][428] = 9'b111111111;
assign micromatrizz[14][429] = 9'b111111111;
assign micromatrizz[14][430] = 9'b111111111;
assign micromatrizz[14][431] = 9'b111111111;
assign micromatrizz[14][432] = 9'b111111111;
assign micromatrizz[14][433] = 9'b111111111;
assign micromatrizz[14][434] = 9'b111111111;
assign micromatrizz[14][435] = 9'b111111111;
assign micromatrizz[14][436] = 9'b111111111;
assign micromatrizz[14][437] = 9'b111111111;
assign micromatrizz[14][438] = 9'b111111111;
assign micromatrizz[14][439] = 9'b111111111;
assign micromatrizz[14][440] = 9'b111111111;
assign micromatrizz[14][441] = 9'b111111111;
assign micromatrizz[14][442] = 9'b111111111;
assign micromatrizz[14][443] = 9'b111111111;
assign micromatrizz[14][444] = 9'b111111111;
assign micromatrizz[14][445] = 9'b111111111;
assign micromatrizz[14][446] = 9'b111111111;
assign micromatrizz[14][447] = 9'b111111111;
assign micromatrizz[14][448] = 9'b111111111;
assign micromatrizz[14][449] = 9'b111111111;
assign micromatrizz[14][450] = 9'b111111111;
assign micromatrizz[14][451] = 9'b111111111;
assign micromatrizz[14][452] = 9'b111111111;
assign micromatrizz[14][453] = 9'b111111111;
assign micromatrizz[14][454] = 9'b111111111;
assign micromatrizz[14][455] = 9'b111111111;
assign micromatrizz[14][456] = 9'b111111111;
assign micromatrizz[14][457] = 9'b111111111;
assign micromatrizz[14][458] = 9'b111111111;
assign micromatrizz[14][459] = 9'b111111111;
assign micromatrizz[14][460] = 9'b111111111;
assign micromatrizz[14][461] = 9'b111111111;
assign micromatrizz[14][462] = 9'b111111111;
assign micromatrizz[14][463] = 9'b111111111;
assign micromatrizz[14][464] = 9'b111111111;
assign micromatrizz[14][465] = 9'b111111111;
assign micromatrizz[14][466] = 9'b111111111;
assign micromatrizz[14][467] = 9'b111111111;
assign micromatrizz[14][468] = 9'b111111111;
assign micromatrizz[14][469] = 9'b111111111;
assign micromatrizz[14][470] = 9'b111111111;
assign micromatrizz[14][471] = 9'b111111111;
assign micromatrizz[14][472] = 9'b111111111;
assign micromatrizz[14][473] = 9'b111111111;
assign micromatrizz[14][474] = 9'b111111111;
assign micromatrizz[14][475] = 9'b111111111;
assign micromatrizz[14][476] = 9'b111111111;
assign micromatrizz[14][477] = 9'b111111111;
assign micromatrizz[14][478] = 9'b111111111;
assign micromatrizz[14][479] = 9'b111111111;
assign micromatrizz[14][480] = 9'b111111111;
assign micromatrizz[14][481] = 9'b111111111;
assign micromatrizz[14][482] = 9'b111111111;
assign micromatrizz[14][483] = 9'b111111111;
assign micromatrizz[14][484] = 9'b111111111;
assign micromatrizz[14][485] = 9'b111111111;
assign micromatrizz[14][486] = 9'b111111111;
assign micromatrizz[14][487] = 9'b111111111;
assign micromatrizz[14][488] = 9'b111111111;
assign micromatrizz[14][489] = 9'b111111111;
assign micromatrizz[14][490] = 9'b111111111;
assign micromatrizz[14][491] = 9'b111111111;
assign micromatrizz[14][492] = 9'b111111111;
assign micromatrizz[14][493] = 9'b111111111;
assign micromatrizz[14][494] = 9'b111111111;
assign micromatrizz[14][495] = 9'b111111111;
assign micromatrizz[14][496] = 9'b111111111;
assign micromatrizz[14][497] = 9'b111111111;
assign micromatrizz[14][498] = 9'b111111111;
assign micromatrizz[14][499] = 9'b111111111;
assign micromatrizz[14][500] = 9'b111111111;
assign micromatrizz[14][501] = 9'b111111111;
assign micromatrizz[14][502] = 9'b111111111;
assign micromatrizz[14][503] = 9'b111111111;
assign micromatrizz[14][504] = 9'b111111111;
assign micromatrizz[14][505] = 9'b111111111;
assign micromatrizz[14][506] = 9'b111111111;
assign micromatrizz[14][507] = 9'b111111111;
assign micromatrizz[14][508] = 9'b111111111;
assign micromatrizz[14][509] = 9'b111111111;
assign micromatrizz[14][510] = 9'b111111111;
assign micromatrizz[14][511] = 9'b111111111;
assign micromatrizz[14][512] = 9'b111111111;
assign micromatrizz[14][513] = 9'b111111111;
assign micromatrizz[14][514] = 9'b111111111;
assign micromatrizz[14][515] = 9'b111111111;
assign micromatrizz[14][516] = 9'b111111111;
assign micromatrizz[14][517] = 9'b111111111;
assign micromatrizz[14][518] = 9'b111111111;
assign micromatrizz[14][519] = 9'b111111111;
assign micromatrizz[14][520] = 9'b111111111;
assign micromatrizz[14][521] = 9'b111111111;
assign micromatrizz[14][522] = 9'b111111111;
assign micromatrizz[14][523] = 9'b111111111;
assign micromatrizz[14][524] = 9'b111111111;
assign micromatrizz[14][525] = 9'b111111111;
assign micromatrizz[14][526] = 9'b111111111;
assign micromatrizz[14][527] = 9'b111111111;
assign micromatrizz[14][528] = 9'b111111111;
assign micromatrizz[14][529] = 9'b111111111;
assign micromatrizz[14][530] = 9'b111111111;
assign micromatrizz[14][531] = 9'b111111111;
assign micromatrizz[14][532] = 9'b111111111;
assign micromatrizz[14][533] = 9'b111111111;
assign micromatrizz[14][534] = 9'b111111111;
assign micromatrizz[14][535] = 9'b111111111;
assign micromatrizz[14][536] = 9'b111111111;
assign micromatrizz[14][537] = 9'b111111111;
assign micromatrizz[14][538] = 9'b111111111;
assign micromatrizz[14][539] = 9'b111111111;
assign micromatrizz[14][540] = 9'b111111111;
assign micromatrizz[14][541] = 9'b111111111;
assign micromatrizz[14][542] = 9'b111111111;
assign micromatrizz[14][543] = 9'b111111111;
assign micromatrizz[14][544] = 9'b111111111;
assign micromatrizz[14][545] = 9'b111111111;
assign micromatrizz[14][546] = 9'b111111111;
assign micromatrizz[14][547] = 9'b111111111;
assign micromatrizz[14][548] = 9'b111111111;
assign micromatrizz[14][549] = 9'b111111111;
assign micromatrizz[14][550] = 9'b111111111;
assign micromatrizz[14][551] = 9'b111111111;
assign micromatrizz[14][552] = 9'b111111111;
assign micromatrizz[14][553] = 9'b111111111;
assign micromatrizz[14][554] = 9'b111111111;
assign micromatrizz[14][555] = 9'b111111111;
assign micromatrizz[14][556] = 9'b111111111;
assign micromatrizz[14][557] = 9'b111111111;
assign micromatrizz[14][558] = 9'b111111111;
assign micromatrizz[14][559] = 9'b111111111;
assign micromatrizz[14][560] = 9'b111111111;
assign micromatrizz[14][561] = 9'b111111111;
assign micromatrizz[14][562] = 9'b111111111;
assign micromatrizz[14][563] = 9'b111111111;
assign micromatrizz[14][564] = 9'b111111111;
assign micromatrizz[14][565] = 9'b111111111;
assign micromatrizz[14][566] = 9'b111111111;
assign micromatrizz[14][567] = 9'b111111111;
assign micromatrizz[14][568] = 9'b111111111;
assign micromatrizz[14][569] = 9'b111111111;
assign micromatrizz[14][570] = 9'b111111111;
assign micromatrizz[14][571] = 9'b111111111;
assign micromatrizz[14][572] = 9'b111111111;
assign micromatrizz[14][573] = 9'b111111111;
assign micromatrizz[14][574] = 9'b111111111;
assign micromatrizz[14][575] = 9'b111111111;
assign micromatrizz[14][576] = 9'b111111111;
assign micromatrizz[14][577] = 9'b111111111;
assign micromatrizz[14][578] = 9'b111111111;
assign micromatrizz[14][579] = 9'b111111111;
assign micromatrizz[14][580] = 9'b111111111;
assign micromatrizz[14][581] = 9'b111111111;
assign micromatrizz[14][582] = 9'b111111111;
assign micromatrizz[14][583] = 9'b111111111;
assign micromatrizz[14][584] = 9'b111111111;
assign micromatrizz[14][585] = 9'b111111111;
assign micromatrizz[14][586] = 9'b111111111;
assign micromatrizz[14][587] = 9'b111111111;
assign micromatrizz[14][588] = 9'b111111111;
assign micromatrizz[14][589] = 9'b111111111;
assign micromatrizz[14][590] = 9'b111111111;
assign micromatrizz[14][591] = 9'b111111111;
assign micromatrizz[14][592] = 9'b111111111;
assign micromatrizz[14][593] = 9'b111111111;
assign micromatrizz[14][594] = 9'b111111111;
assign micromatrizz[14][595] = 9'b111111111;
assign micromatrizz[14][596] = 9'b111111111;
assign micromatrizz[14][597] = 9'b111111111;
assign micromatrizz[14][598] = 9'b111111111;
assign micromatrizz[14][599] = 9'b111111111;
assign micromatrizz[14][600] = 9'b111111111;
assign micromatrizz[14][601] = 9'b111111111;
assign micromatrizz[14][602] = 9'b111111111;
assign micromatrizz[14][603] = 9'b111111111;
assign micromatrizz[14][604] = 9'b111111111;
assign micromatrizz[14][605] = 9'b111111111;
assign micromatrizz[14][606] = 9'b111111111;
assign micromatrizz[14][607] = 9'b111111111;
assign micromatrizz[14][608] = 9'b111111111;
assign micromatrizz[14][609] = 9'b111111111;
assign micromatrizz[14][610] = 9'b111111111;
assign micromatrizz[14][611] = 9'b111111111;
assign micromatrizz[14][612] = 9'b111111111;
assign micromatrizz[14][613] = 9'b111111111;
assign micromatrizz[14][614] = 9'b111111111;
assign micromatrizz[14][615] = 9'b111111111;
assign micromatrizz[14][616] = 9'b111111111;
assign micromatrizz[14][617] = 9'b111111111;
assign micromatrizz[14][618] = 9'b111111111;
assign micromatrizz[14][619] = 9'b111111111;
assign micromatrizz[14][620] = 9'b111111111;
assign micromatrizz[14][621] = 9'b111111111;
assign micromatrizz[14][622] = 9'b111111111;
assign micromatrizz[14][623] = 9'b111111111;
assign micromatrizz[14][624] = 9'b111111111;
assign micromatrizz[14][625] = 9'b111111111;
assign micromatrizz[14][626] = 9'b111111111;
assign micromatrizz[14][627] = 9'b111111111;
assign micromatrizz[14][628] = 9'b111111111;
assign micromatrizz[14][629] = 9'b111111111;
assign micromatrizz[14][630] = 9'b111111111;
assign micromatrizz[14][631] = 9'b111111111;
assign micromatrizz[14][632] = 9'b111111111;
assign micromatrizz[14][633] = 9'b111111111;
assign micromatrizz[14][634] = 9'b111111111;
assign micromatrizz[14][635] = 9'b111111111;
assign micromatrizz[14][636] = 9'b111111111;
assign micromatrizz[14][637] = 9'b111111111;
assign micromatrizz[14][638] = 9'b111111111;
assign micromatrizz[14][639] = 9'b111111111;
assign micromatrizz[15][0] = 9'b111111111;
assign micromatrizz[15][1] = 9'b111111111;
assign micromatrizz[15][2] = 9'b111111111;
assign micromatrizz[15][3] = 9'b111111111;
assign micromatrizz[15][4] = 9'b111111111;
assign micromatrizz[15][5] = 9'b111111111;
assign micromatrizz[15][6] = 9'b111111111;
assign micromatrizz[15][7] = 9'b111111111;
assign micromatrizz[15][8] = 9'b111111111;
assign micromatrizz[15][9] = 9'b111111111;
assign micromatrizz[15][10] = 9'b111111111;
assign micromatrizz[15][11] = 9'b111111111;
assign micromatrizz[15][12] = 9'b111111111;
assign micromatrizz[15][13] = 9'b111111111;
assign micromatrizz[15][14] = 9'b111111111;
assign micromatrizz[15][15] = 9'b111111111;
assign micromatrizz[15][16] = 9'b111111111;
assign micromatrizz[15][17] = 9'b111111111;
assign micromatrizz[15][18] = 9'b111111111;
assign micromatrizz[15][19] = 9'b111111111;
assign micromatrizz[15][20] = 9'b111111111;
assign micromatrizz[15][21] = 9'b111111111;
assign micromatrizz[15][22] = 9'b111111111;
assign micromatrizz[15][23] = 9'b111111111;
assign micromatrizz[15][24] = 9'b111111111;
assign micromatrizz[15][25] = 9'b111111111;
assign micromatrizz[15][26] = 9'b111111111;
assign micromatrizz[15][27] = 9'b111111111;
assign micromatrizz[15][28] = 9'b111111111;
assign micromatrizz[15][29] = 9'b111111111;
assign micromatrizz[15][30] = 9'b111111111;
assign micromatrizz[15][31] = 9'b111111111;
assign micromatrizz[15][32] = 9'b111111111;
assign micromatrizz[15][33] = 9'b111111111;
assign micromatrizz[15][34] = 9'b111111111;
assign micromatrizz[15][35] = 9'b111111111;
assign micromatrizz[15][36] = 9'b111111111;
assign micromatrizz[15][37] = 9'b111111111;
assign micromatrizz[15][38] = 9'b111111111;
assign micromatrizz[15][39] = 9'b111111111;
assign micromatrizz[15][40] = 9'b111111111;
assign micromatrizz[15][41] = 9'b111111111;
assign micromatrizz[15][42] = 9'b111111111;
assign micromatrizz[15][43] = 9'b111111111;
assign micromatrizz[15][44] = 9'b111111111;
assign micromatrizz[15][45] = 9'b111111111;
assign micromatrizz[15][46] = 9'b111111111;
assign micromatrizz[15][47] = 9'b111111111;
assign micromatrizz[15][48] = 9'b111111111;
assign micromatrizz[15][49] = 9'b111111111;
assign micromatrizz[15][50] = 9'b111111111;
assign micromatrizz[15][51] = 9'b111111111;
assign micromatrizz[15][52] = 9'b111111111;
assign micromatrizz[15][53] = 9'b111111111;
assign micromatrizz[15][54] = 9'b111111111;
assign micromatrizz[15][55] = 9'b111111111;
assign micromatrizz[15][56] = 9'b111111111;
assign micromatrizz[15][57] = 9'b111111111;
assign micromatrizz[15][58] = 9'b111111111;
assign micromatrizz[15][59] = 9'b111111111;
assign micromatrizz[15][60] = 9'b111111111;
assign micromatrizz[15][61] = 9'b111111111;
assign micromatrizz[15][62] = 9'b111111111;
assign micromatrizz[15][63] = 9'b111111111;
assign micromatrizz[15][64] = 9'b111111111;
assign micromatrizz[15][65] = 9'b111111111;
assign micromatrizz[15][66] = 9'b111111111;
assign micromatrizz[15][67] = 9'b111111111;
assign micromatrizz[15][68] = 9'b111111111;
assign micromatrizz[15][69] = 9'b111111111;
assign micromatrizz[15][70] = 9'b111111111;
assign micromatrizz[15][71] = 9'b111111111;
assign micromatrizz[15][72] = 9'b111111111;
assign micromatrizz[15][73] = 9'b111111111;
assign micromatrizz[15][74] = 9'b111111111;
assign micromatrizz[15][75] = 9'b111111111;
assign micromatrizz[15][76] = 9'b111111111;
assign micromatrizz[15][77] = 9'b111111111;
assign micromatrizz[15][78] = 9'b111111111;
assign micromatrizz[15][79] = 9'b111111111;
assign micromatrizz[15][80] = 9'b111111111;
assign micromatrizz[15][81] = 9'b111111111;
assign micromatrizz[15][82] = 9'b111111111;
assign micromatrizz[15][83] = 9'b111111111;
assign micromatrizz[15][84] = 9'b111111111;
assign micromatrizz[15][85] = 9'b111111111;
assign micromatrizz[15][86] = 9'b111111111;
assign micromatrizz[15][87] = 9'b111111111;
assign micromatrizz[15][88] = 9'b111111111;
assign micromatrizz[15][89] = 9'b111111111;
assign micromatrizz[15][90] = 9'b111111111;
assign micromatrizz[15][91] = 9'b111111111;
assign micromatrizz[15][92] = 9'b111111111;
assign micromatrizz[15][93] = 9'b111111111;
assign micromatrizz[15][94] = 9'b111111111;
assign micromatrizz[15][95] = 9'b111111111;
assign micromatrizz[15][96] = 9'b111111111;
assign micromatrizz[15][97] = 9'b111111111;
assign micromatrizz[15][98] = 9'b111111111;
assign micromatrizz[15][99] = 9'b111111111;
assign micromatrizz[15][100] = 9'b111111111;
assign micromatrizz[15][101] = 9'b111111111;
assign micromatrizz[15][102] = 9'b111111111;
assign micromatrizz[15][103] = 9'b111111111;
assign micromatrizz[15][104] = 9'b111111111;
assign micromatrizz[15][105] = 9'b111111111;
assign micromatrizz[15][106] = 9'b111111111;
assign micromatrizz[15][107] = 9'b111111111;
assign micromatrizz[15][108] = 9'b111111111;
assign micromatrizz[15][109] = 9'b111111111;
assign micromatrizz[15][110] = 9'b111111111;
assign micromatrizz[15][111] = 9'b111111111;
assign micromatrizz[15][112] = 9'b111111111;
assign micromatrizz[15][113] = 9'b111111111;
assign micromatrizz[15][114] = 9'b111111111;
assign micromatrizz[15][115] = 9'b111111111;
assign micromatrizz[15][116] = 9'b111111111;
assign micromatrizz[15][117] = 9'b111111111;
assign micromatrizz[15][118] = 9'b111111111;
assign micromatrizz[15][119] = 9'b111111111;
assign micromatrizz[15][120] = 9'b111111111;
assign micromatrizz[15][121] = 9'b111111111;
assign micromatrizz[15][122] = 9'b111111111;
assign micromatrizz[15][123] = 9'b111111111;
assign micromatrizz[15][124] = 9'b111111111;
assign micromatrizz[15][125] = 9'b111111111;
assign micromatrizz[15][126] = 9'b111111111;
assign micromatrizz[15][127] = 9'b111111111;
assign micromatrizz[15][128] = 9'b111111111;
assign micromatrizz[15][129] = 9'b111111111;
assign micromatrizz[15][130] = 9'b111111111;
assign micromatrizz[15][131] = 9'b111111111;
assign micromatrizz[15][132] = 9'b111111111;
assign micromatrizz[15][133] = 9'b111111111;
assign micromatrizz[15][134] = 9'b111111111;
assign micromatrizz[15][135] = 9'b111111111;
assign micromatrizz[15][136] = 9'b111111111;
assign micromatrizz[15][137] = 9'b111111111;
assign micromatrizz[15][138] = 9'b111111111;
assign micromatrizz[15][139] = 9'b111111111;
assign micromatrizz[15][140] = 9'b111111111;
assign micromatrizz[15][141] = 9'b111111111;
assign micromatrizz[15][142] = 9'b111111111;
assign micromatrizz[15][143] = 9'b111111111;
assign micromatrizz[15][144] = 9'b111111111;
assign micromatrizz[15][145] = 9'b111111111;
assign micromatrizz[15][146] = 9'b111111111;
assign micromatrizz[15][147] = 9'b111111111;
assign micromatrizz[15][148] = 9'b111111111;
assign micromatrizz[15][149] = 9'b111111111;
assign micromatrizz[15][150] = 9'b111111111;
assign micromatrizz[15][151] = 9'b111111111;
assign micromatrizz[15][152] = 9'b111111111;
assign micromatrizz[15][153] = 9'b111111111;
assign micromatrizz[15][154] = 9'b111111111;
assign micromatrizz[15][155] = 9'b111111111;
assign micromatrizz[15][156] = 9'b111111111;
assign micromatrizz[15][157] = 9'b111111111;
assign micromatrizz[15][158] = 9'b111111111;
assign micromatrizz[15][159] = 9'b111111111;
assign micromatrizz[15][160] = 9'b111111111;
assign micromatrizz[15][161] = 9'b111111111;
assign micromatrizz[15][162] = 9'b111111111;
assign micromatrizz[15][163] = 9'b111111111;
assign micromatrizz[15][164] = 9'b111111111;
assign micromatrizz[15][165] = 9'b111111111;
assign micromatrizz[15][166] = 9'b111111111;
assign micromatrizz[15][167] = 9'b111111111;
assign micromatrizz[15][168] = 9'b111111111;
assign micromatrizz[15][169] = 9'b111111111;
assign micromatrizz[15][170] = 9'b111111111;
assign micromatrizz[15][171] = 9'b111111111;
assign micromatrizz[15][172] = 9'b111111111;
assign micromatrizz[15][173] = 9'b111111111;
assign micromatrizz[15][174] = 9'b111111111;
assign micromatrizz[15][175] = 9'b111111111;
assign micromatrizz[15][176] = 9'b111111111;
assign micromatrizz[15][177] = 9'b111111111;
assign micromatrizz[15][178] = 9'b111111111;
assign micromatrizz[15][179] = 9'b111111111;
assign micromatrizz[15][180] = 9'b111111111;
assign micromatrizz[15][181] = 9'b111111111;
assign micromatrizz[15][182] = 9'b111111111;
assign micromatrizz[15][183] = 9'b111111111;
assign micromatrizz[15][184] = 9'b111111111;
assign micromatrizz[15][185] = 9'b111111111;
assign micromatrizz[15][186] = 9'b111111111;
assign micromatrizz[15][187] = 9'b111111111;
assign micromatrizz[15][188] = 9'b111111111;
assign micromatrizz[15][189] = 9'b111111111;
assign micromatrizz[15][190] = 9'b111111111;
assign micromatrizz[15][191] = 9'b111111111;
assign micromatrizz[15][192] = 9'b111111111;
assign micromatrizz[15][193] = 9'b111111111;
assign micromatrizz[15][194] = 9'b111111111;
assign micromatrizz[15][195] = 9'b111111111;
assign micromatrizz[15][196] = 9'b111111111;
assign micromatrizz[15][197] = 9'b111111111;
assign micromatrizz[15][198] = 9'b111111111;
assign micromatrizz[15][199] = 9'b111111111;
assign micromatrizz[15][200] = 9'b111111111;
assign micromatrizz[15][201] = 9'b111111111;
assign micromatrizz[15][202] = 9'b111111111;
assign micromatrizz[15][203] = 9'b111111111;
assign micromatrizz[15][204] = 9'b111111111;
assign micromatrizz[15][205] = 9'b111111111;
assign micromatrizz[15][206] = 9'b111111111;
assign micromatrizz[15][207] = 9'b111111111;
assign micromatrizz[15][208] = 9'b111111111;
assign micromatrizz[15][209] = 9'b111111111;
assign micromatrizz[15][210] = 9'b111111111;
assign micromatrizz[15][211] = 9'b111111111;
assign micromatrizz[15][212] = 9'b111111111;
assign micromatrizz[15][213] = 9'b111111111;
assign micromatrizz[15][214] = 9'b111111111;
assign micromatrizz[15][215] = 9'b111111111;
assign micromatrizz[15][216] = 9'b111111111;
assign micromatrizz[15][217] = 9'b111111111;
assign micromatrizz[15][218] = 9'b111111111;
assign micromatrizz[15][219] = 9'b111111111;
assign micromatrizz[15][220] = 9'b111111111;
assign micromatrizz[15][221] = 9'b111111111;
assign micromatrizz[15][222] = 9'b111111111;
assign micromatrizz[15][223] = 9'b111111111;
assign micromatrizz[15][224] = 9'b111111111;
assign micromatrizz[15][225] = 9'b111111111;
assign micromatrizz[15][226] = 9'b111111111;
assign micromatrizz[15][227] = 9'b111111111;
assign micromatrizz[15][228] = 9'b111111111;
assign micromatrizz[15][229] = 9'b111111111;
assign micromatrizz[15][230] = 9'b111111111;
assign micromatrizz[15][231] = 9'b111111111;
assign micromatrizz[15][232] = 9'b111111111;
assign micromatrizz[15][233] = 9'b111111111;
assign micromatrizz[15][234] = 9'b111111111;
assign micromatrizz[15][235] = 9'b111111111;
assign micromatrizz[15][236] = 9'b111111111;
assign micromatrizz[15][237] = 9'b111111111;
assign micromatrizz[15][238] = 9'b111111111;
assign micromatrizz[15][239] = 9'b111111111;
assign micromatrizz[15][240] = 9'b111111111;
assign micromatrizz[15][241] = 9'b111111111;
assign micromatrizz[15][242] = 9'b111111111;
assign micromatrizz[15][243] = 9'b111111111;
assign micromatrizz[15][244] = 9'b111111111;
assign micromatrizz[15][245] = 9'b111111111;
assign micromatrizz[15][246] = 9'b111111111;
assign micromatrizz[15][247] = 9'b111111111;
assign micromatrizz[15][248] = 9'b111111111;
assign micromatrizz[15][249] = 9'b111111111;
assign micromatrizz[15][250] = 9'b111111111;
assign micromatrizz[15][251] = 9'b111111111;
assign micromatrizz[15][252] = 9'b111111111;
assign micromatrizz[15][253] = 9'b111111111;
assign micromatrizz[15][254] = 9'b111111111;
assign micromatrizz[15][255] = 9'b111111111;
assign micromatrizz[15][256] = 9'b111111111;
assign micromatrizz[15][257] = 9'b111111111;
assign micromatrizz[15][258] = 9'b111111111;
assign micromatrizz[15][259] = 9'b111111111;
assign micromatrizz[15][260] = 9'b111111111;
assign micromatrizz[15][261] = 9'b111111111;
assign micromatrizz[15][262] = 9'b111111111;
assign micromatrizz[15][263] = 9'b111111111;
assign micromatrizz[15][264] = 9'b111111111;
assign micromatrizz[15][265] = 9'b111111111;
assign micromatrizz[15][266] = 9'b111111111;
assign micromatrizz[15][267] = 9'b111111111;
assign micromatrizz[15][268] = 9'b111111111;
assign micromatrizz[15][269] = 9'b111111111;
assign micromatrizz[15][270] = 9'b111111111;
assign micromatrizz[15][271] = 9'b111111111;
assign micromatrizz[15][272] = 9'b111111111;
assign micromatrizz[15][273] = 9'b111111111;
assign micromatrizz[15][274] = 9'b111111111;
assign micromatrizz[15][275] = 9'b111111111;
assign micromatrizz[15][276] = 9'b111111111;
assign micromatrizz[15][277] = 9'b111111111;
assign micromatrizz[15][278] = 9'b111111111;
assign micromatrizz[15][279] = 9'b111111111;
assign micromatrizz[15][280] = 9'b111111111;
assign micromatrizz[15][281] = 9'b111111111;
assign micromatrizz[15][282] = 9'b111111111;
assign micromatrizz[15][283] = 9'b111111111;
assign micromatrizz[15][284] = 9'b111111111;
assign micromatrizz[15][285] = 9'b111111111;
assign micromatrizz[15][286] = 9'b111111111;
assign micromatrizz[15][287] = 9'b111111111;
assign micromatrizz[15][288] = 9'b111111111;
assign micromatrizz[15][289] = 9'b111111111;
assign micromatrizz[15][290] = 9'b111111111;
assign micromatrizz[15][291] = 9'b111111111;
assign micromatrizz[15][292] = 9'b111111111;
assign micromatrizz[15][293] = 9'b111111111;
assign micromatrizz[15][294] = 9'b111111111;
assign micromatrizz[15][295] = 9'b111111111;
assign micromatrizz[15][296] = 9'b111111111;
assign micromatrizz[15][297] = 9'b111111111;
assign micromatrizz[15][298] = 9'b111111111;
assign micromatrizz[15][299] = 9'b111111111;
assign micromatrizz[15][300] = 9'b111111111;
assign micromatrizz[15][301] = 9'b111111111;
assign micromatrizz[15][302] = 9'b111111111;
assign micromatrizz[15][303] = 9'b111111111;
assign micromatrizz[15][304] = 9'b111111111;
assign micromatrizz[15][305] = 9'b111111111;
assign micromatrizz[15][306] = 9'b111111111;
assign micromatrizz[15][307] = 9'b111111111;
assign micromatrizz[15][308] = 9'b111111111;
assign micromatrizz[15][309] = 9'b111111111;
assign micromatrizz[15][310] = 9'b111111111;
assign micromatrizz[15][311] = 9'b111111111;
assign micromatrizz[15][312] = 9'b111111111;
assign micromatrizz[15][313] = 9'b111111111;
assign micromatrizz[15][314] = 9'b111111111;
assign micromatrizz[15][315] = 9'b111111111;
assign micromatrizz[15][316] = 9'b111111111;
assign micromatrizz[15][317] = 9'b111111111;
assign micromatrizz[15][318] = 9'b111111111;
assign micromatrizz[15][319] = 9'b111111111;
assign micromatrizz[15][320] = 9'b111111111;
assign micromatrizz[15][321] = 9'b111111111;
assign micromatrizz[15][322] = 9'b111111111;
assign micromatrizz[15][323] = 9'b111111111;
assign micromatrizz[15][324] = 9'b111111111;
assign micromatrizz[15][325] = 9'b111111111;
assign micromatrizz[15][326] = 9'b111111111;
assign micromatrizz[15][327] = 9'b111111111;
assign micromatrizz[15][328] = 9'b111111111;
assign micromatrizz[15][329] = 9'b111111111;
assign micromatrizz[15][330] = 9'b111111111;
assign micromatrizz[15][331] = 9'b111111111;
assign micromatrizz[15][332] = 9'b111111111;
assign micromatrizz[15][333] = 9'b111111111;
assign micromatrizz[15][334] = 9'b111111111;
assign micromatrizz[15][335] = 9'b111111111;
assign micromatrizz[15][336] = 9'b111111111;
assign micromatrizz[15][337] = 9'b111111111;
assign micromatrizz[15][338] = 9'b111111111;
assign micromatrizz[15][339] = 9'b111111111;
assign micromatrizz[15][340] = 9'b111111111;
assign micromatrizz[15][341] = 9'b111111111;
assign micromatrizz[15][342] = 9'b111111111;
assign micromatrizz[15][343] = 9'b111111111;
assign micromatrizz[15][344] = 9'b111111111;
assign micromatrizz[15][345] = 9'b111111111;
assign micromatrizz[15][346] = 9'b111111111;
assign micromatrizz[15][347] = 9'b111111111;
assign micromatrizz[15][348] = 9'b111111111;
assign micromatrizz[15][349] = 9'b111111111;
assign micromatrizz[15][350] = 9'b111111111;
assign micromatrizz[15][351] = 9'b111111111;
assign micromatrizz[15][352] = 9'b111111111;
assign micromatrizz[15][353] = 9'b111111111;
assign micromatrizz[15][354] = 9'b111111111;
assign micromatrizz[15][355] = 9'b111111111;
assign micromatrizz[15][356] = 9'b111111111;
assign micromatrizz[15][357] = 9'b111111111;
assign micromatrizz[15][358] = 9'b111111111;
assign micromatrizz[15][359] = 9'b111111111;
assign micromatrizz[15][360] = 9'b111111111;
assign micromatrizz[15][361] = 9'b111111111;
assign micromatrizz[15][362] = 9'b111111111;
assign micromatrizz[15][363] = 9'b111111111;
assign micromatrizz[15][364] = 9'b111111111;
assign micromatrizz[15][365] = 9'b111111111;
assign micromatrizz[15][366] = 9'b111111111;
assign micromatrizz[15][367] = 9'b111111111;
assign micromatrizz[15][368] = 9'b111111111;
assign micromatrizz[15][369] = 9'b111111111;
assign micromatrizz[15][370] = 9'b111111111;
assign micromatrizz[15][371] = 9'b111111111;
assign micromatrizz[15][372] = 9'b111111111;
assign micromatrizz[15][373] = 9'b111111111;
assign micromatrizz[15][374] = 9'b111111111;
assign micromatrizz[15][375] = 9'b111111111;
assign micromatrizz[15][376] = 9'b111111111;
assign micromatrizz[15][377] = 9'b111111111;
assign micromatrizz[15][378] = 9'b111111111;
assign micromatrizz[15][379] = 9'b111111111;
assign micromatrizz[15][380] = 9'b111111111;
assign micromatrizz[15][381] = 9'b111111111;
assign micromatrizz[15][382] = 9'b111111111;
assign micromatrizz[15][383] = 9'b111111111;
assign micromatrizz[15][384] = 9'b111111111;
assign micromatrizz[15][385] = 9'b111111111;
assign micromatrizz[15][386] = 9'b111111111;
assign micromatrizz[15][387] = 9'b111111111;
assign micromatrizz[15][388] = 9'b111111111;
assign micromatrizz[15][389] = 9'b111111111;
assign micromatrizz[15][390] = 9'b111111111;
assign micromatrizz[15][391] = 9'b111111111;
assign micromatrizz[15][392] = 9'b111111111;
assign micromatrizz[15][393] = 9'b111111111;
assign micromatrizz[15][394] = 9'b111111111;
assign micromatrizz[15][395] = 9'b111111111;
assign micromatrizz[15][396] = 9'b111111111;
assign micromatrizz[15][397] = 9'b111111111;
assign micromatrizz[15][398] = 9'b111111111;
assign micromatrizz[15][399] = 9'b111111111;
assign micromatrizz[15][400] = 9'b111111111;
assign micromatrizz[15][401] = 9'b111111111;
assign micromatrizz[15][402] = 9'b111111111;
assign micromatrizz[15][403] = 9'b111111111;
assign micromatrizz[15][404] = 9'b111111111;
assign micromatrizz[15][405] = 9'b111111111;
assign micromatrizz[15][406] = 9'b111111111;
assign micromatrizz[15][407] = 9'b111111111;
assign micromatrizz[15][408] = 9'b111111111;
assign micromatrizz[15][409] = 9'b111111111;
assign micromatrizz[15][410] = 9'b111111111;
assign micromatrizz[15][411] = 9'b111111111;
assign micromatrizz[15][412] = 9'b111111111;
assign micromatrizz[15][413] = 9'b111111111;
assign micromatrizz[15][414] = 9'b111111111;
assign micromatrizz[15][415] = 9'b111111111;
assign micromatrizz[15][416] = 9'b111111111;
assign micromatrizz[15][417] = 9'b111111111;
assign micromatrizz[15][418] = 9'b111111111;
assign micromatrizz[15][419] = 9'b111111111;
assign micromatrizz[15][420] = 9'b111111111;
assign micromatrizz[15][421] = 9'b111111111;
assign micromatrizz[15][422] = 9'b111111111;
assign micromatrizz[15][423] = 9'b111111111;
assign micromatrizz[15][424] = 9'b111111111;
assign micromatrizz[15][425] = 9'b111111111;
assign micromatrizz[15][426] = 9'b111111111;
assign micromatrizz[15][427] = 9'b111111111;
assign micromatrizz[15][428] = 9'b111111111;
assign micromatrizz[15][429] = 9'b111111111;
assign micromatrizz[15][430] = 9'b111111111;
assign micromatrizz[15][431] = 9'b111111111;
assign micromatrizz[15][432] = 9'b111111111;
assign micromatrizz[15][433] = 9'b111111111;
assign micromatrizz[15][434] = 9'b111111111;
assign micromatrizz[15][435] = 9'b111111111;
assign micromatrizz[15][436] = 9'b111111111;
assign micromatrizz[15][437] = 9'b111111111;
assign micromatrizz[15][438] = 9'b111111111;
assign micromatrizz[15][439] = 9'b111111111;
assign micromatrizz[15][440] = 9'b111111111;
assign micromatrizz[15][441] = 9'b111111111;
assign micromatrizz[15][442] = 9'b111111111;
assign micromatrizz[15][443] = 9'b111111111;
assign micromatrizz[15][444] = 9'b111111111;
assign micromatrizz[15][445] = 9'b111111111;
assign micromatrizz[15][446] = 9'b111111111;
assign micromatrizz[15][447] = 9'b111111111;
assign micromatrizz[15][448] = 9'b111111111;
assign micromatrizz[15][449] = 9'b111111111;
assign micromatrizz[15][450] = 9'b111111111;
assign micromatrizz[15][451] = 9'b111111111;
assign micromatrizz[15][452] = 9'b111111111;
assign micromatrizz[15][453] = 9'b111111111;
assign micromatrizz[15][454] = 9'b111111111;
assign micromatrizz[15][455] = 9'b111111111;
assign micromatrizz[15][456] = 9'b111111111;
assign micromatrizz[15][457] = 9'b111111111;
assign micromatrizz[15][458] = 9'b111111111;
assign micromatrizz[15][459] = 9'b111111111;
assign micromatrizz[15][460] = 9'b111111111;
assign micromatrizz[15][461] = 9'b111111111;
assign micromatrizz[15][462] = 9'b111111111;
assign micromatrizz[15][463] = 9'b111111111;
assign micromatrizz[15][464] = 9'b111111111;
assign micromatrizz[15][465] = 9'b111111111;
assign micromatrizz[15][466] = 9'b111111111;
assign micromatrizz[15][467] = 9'b111111111;
assign micromatrizz[15][468] = 9'b111111111;
assign micromatrizz[15][469] = 9'b111111111;
assign micromatrizz[15][470] = 9'b111111111;
assign micromatrizz[15][471] = 9'b111111111;
assign micromatrizz[15][472] = 9'b111111111;
assign micromatrizz[15][473] = 9'b111111111;
assign micromatrizz[15][474] = 9'b111111111;
assign micromatrizz[15][475] = 9'b111111111;
assign micromatrizz[15][476] = 9'b111111111;
assign micromatrizz[15][477] = 9'b111111111;
assign micromatrizz[15][478] = 9'b111111111;
assign micromatrizz[15][479] = 9'b111111111;
assign micromatrizz[15][480] = 9'b111111111;
assign micromatrizz[15][481] = 9'b111111111;
assign micromatrizz[15][482] = 9'b111111111;
assign micromatrizz[15][483] = 9'b111111111;
assign micromatrizz[15][484] = 9'b111111111;
assign micromatrizz[15][485] = 9'b111111111;
assign micromatrizz[15][486] = 9'b111111111;
assign micromatrizz[15][487] = 9'b111111111;
assign micromatrizz[15][488] = 9'b111111111;
assign micromatrizz[15][489] = 9'b111111111;
assign micromatrizz[15][490] = 9'b111111111;
assign micromatrizz[15][491] = 9'b111111111;
assign micromatrizz[15][492] = 9'b111111111;
assign micromatrizz[15][493] = 9'b111111111;
assign micromatrizz[15][494] = 9'b111111111;
assign micromatrizz[15][495] = 9'b111111111;
assign micromatrizz[15][496] = 9'b111111111;
assign micromatrizz[15][497] = 9'b111111111;
assign micromatrizz[15][498] = 9'b111111111;
assign micromatrizz[15][499] = 9'b111111111;
assign micromatrizz[15][500] = 9'b111111111;
assign micromatrizz[15][501] = 9'b111111111;
assign micromatrizz[15][502] = 9'b111111111;
assign micromatrizz[15][503] = 9'b111111111;
assign micromatrizz[15][504] = 9'b111111111;
assign micromatrizz[15][505] = 9'b111111111;
assign micromatrizz[15][506] = 9'b111111111;
assign micromatrizz[15][507] = 9'b111111111;
assign micromatrizz[15][508] = 9'b111111111;
assign micromatrizz[15][509] = 9'b111111111;
assign micromatrizz[15][510] = 9'b111111111;
assign micromatrizz[15][511] = 9'b111111111;
assign micromatrizz[15][512] = 9'b111111111;
assign micromatrizz[15][513] = 9'b111111111;
assign micromatrizz[15][514] = 9'b111111111;
assign micromatrizz[15][515] = 9'b111111111;
assign micromatrizz[15][516] = 9'b111111111;
assign micromatrizz[15][517] = 9'b111111111;
assign micromatrizz[15][518] = 9'b111111111;
assign micromatrizz[15][519] = 9'b111111111;
assign micromatrizz[15][520] = 9'b111111111;
assign micromatrizz[15][521] = 9'b111111111;
assign micromatrizz[15][522] = 9'b111111111;
assign micromatrizz[15][523] = 9'b111111111;
assign micromatrizz[15][524] = 9'b111111111;
assign micromatrizz[15][525] = 9'b111111111;
assign micromatrizz[15][526] = 9'b111111111;
assign micromatrizz[15][527] = 9'b111111111;
assign micromatrizz[15][528] = 9'b111111111;
assign micromatrizz[15][529] = 9'b111111111;
assign micromatrizz[15][530] = 9'b111111111;
assign micromatrizz[15][531] = 9'b111111111;
assign micromatrizz[15][532] = 9'b111111111;
assign micromatrizz[15][533] = 9'b111111111;
assign micromatrizz[15][534] = 9'b111111111;
assign micromatrizz[15][535] = 9'b111111111;
assign micromatrizz[15][536] = 9'b111111111;
assign micromatrizz[15][537] = 9'b111111111;
assign micromatrizz[15][538] = 9'b111111111;
assign micromatrizz[15][539] = 9'b111111111;
assign micromatrizz[15][540] = 9'b111111111;
assign micromatrizz[15][541] = 9'b111111111;
assign micromatrizz[15][542] = 9'b111111111;
assign micromatrizz[15][543] = 9'b111111111;
assign micromatrizz[15][544] = 9'b111111111;
assign micromatrizz[15][545] = 9'b111111111;
assign micromatrizz[15][546] = 9'b111111111;
assign micromatrizz[15][547] = 9'b111111111;
assign micromatrizz[15][548] = 9'b111111111;
assign micromatrizz[15][549] = 9'b111111111;
assign micromatrizz[15][550] = 9'b111111111;
assign micromatrizz[15][551] = 9'b111111111;
assign micromatrizz[15][552] = 9'b111111111;
assign micromatrizz[15][553] = 9'b111111111;
assign micromatrizz[15][554] = 9'b111111111;
assign micromatrizz[15][555] = 9'b111111111;
assign micromatrizz[15][556] = 9'b111111111;
assign micromatrizz[15][557] = 9'b111111111;
assign micromatrizz[15][558] = 9'b111111111;
assign micromatrizz[15][559] = 9'b111111111;
assign micromatrizz[15][560] = 9'b111111111;
assign micromatrizz[15][561] = 9'b111111111;
assign micromatrizz[15][562] = 9'b111111111;
assign micromatrizz[15][563] = 9'b111111111;
assign micromatrizz[15][564] = 9'b111111111;
assign micromatrizz[15][565] = 9'b111111111;
assign micromatrizz[15][566] = 9'b111111111;
assign micromatrizz[15][567] = 9'b111111111;
assign micromatrizz[15][568] = 9'b111111111;
assign micromatrizz[15][569] = 9'b111111111;
assign micromatrizz[15][570] = 9'b111111111;
assign micromatrizz[15][571] = 9'b111111111;
assign micromatrizz[15][572] = 9'b111111111;
assign micromatrizz[15][573] = 9'b111111111;
assign micromatrizz[15][574] = 9'b111111111;
assign micromatrizz[15][575] = 9'b111111111;
assign micromatrizz[15][576] = 9'b111111111;
assign micromatrizz[15][577] = 9'b111111111;
assign micromatrizz[15][578] = 9'b111111111;
assign micromatrizz[15][579] = 9'b111111111;
assign micromatrizz[15][580] = 9'b111111111;
assign micromatrizz[15][581] = 9'b111111111;
assign micromatrizz[15][582] = 9'b111111111;
assign micromatrizz[15][583] = 9'b111111111;
assign micromatrizz[15][584] = 9'b111111111;
assign micromatrizz[15][585] = 9'b111111111;
assign micromatrizz[15][586] = 9'b111111111;
assign micromatrizz[15][587] = 9'b111111111;
assign micromatrizz[15][588] = 9'b111111111;
assign micromatrizz[15][589] = 9'b111111111;
assign micromatrizz[15][590] = 9'b111111111;
assign micromatrizz[15][591] = 9'b111111111;
assign micromatrizz[15][592] = 9'b111111111;
assign micromatrizz[15][593] = 9'b111111111;
assign micromatrizz[15][594] = 9'b111111111;
assign micromatrizz[15][595] = 9'b111111111;
assign micromatrizz[15][596] = 9'b111111111;
assign micromatrizz[15][597] = 9'b111111111;
assign micromatrizz[15][598] = 9'b111111111;
assign micromatrizz[15][599] = 9'b111111111;
assign micromatrizz[15][600] = 9'b111111111;
assign micromatrizz[15][601] = 9'b111111111;
assign micromatrizz[15][602] = 9'b111111111;
assign micromatrizz[15][603] = 9'b111111111;
assign micromatrizz[15][604] = 9'b111111111;
assign micromatrizz[15][605] = 9'b111111111;
assign micromatrizz[15][606] = 9'b111111111;
assign micromatrizz[15][607] = 9'b111111111;
assign micromatrizz[15][608] = 9'b111111111;
assign micromatrizz[15][609] = 9'b111111111;
assign micromatrizz[15][610] = 9'b111111111;
assign micromatrizz[15][611] = 9'b111111111;
assign micromatrizz[15][612] = 9'b111111111;
assign micromatrizz[15][613] = 9'b111111111;
assign micromatrizz[15][614] = 9'b111111111;
assign micromatrizz[15][615] = 9'b111111111;
assign micromatrizz[15][616] = 9'b111111111;
assign micromatrizz[15][617] = 9'b111111111;
assign micromatrizz[15][618] = 9'b111111111;
assign micromatrizz[15][619] = 9'b111111111;
assign micromatrizz[15][620] = 9'b111111111;
assign micromatrizz[15][621] = 9'b111111111;
assign micromatrizz[15][622] = 9'b111111111;
assign micromatrizz[15][623] = 9'b111111111;
assign micromatrizz[15][624] = 9'b111111111;
assign micromatrizz[15][625] = 9'b111111111;
assign micromatrizz[15][626] = 9'b111111111;
assign micromatrizz[15][627] = 9'b111111111;
assign micromatrizz[15][628] = 9'b111111111;
assign micromatrizz[15][629] = 9'b111111111;
assign micromatrizz[15][630] = 9'b111111111;
assign micromatrizz[15][631] = 9'b111111111;
assign micromatrizz[15][632] = 9'b111111111;
assign micromatrizz[15][633] = 9'b111111111;
assign micromatrizz[15][634] = 9'b111111111;
assign micromatrizz[15][635] = 9'b111111111;
assign micromatrizz[15][636] = 9'b111111111;
assign micromatrizz[15][637] = 9'b111111111;
assign micromatrizz[15][638] = 9'b111111111;
assign micromatrizz[15][639] = 9'b111111111;
assign micromatrizz[16][0] = 9'b111111111;
assign micromatrizz[16][1] = 9'b111111111;
assign micromatrizz[16][2] = 9'b111111111;
assign micromatrizz[16][3] = 9'b111111111;
assign micromatrizz[16][4] = 9'b111111111;
assign micromatrizz[16][5] = 9'b111111111;
assign micromatrizz[16][6] = 9'b111111111;
assign micromatrizz[16][7] = 9'b111111111;
assign micromatrizz[16][8] = 9'b111111111;
assign micromatrizz[16][9] = 9'b111111111;
assign micromatrizz[16][10] = 9'b111111111;
assign micromatrizz[16][11] = 9'b111111111;
assign micromatrizz[16][12] = 9'b111111111;
assign micromatrizz[16][13] = 9'b111111111;
assign micromatrizz[16][14] = 9'b111111111;
assign micromatrizz[16][15] = 9'b111111111;
assign micromatrizz[16][16] = 9'b111111111;
assign micromatrizz[16][17] = 9'b111111111;
assign micromatrizz[16][18] = 9'b111111111;
assign micromatrizz[16][19] = 9'b111111111;
assign micromatrizz[16][20] = 9'b111111111;
assign micromatrizz[16][21] = 9'b111111111;
assign micromatrizz[16][22] = 9'b111111111;
assign micromatrizz[16][23] = 9'b111111111;
assign micromatrizz[16][24] = 9'b111111111;
assign micromatrizz[16][25] = 9'b111111111;
assign micromatrizz[16][26] = 9'b111111111;
assign micromatrizz[16][27] = 9'b111111111;
assign micromatrizz[16][28] = 9'b111111111;
assign micromatrizz[16][29] = 9'b111111111;
assign micromatrizz[16][30] = 9'b111111111;
assign micromatrizz[16][31] = 9'b111111111;
assign micromatrizz[16][32] = 9'b111111111;
assign micromatrizz[16][33] = 9'b111111111;
assign micromatrizz[16][34] = 9'b111111111;
assign micromatrizz[16][35] = 9'b111111111;
assign micromatrizz[16][36] = 9'b111111111;
assign micromatrizz[16][37] = 9'b111111111;
assign micromatrizz[16][38] = 9'b111111111;
assign micromatrizz[16][39] = 9'b111111111;
assign micromatrizz[16][40] = 9'b111111111;
assign micromatrizz[16][41] = 9'b111111111;
assign micromatrizz[16][42] = 9'b111111111;
assign micromatrizz[16][43] = 9'b111111111;
assign micromatrizz[16][44] = 9'b111111111;
assign micromatrizz[16][45] = 9'b111111111;
assign micromatrizz[16][46] = 9'b111111111;
assign micromatrizz[16][47] = 9'b111111111;
assign micromatrizz[16][48] = 9'b111111111;
assign micromatrizz[16][49] = 9'b111111111;
assign micromatrizz[16][50] = 9'b111111111;
assign micromatrizz[16][51] = 9'b111111111;
assign micromatrizz[16][52] = 9'b111111111;
assign micromatrizz[16][53] = 9'b111111111;
assign micromatrizz[16][54] = 9'b111111111;
assign micromatrizz[16][55] = 9'b111111111;
assign micromatrizz[16][56] = 9'b111111111;
assign micromatrizz[16][57] = 9'b111111111;
assign micromatrizz[16][58] = 9'b111111111;
assign micromatrizz[16][59] = 9'b111111111;
assign micromatrizz[16][60] = 9'b111111111;
assign micromatrizz[16][61] = 9'b111111111;
assign micromatrizz[16][62] = 9'b111111111;
assign micromatrizz[16][63] = 9'b111111111;
assign micromatrizz[16][64] = 9'b111111111;
assign micromatrizz[16][65] = 9'b111111111;
assign micromatrizz[16][66] = 9'b111111111;
assign micromatrizz[16][67] = 9'b111111111;
assign micromatrizz[16][68] = 9'b111111111;
assign micromatrizz[16][69] = 9'b111111111;
assign micromatrizz[16][70] = 9'b111111111;
assign micromatrizz[16][71] = 9'b111111111;
assign micromatrizz[16][72] = 9'b111111111;
assign micromatrizz[16][73] = 9'b111111111;
assign micromatrizz[16][74] = 9'b111111111;
assign micromatrizz[16][75] = 9'b111111111;
assign micromatrizz[16][76] = 9'b111111111;
assign micromatrizz[16][77] = 9'b111111111;
assign micromatrizz[16][78] = 9'b111111111;
assign micromatrizz[16][79] = 9'b111111111;
assign micromatrizz[16][80] = 9'b111111111;
assign micromatrizz[16][81] = 9'b111111111;
assign micromatrizz[16][82] = 9'b111111111;
assign micromatrizz[16][83] = 9'b111111111;
assign micromatrizz[16][84] = 9'b111111111;
assign micromatrizz[16][85] = 9'b111111111;
assign micromatrizz[16][86] = 9'b111111111;
assign micromatrizz[16][87] = 9'b111111111;
assign micromatrizz[16][88] = 9'b111111111;
assign micromatrizz[16][89] = 9'b111111111;
assign micromatrizz[16][90] = 9'b111111111;
assign micromatrizz[16][91] = 9'b111111111;
assign micromatrizz[16][92] = 9'b111111111;
assign micromatrizz[16][93] = 9'b111111111;
assign micromatrizz[16][94] = 9'b111111111;
assign micromatrizz[16][95] = 9'b111111111;
assign micromatrizz[16][96] = 9'b111111111;
assign micromatrizz[16][97] = 9'b111111111;
assign micromatrizz[16][98] = 9'b111111111;
assign micromatrizz[16][99] = 9'b111111111;
assign micromatrizz[16][100] = 9'b111111111;
assign micromatrizz[16][101] = 9'b111111111;
assign micromatrizz[16][102] = 9'b111111111;
assign micromatrizz[16][103] = 9'b111111111;
assign micromatrizz[16][104] = 9'b111111111;
assign micromatrizz[16][105] = 9'b111111111;
assign micromatrizz[16][106] = 9'b111111111;
assign micromatrizz[16][107] = 9'b111111111;
assign micromatrizz[16][108] = 9'b111111111;
assign micromatrizz[16][109] = 9'b111111111;
assign micromatrizz[16][110] = 9'b111111111;
assign micromatrizz[16][111] = 9'b111111111;
assign micromatrizz[16][112] = 9'b111111111;
assign micromatrizz[16][113] = 9'b111111111;
assign micromatrizz[16][114] = 9'b111111111;
assign micromatrizz[16][115] = 9'b111111111;
assign micromatrizz[16][116] = 9'b111111111;
assign micromatrizz[16][117] = 9'b111111111;
assign micromatrizz[16][118] = 9'b111111111;
assign micromatrizz[16][119] = 9'b111111111;
assign micromatrizz[16][120] = 9'b111111111;
assign micromatrizz[16][121] = 9'b111111111;
assign micromatrizz[16][122] = 9'b111111111;
assign micromatrizz[16][123] = 9'b111111111;
assign micromatrizz[16][124] = 9'b111111111;
assign micromatrizz[16][125] = 9'b111111111;
assign micromatrizz[16][126] = 9'b111111111;
assign micromatrizz[16][127] = 9'b111111111;
assign micromatrizz[16][128] = 9'b111111111;
assign micromatrizz[16][129] = 9'b111111111;
assign micromatrizz[16][130] = 9'b111111111;
assign micromatrizz[16][131] = 9'b111111111;
assign micromatrizz[16][132] = 9'b111111111;
assign micromatrizz[16][133] = 9'b111111111;
assign micromatrizz[16][134] = 9'b111111111;
assign micromatrizz[16][135] = 9'b111111111;
assign micromatrizz[16][136] = 9'b111111111;
assign micromatrizz[16][137] = 9'b111111111;
assign micromatrizz[16][138] = 9'b111111111;
assign micromatrizz[16][139] = 9'b111111111;
assign micromatrizz[16][140] = 9'b111111111;
assign micromatrizz[16][141] = 9'b111111111;
assign micromatrizz[16][142] = 9'b111111111;
assign micromatrizz[16][143] = 9'b111111111;
assign micromatrizz[16][144] = 9'b111111111;
assign micromatrizz[16][145] = 9'b111111111;
assign micromatrizz[16][146] = 9'b111111111;
assign micromatrizz[16][147] = 9'b111111111;
assign micromatrizz[16][148] = 9'b111111111;
assign micromatrizz[16][149] = 9'b111111111;
assign micromatrizz[16][150] = 9'b111111111;
assign micromatrizz[16][151] = 9'b111111111;
assign micromatrizz[16][152] = 9'b111111111;
assign micromatrizz[16][153] = 9'b111111111;
assign micromatrizz[16][154] = 9'b111111111;
assign micromatrizz[16][155] = 9'b111111111;
assign micromatrizz[16][156] = 9'b111111111;
assign micromatrizz[16][157] = 9'b111111111;
assign micromatrizz[16][158] = 9'b111111111;
assign micromatrizz[16][159] = 9'b111111111;
assign micromatrizz[16][160] = 9'b111111111;
assign micromatrizz[16][161] = 9'b111111111;
assign micromatrizz[16][162] = 9'b111111111;
assign micromatrizz[16][163] = 9'b111111111;
assign micromatrizz[16][164] = 9'b111111111;
assign micromatrizz[16][165] = 9'b111111111;
assign micromatrizz[16][166] = 9'b111111111;
assign micromatrizz[16][167] = 9'b111111111;
assign micromatrizz[16][168] = 9'b111111111;
assign micromatrizz[16][169] = 9'b111111111;
assign micromatrizz[16][170] = 9'b111111111;
assign micromatrizz[16][171] = 9'b111111111;
assign micromatrizz[16][172] = 9'b111111111;
assign micromatrizz[16][173] = 9'b111111111;
assign micromatrizz[16][174] = 9'b111111111;
assign micromatrizz[16][175] = 9'b111111111;
assign micromatrizz[16][176] = 9'b111111111;
assign micromatrizz[16][177] = 9'b111111111;
assign micromatrizz[16][178] = 9'b111111111;
assign micromatrizz[16][179] = 9'b111111111;
assign micromatrizz[16][180] = 9'b111111111;
assign micromatrizz[16][181] = 9'b111111111;
assign micromatrizz[16][182] = 9'b111111111;
assign micromatrizz[16][183] = 9'b111111111;
assign micromatrizz[16][184] = 9'b111111111;
assign micromatrizz[16][185] = 9'b111111111;
assign micromatrizz[16][186] = 9'b111111111;
assign micromatrizz[16][187] = 9'b111111111;
assign micromatrizz[16][188] = 9'b111111111;
assign micromatrizz[16][189] = 9'b111111111;
assign micromatrizz[16][190] = 9'b111111111;
assign micromatrizz[16][191] = 9'b111111111;
assign micromatrizz[16][192] = 9'b111111111;
assign micromatrizz[16][193] = 9'b111111111;
assign micromatrizz[16][194] = 9'b111111111;
assign micromatrizz[16][195] = 9'b111111111;
assign micromatrizz[16][196] = 9'b111111111;
assign micromatrizz[16][197] = 9'b111111111;
assign micromatrizz[16][198] = 9'b111111111;
assign micromatrizz[16][199] = 9'b111111111;
assign micromatrizz[16][200] = 9'b111111111;
assign micromatrizz[16][201] = 9'b111111111;
assign micromatrizz[16][202] = 9'b111111111;
assign micromatrizz[16][203] = 9'b111111111;
assign micromatrizz[16][204] = 9'b111111111;
assign micromatrizz[16][205] = 9'b111111111;
assign micromatrizz[16][206] = 9'b111111111;
assign micromatrizz[16][207] = 9'b111111111;
assign micromatrizz[16][208] = 9'b111111111;
assign micromatrizz[16][209] = 9'b111111111;
assign micromatrizz[16][210] = 9'b111111111;
assign micromatrizz[16][211] = 9'b111111111;
assign micromatrizz[16][212] = 9'b111111111;
assign micromatrizz[16][213] = 9'b111111111;
assign micromatrizz[16][214] = 9'b111111111;
assign micromatrizz[16][215] = 9'b111111111;
assign micromatrizz[16][216] = 9'b111111111;
assign micromatrizz[16][217] = 9'b111111111;
assign micromatrizz[16][218] = 9'b111111111;
assign micromatrizz[16][219] = 9'b111111111;
assign micromatrizz[16][220] = 9'b111111111;
assign micromatrizz[16][221] = 9'b111111111;
assign micromatrizz[16][222] = 9'b111111111;
assign micromatrizz[16][223] = 9'b111111111;
assign micromatrizz[16][224] = 9'b111111111;
assign micromatrizz[16][225] = 9'b111111111;
assign micromatrizz[16][226] = 9'b111111111;
assign micromatrizz[16][227] = 9'b111111111;
assign micromatrizz[16][228] = 9'b111111111;
assign micromatrizz[16][229] = 9'b111111111;
assign micromatrizz[16][230] = 9'b111111111;
assign micromatrizz[16][231] = 9'b111111111;
assign micromatrizz[16][232] = 9'b111111111;
assign micromatrizz[16][233] = 9'b111111111;
assign micromatrizz[16][234] = 9'b111111111;
assign micromatrizz[16][235] = 9'b111111111;
assign micromatrizz[16][236] = 9'b111111111;
assign micromatrizz[16][237] = 9'b111111111;
assign micromatrizz[16][238] = 9'b111111111;
assign micromatrizz[16][239] = 9'b111111111;
assign micromatrizz[16][240] = 9'b111111111;
assign micromatrizz[16][241] = 9'b111111111;
assign micromatrizz[16][242] = 9'b111111111;
assign micromatrizz[16][243] = 9'b111111111;
assign micromatrizz[16][244] = 9'b111111111;
assign micromatrizz[16][245] = 9'b111111111;
assign micromatrizz[16][246] = 9'b111111111;
assign micromatrizz[16][247] = 9'b111111111;
assign micromatrizz[16][248] = 9'b111111111;
assign micromatrizz[16][249] = 9'b111111111;
assign micromatrizz[16][250] = 9'b111111111;
assign micromatrizz[16][251] = 9'b111111111;
assign micromatrizz[16][252] = 9'b111111111;
assign micromatrizz[16][253] = 9'b111111111;
assign micromatrizz[16][254] = 9'b111111111;
assign micromatrizz[16][255] = 9'b111111111;
assign micromatrizz[16][256] = 9'b111111111;
assign micromatrizz[16][257] = 9'b111111111;
assign micromatrizz[16][258] = 9'b111111111;
assign micromatrizz[16][259] = 9'b111111111;
assign micromatrizz[16][260] = 9'b111111111;
assign micromatrizz[16][261] = 9'b111111111;
assign micromatrizz[16][262] = 9'b111111111;
assign micromatrizz[16][263] = 9'b111111111;
assign micromatrizz[16][264] = 9'b111111111;
assign micromatrizz[16][265] = 9'b111111111;
assign micromatrizz[16][266] = 9'b111111111;
assign micromatrizz[16][267] = 9'b111111111;
assign micromatrizz[16][268] = 9'b111111111;
assign micromatrizz[16][269] = 9'b111111111;
assign micromatrizz[16][270] = 9'b111111111;
assign micromatrizz[16][271] = 9'b111111111;
assign micromatrizz[16][272] = 9'b111111111;
assign micromatrizz[16][273] = 9'b111111111;
assign micromatrizz[16][274] = 9'b111111111;
assign micromatrizz[16][275] = 9'b111111111;
assign micromatrizz[16][276] = 9'b111111111;
assign micromatrizz[16][277] = 9'b111111111;
assign micromatrizz[16][278] = 9'b111111111;
assign micromatrizz[16][279] = 9'b111111111;
assign micromatrizz[16][280] = 9'b111111111;
assign micromatrizz[16][281] = 9'b111111111;
assign micromatrizz[16][282] = 9'b111111111;
assign micromatrizz[16][283] = 9'b111111111;
assign micromatrizz[16][284] = 9'b111111111;
assign micromatrizz[16][285] = 9'b111111111;
assign micromatrizz[16][286] = 9'b111111111;
assign micromatrizz[16][287] = 9'b111111111;
assign micromatrizz[16][288] = 9'b111111111;
assign micromatrizz[16][289] = 9'b111111111;
assign micromatrizz[16][290] = 9'b111111111;
assign micromatrizz[16][291] = 9'b111111111;
assign micromatrizz[16][292] = 9'b111111111;
assign micromatrizz[16][293] = 9'b111111111;
assign micromatrizz[16][294] = 9'b111111111;
assign micromatrizz[16][295] = 9'b111111111;
assign micromatrizz[16][296] = 9'b111111111;
assign micromatrizz[16][297] = 9'b111111111;
assign micromatrizz[16][298] = 9'b111111111;
assign micromatrizz[16][299] = 9'b111111111;
assign micromatrizz[16][300] = 9'b111111111;
assign micromatrizz[16][301] = 9'b111111111;
assign micromatrizz[16][302] = 9'b111111111;
assign micromatrizz[16][303] = 9'b111111111;
assign micromatrizz[16][304] = 9'b111111111;
assign micromatrizz[16][305] = 9'b111111111;
assign micromatrizz[16][306] = 9'b111111111;
assign micromatrizz[16][307] = 9'b111111111;
assign micromatrizz[16][308] = 9'b111111111;
assign micromatrizz[16][309] = 9'b111111111;
assign micromatrizz[16][310] = 9'b111111111;
assign micromatrizz[16][311] = 9'b111111111;
assign micromatrizz[16][312] = 9'b111111111;
assign micromatrizz[16][313] = 9'b111111111;
assign micromatrizz[16][314] = 9'b111111111;
assign micromatrizz[16][315] = 9'b111111111;
assign micromatrizz[16][316] = 9'b111111111;
assign micromatrizz[16][317] = 9'b111111111;
assign micromatrizz[16][318] = 9'b111111111;
assign micromatrizz[16][319] = 9'b111111111;
assign micromatrizz[16][320] = 9'b111111111;
assign micromatrizz[16][321] = 9'b111111111;
assign micromatrizz[16][322] = 9'b111111111;
assign micromatrizz[16][323] = 9'b111111111;
assign micromatrizz[16][324] = 9'b111111111;
assign micromatrizz[16][325] = 9'b111111111;
assign micromatrizz[16][326] = 9'b111111111;
assign micromatrizz[16][327] = 9'b111111111;
assign micromatrizz[16][328] = 9'b111111111;
assign micromatrizz[16][329] = 9'b111111111;
assign micromatrizz[16][330] = 9'b111111111;
assign micromatrizz[16][331] = 9'b111111111;
assign micromatrizz[16][332] = 9'b111111111;
assign micromatrizz[16][333] = 9'b111111111;
assign micromatrizz[16][334] = 9'b111111111;
assign micromatrizz[16][335] = 9'b111111111;
assign micromatrizz[16][336] = 9'b111111111;
assign micromatrizz[16][337] = 9'b111111111;
assign micromatrizz[16][338] = 9'b111111111;
assign micromatrizz[16][339] = 9'b111111111;
assign micromatrizz[16][340] = 9'b111111111;
assign micromatrizz[16][341] = 9'b111111111;
assign micromatrizz[16][342] = 9'b111111111;
assign micromatrizz[16][343] = 9'b111111111;
assign micromatrizz[16][344] = 9'b111111111;
assign micromatrizz[16][345] = 9'b111111111;
assign micromatrizz[16][346] = 9'b111111111;
assign micromatrizz[16][347] = 9'b111111111;
assign micromatrizz[16][348] = 9'b111111111;
assign micromatrizz[16][349] = 9'b111111111;
assign micromatrizz[16][350] = 9'b111111111;
assign micromatrizz[16][351] = 9'b111111111;
assign micromatrizz[16][352] = 9'b111111111;
assign micromatrizz[16][353] = 9'b111111111;
assign micromatrizz[16][354] = 9'b111111111;
assign micromatrizz[16][355] = 9'b111111111;
assign micromatrizz[16][356] = 9'b111111111;
assign micromatrizz[16][357] = 9'b111111111;
assign micromatrizz[16][358] = 9'b111111111;
assign micromatrizz[16][359] = 9'b111111111;
assign micromatrizz[16][360] = 9'b111111111;
assign micromatrizz[16][361] = 9'b111111111;
assign micromatrizz[16][362] = 9'b111111111;
assign micromatrizz[16][363] = 9'b111111111;
assign micromatrizz[16][364] = 9'b111111111;
assign micromatrizz[16][365] = 9'b111111111;
assign micromatrizz[16][366] = 9'b111111111;
assign micromatrizz[16][367] = 9'b111111111;
assign micromatrizz[16][368] = 9'b111111111;
assign micromatrizz[16][369] = 9'b111111111;
assign micromatrizz[16][370] = 9'b111111111;
assign micromatrizz[16][371] = 9'b111111111;
assign micromatrizz[16][372] = 9'b111111111;
assign micromatrizz[16][373] = 9'b111111111;
assign micromatrizz[16][374] = 9'b111111111;
assign micromatrizz[16][375] = 9'b111111111;
assign micromatrizz[16][376] = 9'b111111111;
assign micromatrizz[16][377] = 9'b111111111;
assign micromatrizz[16][378] = 9'b111111111;
assign micromatrizz[16][379] = 9'b111111111;
assign micromatrizz[16][380] = 9'b111111111;
assign micromatrizz[16][381] = 9'b111111111;
assign micromatrizz[16][382] = 9'b111111111;
assign micromatrizz[16][383] = 9'b111111111;
assign micromatrizz[16][384] = 9'b111111111;
assign micromatrizz[16][385] = 9'b111111111;
assign micromatrizz[16][386] = 9'b111111111;
assign micromatrizz[16][387] = 9'b111111111;
assign micromatrizz[16][388] = 9'b111111111;
assign micromatrizz[16][389] = 9'b111111111;
assign micromatrizz[16][390] = 9'b111111111;
assign micromatrizz[16][391] = 9'b111111111;
assign micromatrizz[16][392] = 9'b111111111;
assign micromatrizz[16][393] = 9'b111111111;
assign micromatrizz[16][394] = 9'b111111111;
assign micromatrizz[16][395] = 9'b111111111;
assign micromatrizz[16][396] = 9'b111111111;
assign micromatrizz[16][397] = 9'b111111111;
assign micromatrizz[16][398] = 9'b111111111;
assign micromatrizz[16][399] = 9'b111111111;
assign micromatrizz[16][400] = 9'b111111111;
assign micromatrizz[16][401] = 9'b111111111;
assign micromatrizz[16][402] = 9'b111111111;
assign micromatrizz[16][403] = 9'b111111111;
assign micromatrizz[16][404] = 9'b111111111;
assign micromatrizz[16][405] = 9'b111111111;
assign micromatrizz[16][406] = 9'b111111111;
assign micromatrizz[16][407] = 9'b111111111;
assign micromatrizz[16][408] = 9'b111111111;
assign micromatrizz[16][409] = 9'b111111111;
assign micromatrizz[16][410] = 9'b111111111;
assign micromatrizz[16][411] = 9'b111111111;
assign micromatrizz[16][412] = 9'b111111111;
assign micromatrizz[16][413] = 9'b111111111;
assign micromatrizz[16][414] = 9'b111111111;
assign micromatrizz[16][415] = 9'b111111111;
assign micromatrizz[16][416] = 9'b111111111;
assign micromatrizz[16][417] = 9'b111111111;
assign micromatrizz[16][418] = 9'b111111111;
assign micromatrizz[16][419] = 9'b111111111;
assign micromatrizz[16][420] = 9'b111111111;
assign micromatrizz[16][421] = 9'b111111111;
assign micromatrizz[16][422] = 9'b111111111;
assign micromatrizz[16][423] = 9'b111111111;
assign micromatrizz[16][424] = 9'b111111111;
assign micromatrizz[16][425] = 9'b111111111;
assign micromatrizz[16][426] = 9'b111111111;
assign micromatrizz[16][427] = 9'b111111111;
assign micromatrizz[16][428] = 9'b111111111;
assign micromatrizz[16][429] = 9'b111111111;
assign micromatrizz[16][430] = 9'b111111111;
assign micromatrizz[16][431] = 9'b111111111;
assign micromatrizz[16][432] = 9'b111111111;
assign micromatrizz[16][433] = 9'b111111111;
assign micromatrizz[16][434] = 9'b111111111;
assign micromatrizz[16][435] = 9'b111111111;
assign micromatrizz[16][436] = 9'b111111111;
assign micromatrizz[16][437] = 9'b111111111;
assign micromatrizz[16][438] = 9'b111111111;
assign micromatrizz[16][439] = 9'b111111111;
assign micromatrizz[16][440] = 9'b111111111;
assign micromatrizz[16][441] = 9'b111111111;
assign micromatrizz[16][442] = 9'b111111111;
assign micromatrizz[16][443] = 9'b111111111;
assign micromatrizz[16][444] = 9'b111111111;
assign micromatrizz[16][445] = 9'b111111111;
assign micromatrizz[16][446] = 9'b111111111;
assign micromatrizz[16][447] = 9'b111111111;
assign micromatrizz[16][448] = 9'b111111111;
assign micromatrizz[16][449] = 9'b111111111;
assign micromatrizz[16][450] = 9'b111111111;
assign micromatrizz[16][451] = 9'b111111111;
assign micromatrizz[16][452] = 9'b111111111;
assign micromatrizz[16][453] = 9'b111111111;
assign micromatrizz[16][454] = 9'b111111111;
assign micromatrizz[16][455] = 9'b111111111;
assign micromatrizz[16][456] = 9'b111111111;
assign micromatrizz[16][457] = 9'b111111111;
assign micromatrizz[16][458] = 9'b111111111;
assign micromatrizz[16][459] = 9'b111111111;
assign micromatrizz[16][460] = 9'b111111111;
assign micromatrizz[16][461] = 9'b111111111;
assign micromatrizz[16][462] = 9'b111111111;
assign micromatrizz[16][463] = 9'b111111111;
assign micromatrizz[16][464] = 9'b111111111;
assign micromatrizz[16][465] = 9'b111111111;
assign micromatrizz[16][466] = 9'b111111111;
assign micromatrizz[16][467] = 9'b111111111;
assign micromatrizz[16][468] = 9'b111111111;
assign micromatrizz[16][469] = 9'b111111111;
assign micromatrizz[16][470] = 9'b111111111;
assign micromatrizz[16][471] = 9'b111111111;
assign micromatrizz[16][472] = 9'b111111111;
assign micromatrizz[16][473] = 9'b111111111;
assign micromatrizz[16][474] = 9'b111111111;
assign micromatrizz[16][475] = 9'b111111111;
assign micromatrizz[16][476] = 9'b111111111;
assign micromatrizz[16][477] = 9'b111111111;
assign micromatrizz[16][478] = 9'b111111111;
assign micromatrizz[16][479] = 9'b111111111;
assign micromatrizz[16][480] = 9'b111111111;
assign micromatrizz[16][481] = 9'b111111111;
assign micromatrizz[16][482] = 9'b111111111;
assign micromatrizz[16][483] = 9'b111111111;
assign micromatrizz[16][484] = 9'b111111111;
assign micromatrizz[16][485] = 9'b111111111;
assign micromatrizz[16][486] = 9'b111111111;
assign micromatrizz[16][487] = 9'b111111111;
assign micromatrizz[16][488] = 9'b111111111;
assign micromatrizz[16][489] = 9'b111111111;
assign micromatrizz[16][490] = 9'b111111111;
assign micromatrizz[16][491] = 9'b111111111;
assign micromatrizz[16][492] = 9'b111111111;
assign micromatrizz[16][493] = 9'b111111111;
assign micromatrizz[16][494] = 9'b111111111;
assign micromatrizz[16][495] = 9'b111111111;
assign micromatrizz[16][496] = 9'b111111111;
assign micromatrizz[16][497] = 9'b111111111;
assign micromatrizz[16][498] = 9'b111111111;
assign micromatrizz[16][499] = 9'b111111111;
assign micromatrizz[16][500] = 9'b111111111;
assign micromatrizz[16][501] = 9'b111111111;
assign micromatrizz[16][502] = 9'b111111111;
assign micromatrizz[16][503] = 9'b111111111;
assign micromatrizz[16][504] = 9'b111111111;
assign micromatrizz[16][505] = 9'b111111111;
assign micromatrizz[16][506] = 9'b111111111;
assign micromatrizz[16][507] = 9'b111111111;
assign micromatrizz[16][508] = 9'b111111111;
assign micromatrizz[16][509] = 9'b111111111;
assign micromatrizz[16][510] = 9'b111111111;
assign micromatrizz[16][511] = 9'b111111111;
assign micromatrizz[16][512] = 9'b111111111;
assign micromatrizz[16][513] = 9'b111111111;
assign micromatrizz[16][514] = 9'b111111111;
assign micromatrizz[16][515] = 9'b111111111;
assign micromatrizz[16][516] = 9'b111111111;
assign micromatrizz[16][517] = 9'b111111111;
assign micromatrizz[16][518] = 9'b111111111;
assign micromatrizz[16][519] = 9'b111111111;
assign micromatrizz[16][520] = 9'b111111111;
assign micromatrizz[16][521] = 9'b111111111;
assign micromatrizz[16][522] = 9'b111111111;
assign micromatrizz[16][523] = 9'b111111111;
assign micromatrizz[16][524] = 9'b111111111;
assign micromatrizz[16][525] = 9'b111111111;
assign micromatrizz[16][526] = 9'b111111111;
assign micromatrizz[16][527] = 9'b111111111;
assign micromatrizz[16][528] = 9'b111111111;
assign micromatrizz[16][529] = 9'b111111111;
assign micromatrizz[16][530] = 9'b111111111;
assign micromatrizz[16][531] = 9'b111111111;
assign micromatrizz[16][532] = 9'b111111111;
assign micromatrizz[16][533] = 9'b111111111;
assign micromatrizz[16][534] = 9'b111111111;
assign micromatrizz[16][535] = 9'b111111111;
assign micromatrizz[16][536] = 9'b111111111;
assign micromatrizz[16][537] = 9'b111111111;
assign micromatrizz[16][538] = 9'b111111111;
assign micromatrizz[16][539] = 9'b111111111;
assign micromatrizz[16][540] = 9'b111111111;
assign micromatrizz[16][541] = 9'b111111111;
assign micromatrizz[16][542] = 9'b111111111;
assign micromatrizz[16][543] = 9'b111111111;
assign micromatrizz[16][544] = 9'b111111111;
assign micromatrizz[16][545] = 9'b111111111;
assign micromatrizz[16][546] = 9'b111111111;
assign micromatrizz[16][547] = 9'b111111111;
assign micromatrizz[16][548] = 9'b111111111;
assign micromatrizz[16][549] = 9'b111111111;
assign micromatrizz[16][550] = 9'b111111111;
assign micromatrizz[16][551] = 9'b111111111;
assign micromatrizz[16][552] = 9'b111111111;
assign micromatrizz[16][553] = 9'b111111111;
assign micromatrizz[16][554] = 9'b111111111;
assign micromatrizz[16][555] = 9'b111111111;
assign micromatrizz[16][556] = 9'b111111111;
assign micromatrizz[16][557] = 9'b111111111;
assign micromatrizz[16][558] = 9'b111111111;
assign micromatrizz[16][559] = 9'b111111111;
assign micromatrizz[16][560] = 9'b111111111;
assign micromatrizz[16][561] = 9'b111111111;
assign micromatrizz[16][562] = 9'b111111111;
assign micromatrizz[16][563] = 9'b111111111;
assign micromatrizz[16][564] = 9'b111111111;
assign micromatrizz[16][565] = 9'b111111111;
assign micromatrizz[16][566] = 9'b111111111;
assign micromatrizz[16][567] = 9'b111111111;
assign micromatrizz[16][568] = 9'b111111111;
assign micromatrizz[16][569] = 9'b111111111;
assign micromatrizz[16][570] = 9'b111111111;
assign micromatrizz[16][571] = 9'b111111111;
assign micromatrizz[16][572] = 9'b111111111;
assign micromatrizz[16][573] = 9'b111111111;
assign micromatrizz[16][574] = 9'b111111111;
assign micromatrizz[16][575] = 9'b111111111;
assign micromatrizz[16][576] = 9'b111111111;
assign micromatrizz[16][577] = 9'b111111111;
assign micromatrizz[16][578] = 9'b111111111;
assign micromatrizz[16][579] = 9'b111111111;
assign micromatrizz[16][580] = 9'b111111111;
assign micromatrizz[16][581] = 9'b111111111;
assign micromatrizz[16][582] = 9'b111111111;
assign micromatrizz[16][583] = 9'b111111111;
assign micromatrizz[16][584] = 9'b111111111;
assign micromatrizz[16][585] = 9'b111111111;
assign micromatrizz[16][586] = 9'b111111111;
assign micromatrizz[16][587] = 9'b111111111;
assign micromatrizz[16][588] = 9'b111111111;
assign micromatrizz[16][589] = 9'b111111111;
assign micromatrizz[16][590] = 9'b111111111;
assign micromatrizz[16][591] = 9'b111111111;
assign micromatrizz[16][592] = 9'b111111111;
assign micromatrizz[16][593] = 9'b111111111;
assign micromatrizz[16][594] = 9'b111111111;
assign micromatrizz[16][595] = 9'b111111111;
assign micromatrizz[16][596] = 9'b111111111;
assign micromatrizz[16][597] = 9'b111111111;
assign micromatrizz[16][598] = 9'b111111111;
assign micromatrizz[16][599] = 9'b111111111;
assign micromatrizz[16][600] = 9'b111111111;
assign micromatrizz[16][601] = 9'b111111111;
assign micromatrizz[16][602] = 9'b111111111;
assign micromatrizz[16][603] = 9'b111111111;
assign micromatrizz[16][604] = 9'b111111111;
assign micromatrizz[16][605] = 9'b111111111;
assign micromatrizz[16][606] = 9'b111111111;
assign micromatrizz[16][607] = 9'b111111111;
assign micromatrizz[16][608] = 9'b111111111;
assign micromatrizz[16][609] = 9'b111111111;
assign micromatrizz[16][610] = 9'b111111111;
assign micromatrizz[16][611] = 9'b111111111;
assign micromatrizz[16][612] = 9'b111111111;
assign micromatrizz[16][613] = 9'b111111111;
assign micromatrizz[16][614] = 9'b111111111;
assign micromatrizz[16][615] = 9'b111111111;
assign micromatrizz[16][616] = 9'b111111111;
assign micromatrizz[16][617] = 9'b111111111;
assign micromatrizz[16][618] = 9'b111111111;
assign micromatrizz[16][619] = 9'b111111111;
assign micromatrizz[16][620] = 9'b111111111;
assign micromatrizz[16][621] = 9'b111111111;
assign micromatrizz[16][622] = 9'b111111111;
assign micromatrizz[16][623] = 9'b111111111;
assign micromatrizz[16][624] = 9'b111111111;
assign micromatrizz[16][625] = 9'b111111111;
assign micromatrizz[16][626] = 9'b111111111;
assign micromatrizz[16][627] = 9'b111111111;
assign micromatrizz[16][628] = 9'b111111111;
assign micromatrizz[16][629] = 9'b111111111;
assign micromatrizz[16][630] = 9'b111111111;
assign micromatrizz[16][631] = 9'b111111111;
assign micromatrizz[16][632] = 9'b111111111;
assign micromatrizz[16][633] = 9'b111111111;
assign micromatrizz[16][634] = 9'b111111111;
assign micromatrizz[16][635] = 9'b111111111;
assign micromatrizz[16][636] = 9'b111111111;
assign micromatrizz[16][637] = 9'b111111111;
assign micromatrizz[16][638] = 9'b111111111;
assign micromatrizz[16][639] = 9'b111111111;
assign micromatrizz[17][0] = 9'b111111111;
assign micromatrizz[17][1] = 9'b111111111;
assign micromatrizz[17][2] = 9'b111111111;
assign micromatrizz[17][3] = 9'b111111111;
assign micromatrizz[17][4] = 9'b111111111;
assign micromatrizz[17][5] = 9'b111111111;
assign micromatrizz[17][6] = 9'b111111111;
assign micromatrizz[17][7] = 9'b111111111;
assign micromatrizz[17][8] = 9'b111111111;
assign micromatrizz[17][9] = 9'b111111111;
assign micromatrizz[17][10] = 9'b111111111;
assign micromatrizz[17][11] = 9'b111111111;
assign micromatrizz[17][12] = 9'b111111111;
assign micromatrizz[17][13] = 9'b111111111;
assign micromatrizz[17][14] = 9'b111111111;
assign micromatrizz[17][15] = 9'b111111111;
assign micromatrizz[17][16] = 9'b111111111;
assign micromatrizz[17][17] = 9'b111111111;
assign micromatrizz[17][18] = 9'b111111111;
assign micromatrizz[17][19] = 9'b111111111;
assign micromatrizz[17][20] = 9'b111111111;
assign micromatrizz[17][21] = 9'b111111111;
assign micromatrizz[17][22] = 9'b111111111;
assign micromatrizz[17][23] = 9'b111111111;
assign micromatrizz[17][24] = 9'b111111111;
assign micromatrizz[17][25] = 9'b111111111;
assign micromatrizz[17][26] = 9'b111111111;
assign micromatrizz[17][27] = 9'b111111111;
assign micromatrizz[17][28] = 9'b111111111;
assign micromatrizz[17][29] = 9'b111111111;
assign micromatrizz[17][30] = 9'b111111111;
assign micromatrizz[17][31] = 9'b111111111;
assign micromatrizz[17][32] = 9'b111111111;
assign micromatrizz[17][33] = 9'b111111111;
assign micromatrizz[17][34] = 9'b111111111;
assign micromatrizz[17][35] = 9'b111111111;
assign micromatrizz[17][36] = 9'b111111111;
assign micromatrizz[17][37] = 9'b111111111;
assign micromatrizz[17][38] = 9'b111111111;
assign micromatrizz[17][39] = 9'b111111111;
assign micromatrizz[17][40] = 9'b111111111;
assign micromatrizz[17][41] = 9'b111111111;
assign micromatrizz[17][42] = 9'b111111111;
assign micromatrizz[17][43] = 9'b111111111;
assign micromatrizz[17][44] = 9'b111111111;
assign micromatrizz[17][45] = 9'b111111111;
assign micromatrizz[17][46] = 9'b111111111;
assign micromatrizz[17][47] = 9'b111111111;
assign micromatrizz[17][48] = 9'b111111111;
assign micromatrizz[17][49] = 9'b111111111;
assign micromatrizz[17][50] = 9'b111111111;
assign micromatrizz[17][51] = 9'b111111111;
assign micromatrizz[17][52] = 9'b111111111;
assign micromatrizz[17][53] = 9'b111111111;
assign micromatrizz[17][54] = 9'b111111111;
assign micromatrizz[17][55] = 9'b111111111;
assign micromatrizz[17][56] = 9'b111111111;
assign micromatrizz[17][57] = 9'b111111111;
assign micromatrizz[17][58] = 9'b111111111;
assign micromatrizz[17][59] = 9'b111111111;
assign micromatrizz[17][60] = 9'b111111111;
assign micromatrizz[17][61] = 9'b111111111;
assign micromatrizz[17][62] = 9'b111111111;
assign micromatrizz[17][63] = 9'b111111111;
assign micromatrizz[17][64] = 9'b111111111;
assign micromatrizz[17][65] = 9'b111111111;
assign micromatrizz[17][66] = 9'b111111111;
assign micromatrizz[17][67] = 9'b111111111;
assign micromatrizz[17][68] = 9'b111111111;
assign micromatrizz[17][69] = 9'b111111111;
assign micromatrizz[17][70] = 9'b111111111;
assign micromatrizz[17][71] = 9'b111111111;
assign micromatrizz[17][72] = 9'b111111111;
assign micromatrizz[17][73] = 9'b111111111;
assign micromatrizz[17][74] = 9'b111111111;
assign micromatrizz[17][75] = 9'b111111111;
assign micromatrizz[17][76] = 9'b111111111;
assign micromatrizz[17][77] = 9'b111111111;
assign micromatrizz[17][78] = 9'b111111111;
assign micromatrizz[17][79] = 9'b111111111;
assign micromatrizz[17][80] = 9'b111111111;
assign micromatrizz[17][81] = 9'b111111111;
assign micromatrizz[17][82] = 9'b111111111;
assign micromatrizz[17][83] = 9'b111111111;
assign micromatrizz[17][84] = 9'b111111111;
assign micromatrizz[17][85] = 9'b111111111;
assign micromatrizz[17][86] = 9'b111111111;
assign micromatrizz[17][87] = 9'b111111111;
assign micromatrizz[17][88] = 9'b111111111;
assign micromatrizz[17][89] = 9'b111111111;
assign micromatrizz[17][90] = 9'b111111111;
assign micromatrizz[17][91] = 9'b111111111;
assign micromatrizz[17][92] = 9'b111111111;
assign micromatrizz[17][93] = 9'b111111111;
assign micromatrizz[17][94] = 9'b111111111;
assign micromatrizz[17][95] = 9'b111111111;
assign micromatrizz[17][96] = 9'b111111111;
assign micromatrizz[17][97] = 9'b111111111;
assign micromatrizz[17][98] = 9'b111111111;
assign micromatrizz[17][99] = 9'b111111111;
assign micromatrizz[17][100] = 9'b111111111;
assign micromatrizz[17][101] = 9'b111111111;
assign micromatrizz[17][102] = 9'b111111111;
assign micromatrizz[17][103] = 9'b111111111;
assign micromatrizz[17][104] = 9'b111111111;
assign micromatrizz[17][105] = 9'b111111111;
assign micromatrizz[17][106] = 9'b111111111;
assign micromatrizz[17][107] = 9'b111111111;
assign micromatrizz[17][108] = 9'b111111111;
assign micromatrizz[17][109] = 9'b111111111;
assign micromatrizz[17][110] = 9'b111111111;
assign micromatrizz[17][111] = 9'b111111111;
assign micromatrizz[17][112] = 9'b111111111;
assign micromatrizz[17][113] = 9'b111111111;
assign micromatrizz[17][114] = 9'b111111111;
assign micromatrizz[17][115] = 9'b111111111;
assign micromatrizz[17][116] = 9'b111111111;
assign micromatrizz[17][117] = 9'b111111111;
assign micromatrizz[17][118] = 9'b111111111;
assign micromatrizz[17][119] = 9'b111111111;
assign micromatrizz[17][120] = 9'b111111111;
assign micromatrizz[17][121] = 9'b111111111;
assign micromatrizz[17][122] = 9'b111111111;
assign micromatrizz[17][123] = 9'b111111111;
assign micromatrizz[17][124] = 9'b111111111;
assign micromatrizz[17][125] = 9'b111111111;
assign micromatrizz[17][126] = 9'b111111111;
assign micromatrizz[17][127] = 9'b111111111;
assign micromatrizz[17][128] = 9'b111111111;
assign micromatrizz[17][129] = 9'b111111111;
assign micromatrizz[17][130] = 9'b111111111;
assign micromatrizz[17][131] = 9'b111111111;
assign micromatrizz[17][132] = 9'b111111111;
assign micromatrizz[17][133] = 9'b111111111;
assign micromatrizz[17][134] = 9'b111111111;
assign micromatrizz[17][135] = 9'b111111111;
assign micromatrizz[17][136] = 9'b111111111;
assign micromatrizz[17][137] = 9'b111111111;
assign micromatrizz[17][138] = 9'b111111111;
assign micromatrizz[17][139] = 9'b111111111;
assign micromatrizz[17][140] = 9'b111111111;
assign micromatrizz[17][141] = 9'b111111111;
assign micromatrizz[17][142] = 9'b111111111;
assign micromatrizz[17][143] = 9'b111111111;
assign micromatrizz[17][144] = 9'b111111111;
assign micromatrizz[17][145] = 9'b111111111;
assign micromatrizz[17][146] = 9'b111111111;
assign micromatrizz[17][147] = 9'b111111111;
assign micromatrizz[17][148] = 9'b111111111;
assign micromatrizz[17][149] = 9'b111111111;
assign micromatrizz[17][150] = 9'b111111111;
assign micromatrizz[17][151] = 9'b111111111;
assign micromatrizz[17][152] = 9'b111111111;
assign micromatrizz[17][153] = 9'b111111111;
assign micromatrizz[17][154] = 9'b111111111;
assign micromatrizz[17][155] = 9'b111111111;
assign micromatrizz[17][156] = 9'b111111111;
assign micromatrizz[17][157] = 9'b111111111;
assign micromatrizz[17][158] = 9'b111111111;
assign micromatrizz[17][159] = 9'b111111111;
assign micromatrizz[17][160] = 9'b111111111;
assign micromatrizz[17][161] = 9'b111111111;
assign micromatrizz[17][162] = 9'b111111111;
assign micromatrizz[17][163] = 9'b111111111;
assign micromatrizz[17][164] = 9'b111111111;
assign micromatrizz[17][165] = 9'b111111111;
assign micromatrizz[17][166] = 9'b111111111;
assign micromatrizz[17][167] = 9'b111111111;
assign micromatrizz[17][168] = 9'b111111111;
assign micromatrizz[17][169] = 9'b111111111;
assign micromatrizz[17][170] = 9'b111111111;
assign micromatrizz[17][171] = 9'b111111111;
assign micromatrizz[17][172] = 9'b111111111;
assign micromatrizz[17][173] = 9'b111111111;
assign micromatrizz[17][174] = 9'b111111111;
assign micromatrizz[17][175] = 9'b111111111;
assign micromatrizz[17][176] = 9'b111111111;
assign micromatrizz[17][177] = 9'b111111111;
assign micromatrizz[17][178] = 9'b111111111;
assign micromatrizz[17][179] = 9'b111111111;
assign micromatrizz[17][180] = 9'b111111111;
assign micromatrizz[17][181] = 9'b111111111;
assign micromatrizz[17][182] = 9'b111111111;
assign micromatrizz[17][183] = 9'b111111111;
assign micromatrizz[17][184] = 9'b111111111;
assign micromatrizz[17][185] = 9'b111111111;
assign micromatrizz[17][186] = 9'b111111111;
assign micromatrizz[17][187] = 9'b111111111;
assign micromatrizz[17][188] = 9'b111111111;
assign micromatrizz[17][189] = 9'b111111111;
assign micromatrizz[17][190] = 9'b111111111;
assign micromatrizz[17][191] = 9'b111111111;
assign micromatrizz[17][192] = 9'b111111111;
assign micromatrizz[17][193] = 9'b111111111;
assign micromatrizz[17][194] = 9'b111111111;
assign micromatrizz[17][195] = 9'b111111111;
assign micromatrizz[17][196] = 9'b111111111;
assign micromatrizz[17][197] = 9'b111111111;
assign micromatrizz[17][198] = 9'b111111111;
assign micromatrizz[17][199] = 9'b111111111;
assign micromatrizz[17][200] = 9'b111111111;
assign micromatrizz[17][201] = 9'b111111111;
assign micromatrizz[17][202] = 9'b111111111;
assign micromatrizz[17][203] = 9'b111111111;
assign micromatrizz[17][204] = 9'b111111111;
assign micromatrizz[17][205] = 9'b111111111;
assign micromatrizz[17][206] = 9'b111111111;
assign micromatrizz[17][207] = 9'b111111111;
assign micromatrizz[17][208] = 9'b111111111;
assign micromatrizz[17][209] = 9'b111111111;
assign micromatrizz[17][210] = 9'b111111111;
assign micromatrizz[17][211] = 9'b111111111;
assign micromatrizz[17][212] = 9'b111111111;
assign micromatrizz[17][213] = 9'b111111111;
assign micromatrizz[17][214] = 9'b111111111;
assign micromatrizz[17][215] = 9'b111111111;
assign micromatrizz[17][216] = 9'b111111111;
assign micromatrizz[17][217] = 9'b111111111;
assign micromatrizz[17][218] = 9'b111111111;
assign micromatrizz[17][219] = 9'b111111111;
assign micromatrizz[17][220] = 9'b111111111;
assign micromatrizz[17][221] = 9'b111111111;
assign micromatrizz[17][222] = 9'b111111111;
assign micromatrizz[17][223] = 9'b111111111;
assign micromatrizz[17][224] = 9'b111111111;
assign micromatrizz[17][225] = 9'b111111111;
assign micromatrizz[17][226] = 9'b111111111;
assign micromatrizz[17][227] = 9'b111111111;
assign micromatrizz[17][228] = 9'b111111111;
assign micromatrizz[17][229] = 9'b111111111;
assign micromatrizz[17][230] = 9'b111111111;
assign micromatrizz[17][231] = 9'b111111111;
assign micromatrizz[17][232] = 9'b111111111;
assign micromatrizz[17][233] = 9'b111111111;
assign micromatrizz[17][234] = 9'b111111111;
assign micromatrizz[17][235] = 9'b111111111;
assign micromatrizz[17][236] = 9'b111111111;
assign micromatrizz[17][237] = 9'b111111111;
assign micromatrizz[17][238] = 9'b111111111;
assign micromatrizz[17][239] = 9'b111111111;
assign micromatrizz[17][240] = 9'b111111111;
assign micromatrizz[17][241] = 9'b111111111;
assign micromatrizz[17][242] = 9'b111111111;
assign micromatrizz[17][243] = 9'b111111111;
assign micromatrizz[17][244] = 9'b111111111;
assign micromatrizz[17][245] = 9'b111111111;
assign micromatrizz[17][246] = 9'b111111111;
assign micromatrizz[17][247] = 9'b111111111;
assign micromatrizz[17][248] = 9'b111111111;
assign micromatrizz[17][249] = 9'b111111111;
assign micromatrizz[17][250] = 9'b111111111;
assign micromatrizz[17][251] = 9'b111111111;
assign micromatrizz[17][252] = 9'b111111111;
assign micromatrizz[17][253] = 9'b111111111;
assign micromatrizz[17][254] = 9'b111111111;
assign micromatrizz[17][255] = 9'b111111111;
assign micromatrizz[17][256] = 9'b111111111;
assign micromatrizz[17][257] = 9'b111111111;
assign micromatrizz[17][258] = 9'b111111111;
assign micromatrizz[17][259] = 9'b111111111;
assign micromatrizz[17][260] = 9'b111111111;
assign micromatrizz[17][261] = 9'b111111111;
assign micromatrizz[17][262] = 9'b111111111;
assign micromatrizz[17][263] = 9'b111111111;
assign micromatrizz[17][264] = 9'b111111111;
assign micromatrizz[17][265] = 9'b111111111;
assign micromatrizz[17][266] = 9'b111111111;
assign micromatrizz[17][267] = 9'b111111111;
assign micromatrizz[17][268] = 9'b111111111;
assign micromatrizz[17][269] = 9'b111111111;
assign micromatrizz[17][270] = 9'b111111111;
assign micromatrizz[17][271] = 9'b111111111;
assign micromatrizz[17][272] = 9'b111111111;
assign micromatrizz[17][273] = 9'b111111111;
assign micromatrizz[17][274] = 9'b111111111;
assign micromatrizz[17][275] = 9'b111111111;
assign micromatrizz[17][276] = 9'b111111111;
assign micromatrizz[17][277] = 9'b111111111;
assign micromatrizz[17][278] = 9'b111111111;
assign micromatrizz[17][279] = 9'b111111111;
assign micromatrizz[17][280] = 9'b111111111;
assign micromatrizz[17][281] = 9'b111111111;
assign micromatrizz[17][282] = 9'b111111111;
assign micromatrizz[17][283] = 9'b111111111;
assign micromatrizz[17][284] = 9'b111111111;
assign micromatrizz[17][285] = 9'b111111111;
assign micromatrizz[17][286] = 9'b111111111;
assign micromatrizz[17][287] = 9'b111111111;
assign micromatrizz[17][288] = 9'b111111111;
assign micromatrizz[17][289] = 9'b111111111;
assign micromatrizz[17][290] = 9'b111111111;
assign micromatrizz[17][291] = 9'b111111111;
assign micromatrizz[17][292] = 9'b111111111;
assign micromatrizz[17][293] = 9'b111111111;
assign micromatrizz[17][294] = 9'b111111111;
assign micromatrizz[17][295] = 9'b111111111;
assign micromatrizz[17][296] = 9'b111111111;
assign micromatrizz[17][297] = 9'b111111111;
assign micromatrizz[17][298] = 9'b111111111;
assign micromatrizz[17][299] = 9'b111111111;
assign micromatrizz[17][300] = 9'b111111111;
assign micromatrizz[17][301] = 9'b111111111;
assign micromatrizz[17][302] = 9'b111111111;
assign micromatrizz[17][303] = 9'b111111111;
assign micromatrizz[17][304] = 9'b111111111;
assign micromatrizz[17][305] = 9'b111111111;
assign micromatrizz[17][306] = 9'b111111111;
assign micromatrizz[17][307] = 9'b111111111;
assign micromatrizz[17][308] = 9'b111111111;
assign micromatrizz[17][309] = 9'b111111111;
assign micromatrizz[17][310] = 9'b111111111;
assign micromatrizz[17][311] = 9'b111111111;
assign micromatrizz[17][312] = 9'b111111111;
assign micromatrizz[17][313] = 9'b111111111;
assign micromatrizz[17][314] = 9'b111111111;
assign micromatrizz[17][315] = 9'b111111111;
assign micromatrizz[17][316] = 9'b111111111;
assign micromatrizz[17][317] = 9'b111111111;
assign micromatrizz[17][318] = 9'b111111111;
assign micromatrizz[17][319] = 9'b111111111;
assign micromatrizz[17][320] = 9'b111111111;
assign micromatrizz[17][321] = 9'b111111111;
assign micromatrizz[17][322] = 9'b111111111;
assign micromatrizz[17][323] = 9'b111111111;
assign micromatrizz[17][324] = 9'b111111111;
assign micromatrizz[17][325] = 9'b111111111;
assign micromatrizz[17][326] = 9'b111111111;
assign micromatrizz[17][327] = 9'b111111111;
assign micromatrizz[17][328] = 9'b111111111;
assign micromatrizz[17][329] = 9'b111111111;
assign micromatrizz[17][330] = 9'b111111111;
assign micromatrizz[17][331] = 9'b111111111;
assign micromatrizz[17][332] = 9'b111111111;
assign micromatrizz[17][333] = 9'b111111111;
assign micromatrizz[17][334] = 9'b111111111;
assign micromatrizz[17][335] = 9'b111111111;
assign micromatrizz[17][336] = 9'b111111111;
assign micromatrizz[17][337] = 9'b111111111;
assign micromatrizz[17][338] = 9'b111111111;
assign micromatrizz[17][339] = 9'b111111111;
assign micromatrizz[17][340] = 9'b111111111;
assign micromatrizz[17][341] = 9'b111111111;
assign micromatrizz[17][342] = 9'b111111111;
assign micromatrizz[17][343] = 9'b111111111;
assign micromatrizz[17][344] = 9'b111111111;
assign micromatrizz[17][345] = 9'b111111111;
assign micromatrizz[17][346] = 9'b111111111;
assign micromatrizz[17][347] = 9'b111111111;
assign micromatrizz[17][348] = 9'b111111111;
assign micromatrizz[17][349] = 9'b111111111;
assign micromatrizz[17][350] = 9'b111111111;
assign micromatrizz[17][351] = 9'b111111111;
assign micromatrizz[17][352] = 9'b111111111;
assign micromatrizz[17][353] = 9'b111111111;
assign micromatrizz[17][354] = 9'b111111111;
assign micromatrizz[17][355] = 9'b111111111;
assign micromatrizz[17][356] = 9'b111111111;
assign micromatrizz[17][357] = 9'b111111111;
assign micromatrizz[17][358] = 9'b111111111;
assign micromatrizz[17][359] = 9'b111111111;
assign micromatrizz[17][360] = 9'b111111111;
assign micromatrizz[17][361] = 9'b111111111;
assign micromatrizz[17][362] = 9'b111111111;
assign micromatrizz[17][363] = 9'b111111111;
assign micromatrizz[17][364] = 9'b111111111;
assign micromatrizz[17][365] = 9'b111111111;
assign micromatrizz[17][366] = 9'b111111111;
assign micromatrizz[17][367] = 9'b111111111;
assign micromatrizz[17][368] = 9'b111111111;
assign micromatrizz[17][369] = 9'b111111111;
assign micromatrizz[17][370] = 9'b111111111;
assign micromatrizz[17][371] = 9'b111111111;
assign micromatrizz[17][372] = 9'b111111111;
assign micromatrizz[17][373] = 9'b111111111;
assign micromatrizz[17][374] = 9'b111111111;
assign micromatrizz[17][375] = 9'b111111111;
assign micromatrizz[17][376] = 9'b111111111;
assign micromatrizz[17][377] = 9'b111111111;
assign micromatrizz[17][378] = 9'b111111111;
assign micromatrizz[17][379] = 9'b111111111;
assign micromatrizz[17][380] = 9'b111111111;
assign micromatrizz[17][381] = 9'b111111111;
assign micromatrizz[17][382] = 9'b111111111;
assign micromatrizz[17][383] = 9'b111111111;
assign micromatrizz[17][384] = 9'b111111111;
assign micromatrizz[17][385] = 9'b111111111;
assign micromatrizz[17][386] = 9'b111111111;
assign micromatrizz[17][387] = 9'b111111111;
assign micromatrizz[17][388] = 9'b111111111;
assign micromatrizz[17][389] = 9'b111111111;
assign micromatrizz[17][390] = 9'b111111111;
assign micromatrizz[17][391] = 9'b111111111;
assign micromatrizz[17][392] = 9'b111111111;
assign micromatrizz[17][393] = 9'b111111111;
assign micromatrizz[17][394] = 9'b111111111;
assign micromatrizz[17][395] = 9'b111111111;
assign micromatrizz[17][396] = 9'b111111111;
assign micromatrizz[17][397] = 9'b111111111;
assign micromatrizz[17][398] = 9'b111111111;
assign micromatrizz[17][399] = 9'b111111111;
assign micromatrizz[17][400] = 9'b111111111;
assign micromatrizz[17][401] = 9'b111111111;
assign micromatrizz[17][402] = 9'b111111111;
assign micromatrizz[17][403] = 9'b111111111;
assign micromatrizz[17][404] = 9'b111111111;
assign micromatrizz[17][405] = 9'b111111111;
assign micromatrizz[17][406] = 9'b111111111;
assign micromatrizz[17][407] = 9'b111111111;
assign micromatrizz[17][408] = 9'b111111111;
assign micromatrizz[17][409] = 9'b111111111;
assign micromatrizz[17][410] = 9'b111111111;
assign micromatrizz[17][411] = 9'b111111111;
assign micromatrizz[17][412] = 9'b111111111;
assign micromatrizz[17][413] = 9'b111111111;
assign micromatrizz[17][414] = 9'b111111111;
assign micromatrizz[17][415] = 9'b111111111;
assign micromatrizz[17][416] = 9'b111111111;
assign micromatrizz[17][417] = 9'b111111111;
assign micromatrizz[17][418] = 9'b111111111;
assign micromatrizz[17][419] = 9'b111111111;
assign micromatrizz[17][420] = 9'b111111111;
assign micromatrizz[17][421] = 9'b111111111;
assign micromatrizz[17][422] = 9'b111111111;
assign micromatrizz[17][423] = 9'b111111111;
assign micromatrizz[17][424] = 9'b111111111;
assign micromatrizz[17][425] = 9'b111111111;
assign micromatrizz[17][426] = 9'b111111111;
assign micromatrizz[17][427] = 9'b111111111;
assign micromatrizz[17][428] = 9'b111111111;
assign micromatrizz[17][429] = 9'b111111111;
assign micromatrizz[17][430] = 9'b111111111;
assign micromatrizz[17][431] = 9'b111111111;
assign micromatrizz[17][432] = 9'b111111111;
assign micromatrizz[17][433] = 9'b111111111;
assign micromatrizz[17][434] = 9'b111111111;
assign micromatrizz[17][435] = 9'b111111111;
assign micromatrizz[17][436] = 9'b111111111;
assign micromatrizz[17][437] = 9'b111111111;
assign micromatrizz[17][438] = 9'b111111111;
assign micromatrizz[17][439] = 9'b111111111;
assign micromatrizz[17][440] = 9'b111111111;
assign micromatrizz[17][441] = 9'b111111111;
assign micromatrizz[17][442] = 9'b111111111;
assign micromatrizz[17][443] = 9'b111111111;
assign micromatrizz[17][444] = 9'b111111111;
assign micromatrizz[17][445] = 9'b111111111;
assign micromatrizz[17][446] = 9'b111111111;
assign micromatrizz[17][447] = 9'b111111111;
assign micromatrizz[17][448] = 9'b111111111;
assign micromatrizz[17][449] = 9'b111111111;
assign micromatrizz[17][450] = 9'b111111111;
assign micromatrizz[17][451] = 9'b111111111;
assign micromatrizz[17][452] = 9'b111111111;
assign micromatrizz[17][453] = 9'b111111111;
assign micromatrizz[17][454] = 9'b111111111;
assign micromatrizz[17][455] = 9'b111111111;
assign micromatrizz[17][456] = 9'b111111111;
assign micromatrizz[17][457] = 9'b111111111;
assign micromatrizz[17][458] = 9'b111111111;
assign micromatrizz[17][459] = 9'b111111111;
assign micromatrizz[17][460] = 9'b111111111;
assign micromatrizz[17][461] = 9'b111111111;
assign micromatrizz[17][462] = 9'b111111111;
assign micromatrizz[17][463] = 9'b111111111;
assign micromatrizz[17][464] = 9'b111111111;
assign micromatrizz[17][465] = 9'b111111111;
assign micromatrizz[17][466] = 9'b111111111;
assign micromatrizz[17][467] = 9'b111111111;
assign micromatrizz[17][468] = 9'b111111111;
assign micromatrizz[17][469] = 9'b111111111;
assign micromatrizz[17][470] = 9'b111111111;
assign micromatrizz[17][471] = 9'b111111111;
assign micromatrizz[17][472] = 9'b111111111;
assign micromatrizz[17][473] = 9'b111111111;
assign micromatrizz[17][474] = 9'b111111111;
assign micromatrizz[17][475] = 9'b111111111;
assign micromatrizz[17][476] = 9'b111111111;
assign micromatrizz[17][477] = 9'b111111111;
assign micromatrizz[17][478] = 9'b111111111;
assign micromatrizz[17][479] = 9'b111111111;
assign micromatrizz[17][480] = 9'b111111111;
assign micromatrizz[17][481] = 9'b111111111;
assign micromatrizz[17][482] = 9'b111111111;
assign micromatrizz[17][483] = 9'b111111111;
assign micromatrizz[17][484] = 9'b111111111;
assign micromatrizz[17][485] = 9'b111111111;
assign micromatrizz[17][486] = 9'b111111111;
assign micromatrizz[17][487] = 9'b111111111;
assign micromatrizz[17][488] = 9'b111111111;
assign micromatrizz[17][489] = 9'b111111111;
assign micromatrizz[17][490] = 9'b111111111;
assign micromatrizz[17][491] = 9'b111111111;
assign micromatrizz[17][492] = 9'b111111111;
assign micromatrizz[17][493] = 9'b111111111;
assign micromatrizz[17][494] = 9'b111111111;
assign micromatrizz[17][495] = 9'b111111111;
assign micromatrizz[17][496] = 9'b111111111;
assign micromatrizz[17][497] = 9'b111111111;
assign micromatrizz[17][498] = 9'b111111111;
assign micromatrizz[17][499] = 9'b111111111;
assign micromatrizz[17][500] = 9'b111111111;
assign micromatrizz[17][501] = 9'b111111111;
assign micromatrizz[17][502] = 9'b111111111;
assign micromatrizz[17][503] = 9'b111111111;
assign micromatrizz[17][504] = 9'b111111111;
assign micromatrizz[17][505] = 9'b111111111;
assign micromatrizz[17][506] = 9'b111111111;
assign micromatrizz[17][507] = 9'b111111111;
assign micromatrizz[17][508] = 9'b111111111;
assign micromatrizz[17][509] = 9'b111111111;
assign micromatrizz[17][510] = 9'b111111111;
assign micromatrizz[17][511] = 9'b111111111;
assign micromatrizz[17][512] = 9'b111111111;
assign micromatrizz[17][513] = 9'b111111111;
assign micromatrizz[17][514] = 9'b111111111;
assign micromatrizz[17][515] = 9'b111111111;
assign micromatrizz[17][516] = 9'b111111111;
assign micromatrizz[17][517] = 9'b111111111;
assign micromatrizz[17][518] = 9'b111111111;
assign micromatrizz[17][519] = 9'b111111111;
assign micromatrizz[17][520] = 9'b111111111;
assign micromatrizz[17][521] = 9'b111111111;
assign micromatrizz[17][522] = 9'b111111111;
assign micromatrizz[17][523] = 9'b111111111;
assign micromatrizz[17][524] = 9'b111111111;
assign micromatrizz[17][525] = 9'b111111111;
assign micromatrizz[17][526] = 9'b111111111;
assign micromatrizz[17][527] = 9'b111111111;
assign micromatrizz[17][528] = 9'b111111111;
assign micromatrizz[17][529] = 9'b111111111;
assign micromatrizz[17][530] = 9'b111111111;
assign micromatrizz[17][531] = 9'b111111111;
assign micromatrizz[17][532] = 9'b111111111;
assign micromatrizz[17][533] = 9'b111111111;
assign micromatrizz[17][534] = 9'b111111111;
assign micromatrizz[17][535] = 9'b111111111;
assign micromatrizz[17][536] = 9'b111111111;
assign micromatrizz[17][537] = 9'b111111111;
assign micromatrizz[17][538] = 9'b111111111;
assign micromatrizz[17][539] = 9'b111111111;
assign micromatrizz[17][540] = 9'b111111111;
assign micromatrizz[17][541] = 9'b111111111;
assign micromatrizz[17][542] = 9'b111111111;
assign micromatrizz[17][543] = 9'b111111111;
assign micromatrizz[17][544] = 9'b111111111;
assign micromatrizz[17][545] = 9'b111111111;
assign micromatrizz[17][546] = 9'b111111111;
assign micromatrizz[17][547] = 9'b111111111;
assign micromatrizz[17][548] = 9'b111111111;
assign micromatrizz[17][549] = 9'b111111111;
assign micromatrizz[17][550] = 9'b111111111;
assign micromatrizz[17][551] = 9'b111111111;
assign micromatrizz[17][552] = 9'b111111111;
assign micromatrizz[17][553] = 9'b111111111;
assign micromatrizz[17][554] = 9'b111111111;
assign micromatrizz[17][555] = 9'b111111111;
assign micromatrizz[17][556] = 9'b111111111;
assign micromatrizz[17][557] = 9'b111111111;
assign micromatrizz[17][558] = 9'b111111111;
assign micromatrizz[17][559] = 9'b111111111;
assign micromatrizz[17][560] = 9'b111111111;
assign micromatrizz[17][561] = 9'b111111111;
assign micromatrizz[17][562] = 9'b111111111;
assign micromatrizz[17][563] = 9'b111111111;
assign micromatrizz[17][564] = 9'b111111111;
assign micromatrizz[17][565] = 9'b111111111;
assign micromatrizz[17][566] = 9'b111111111;
assign micromatrizz[17][567] = 9'b111111111;
assign micromatrizz[17][568] = 9'b111111111;
assign micromatrizz[17][569] = 9'b111111111;
assign micromatrizz[17][570] = 9'b111111111;
assign micromatrizz[17][571] = 9'b111111111;
assign micromatrizz[17][572] = 9'b111111111;
assign micromatrizz[17][573] = 9'b111111111;
assign micromatrizz[17][574] = 9'b111111111;
assign micromatrizz[17][575] = 9'b111111111;
assign micromatrizz[17][576] = 9'b111111111;
assign micromatrizz[17][577] = 9'b111111111;
assign micromatrizz[17][578] = 9'b111111111;
assign micromatrizz[17][579] = 9'b111111111;
assign micromatrizz[17][580] = 9'b111111111;
assign micromatrizz[17][581] = 9'b111111111;
assign micromatrizz[17][582] = 9'b111111111;
assign micromatrizz[17][583] = 9'b111111111;
assign micromatrizz[17][584] = 9'b111111111;
assign micromatrizz[17][585] = 9'b111111111;
assign micromatrizz[17][586] = 9'b111111111;
assign micromatrizz[17][587] = 9'b111111111;
assign micromatrizz[17][588] = 9'b111111111;
assign micromatrizz[17][589] = 9'b111111111;
assign micromatrizz[17][590] = 9'b111111111;
assign micromatrizz[17][591] = 9'b111111111;
assign micromatrizz[17][592] = 9'b111111111;
assign micromatrizz[17][593] = 9'b111111111;
assign micromatrizz[17][594] = 9'b111111111;
assign micromatrizz[17][595] = 9'b111111111;
assign micromatrizz[17][596] = 9'b111111111;
assign micromatrizz[17][597] = 9'b111111111;
assign micromatrizz[17][598] = 9'b111111111;
assign micromatrizz[17][599] = 9'b111111111;
assign micromatrizz[17][600] = 9'b111111111;
assign micromatrizz[17][601] = 9'b111111111;
assign micromatrizz[17][602] = 9'b111111111;
assign micromatrizz[17][603] = 9'b111111111;
assign micromatrizz[17][604] = 9'b111111111;
assign micromatrizz[17][605] = 9'b111111111;
assign micromatrizz[17][606] = 9'b111111111;
assign micromatrizz[17][607] = 9'b111111111;
assign micromatrizz[17][608] = 9'b111111111;
assign micromatrizz[17][609] = 9'b111111111;
assign micromatrizz[17][610] = 9'b111111111;
assign micromatrizz[17][611] = 9'b111111111;
assign micromatrizz[17][612] = 9'b111111111;
assign micromatrizz[17][613] = 9'b111111111;
assign micromatrizz[17][614] = 9'b111111111;
assign micromatrizz[17][615] = 9'b111111111;
assign micromatrizz[17][616] = 9'b111111111;
assign micromatrizz[17][617] = 9'b111111111;
assign micromatrizz[17][618] = 9'b111111111;
assign micromatrizz[17][619] = 9'b111111111;
assign micromatrizz[17][620] = 9'b111111111;
assign micromatrizz[17][621] = 9'b111111111;
assign micromatrizz[17][622] = 9'b111111111;
assign micromatrizz[17][623] = 9'b111111111;
assign micromatrizz[17][624] = 9'b111111111;
assign micromatrizz[17][625] = 9'b111111111;
assign micromatrizz[17][626] = 9'b111111111;
assign micromatrizz[17][627] = 9'b111111111;
assign micromatrizz[17][628] = 9'b111111111;
assign micromatrizz[17][629] = 9'b111111111;
assign micromatrizz[17][630] = 9'b111111111;
assign micromatrizz[17][631] = 9'b111111111;
assign micromatrizz[17][632] = 9'b111111111;
assign micromatrizz[17][633] = 9'b111111111;
assign micromatrizz[17][634] = 9'b111111111;
assign micromatrizz[17][635] = 9'b111111111;
assign micromatrizz[17][636] = 9'b111111111;
assign micromatrizz[17][637] = 9'b111111111;
assign micromatrizz[17][638] = 9'b111111111;
assign micromatrizz[17][639] = 9'b111111111;
assign micromatrizz[18][0] = 9'b111111111;
assign micromatrizz[18][1] = 9'b111111111;
assign micromatrizz[18][2] = 9'b111111111;
assign micromatrizz[18][3] = 9'b111111111;
assign micromatrizz[18][4] = 9'b111111111;
assign micromatrizz[18][5] = 9'b111111111;
assign micromatrizz[18][6] = 9'b111111111;
assign micromatrizz[18][7] = 9'b111111111;
assign micromatrizz[18][8] = 9'b111111111;
assign micromatrizz[18][9] = 9'b111111111;
assign micromatrizz[18][10] = 9'b111111111;
assign micromatrizz[18][11] = 9'b111111111;
assign micromatrizz[18][12] = 9'b111111111;
assign micromatrizz[18][13] = 9'b111111111;
assign micromatrizz[18][14] = 9'b111111111;
assign micromatrizz[18][15] = 9'b111111111;
assign micromatrizz[18][16] = 9'b111111111;
assign micromatrizz[18][17] = 9'b111111111;
assign micromatrizz[18][18] = 9'b111111111;
assign micromatrizz[18][19] = 9'b111111111;
assign micromatrizz[18][20] = 9'b111111111;
assign micromatrizz[18][21] = 9'b111111111;
assign micromatrizz[18][22] = 9'b111111111;
assign micromatrizz[18][23] = 9'b111111111;
assign micromatrizz[18][24] = 9'b111111111;
assign micromatrizz[18][25] = 9'b111111111;
assign micromatrizz[18][26] = 9'b111111111;
assign micromatrizz[18][27] = 9'b111111111;
assign micromatrizz[18][28] = 9'b111111111;
assign micromatrizz[18][29] = 9'b111111111;
assign micromatrizz[18][30] = 9'b111111111;
assign micromatrizz[18][31] = 9'b111111111;
assign micromatrizz[18][32] = 9'b111111111;
assign micromatrizz[18][33] = 9'b111111111;
assign micromatrizz[18][34] = 9'b111111111;
assign micromatrizz[18][35] = 9'b111111111;
assign micromatrizz[18][36] = 9'b111111111;
assign micromatrizz[18][37] = 9'b111111111;
assign micromatrizz[18][38] = 9'b111111111;
assign micromatrizz[18][39] = 9'b111111111;
assign micromatrizz[18][40] = 9'b111111111;
assign micromatrizz[18][41] = 9'b111111111;
assign micromatrizz[18][42] = 9'b111111111;
assign micromatrizz[18][43] = 9'b111111111;
assign micromatrizz[18][44] = 9'b111111111;
assign micromatrizz[18][45] = 9'b111111111;
assign micromatrizz[18][46] = 9'b111111111;
assign micromatrizz[18][47] = 9'b111111111;
assign micromatrizz[18][48] = 9'b111111111;
assign micromatrizz[18][49] = 9'b111111111;
assign micromatrizz[18][50] = 9'b111111111;
assign micromatrizz[18][51] = 9'b111111111;
assign micromatrizz[18][52] = 9'b111111111;
assign micromatrizz[18][53] = 9'b111111111;
assign micromatrizz[18][54] = 9'b111111111;
assign micromatrizz[18][55] = 9'b111111111;
assign micromatrizz[18][56] = 9'b111111111;
assign micromatrizz[18][57] = 9'b111111111;
assign micromatrizz[18][58] = 9'b111111111;
assign micromatrizz[18][59] = 9'b111111111;
assign micromatrizz[18][60] = 9'b111111111;
assign micromatrizz[18][61] = 9'b111111111;
assign micromatrizz[18][62] = 9'b111111111;
assign micromatrizz[18][63] = 9'b111111111;
assign micromatrizz[18][64] = 9'b111111111;
assign micromatrizz[18][65] = 9'b111111111;
assign micromatrizz[18][66] = 9'b111111111;
assign micromatrizz[18][67] = 9'b111111111;
assign micromatrizz[18][68] = 9'b111111111;
assign micromatrizz[18][69] = 9'b111111111;
assign micromatrizz[18][70] = 9'b111111111;
assign micromatrizz[18][71] = 9'b111111111;
assign micromatrizz[18][72] = 9'b111111111;
assign micromatrizz[18][73] = 9'b111111111;
assign micromatrizz[18][74] = 9'b111111111;
assign micromatrizz[18][75] = 9'b111111111;
assign micromatrizz[18][76] = 9'b111111111;
assign micromatrizz[18][77] = 9'b111111111;
assign micromatrizz[18][78] = 9'b111111111;
assign micromatrizz[18][79] = 9'b111111111;
assign micromatrizz[18][80] = 9'b111111111;
assign micromatrizz[18][81] = 9'b111111111;
assign micromatrizz[18][82] = 9'b111111111;
assign micromatrizz[18][83] = 9'b111111111;
assign micromatrizz[18][84] = 9'b111111111;
assign micromatrizz[18][85] = 9'b111111111;
assign micromatrizz[18][86] = 9'b111111111;
assign micromatrizz[18][87] = 9'b111111111;
assign micromatrizz[18][88] = 9'b111111111;
assign micromatrizz[18][89] = 9'b111111111;
assign micromatrizz[18][90] = 9'b111111111;
assign micromatrizz[18][91] = 9'b111111111;
assign micromatrizz[18][92] = 9'b111111111;
assign micromatrizz[18][93] = 9'b111111111;
assign micromatrizz[18][94] = 9'b111111111;
assign micromatrizz[18][95] = 9'b111111111;
assign micromatrizz[18][96] = 9'b111111111;
assign micromatrizz[18][97] = 9'b111111111;
assign micromatrizz[18][98] = 9'b111111111;
assign micromatrizz[18][99] = 9'b111111111;
assign micromatrizz[18][100] = 9'b111111111;
assign micromatrizz[18][101] = 9'b111111111;
assign micromatrizz[18][102] = 9'b111111111;
assign micromatrizz[18][103] = 9'b111111111;
assign micromatrizz[18][104] = 9'b111111111;
assign micromatrizz[18][105] = 9'b111111111;
assign micromatrizz[18][106] = 9'b111111111;
assign micromatrizz[18][107] = 9'b111111111;
assign micromatrizz[18][108] = 9'b111111111;
assign micromatrizz[18][109] = 9'b111111111;
assign micromatrizz[18][110] = 9'b111111111;
assign micromatrizz[18][111] = 9'b111111111;
assign micromatrizz[18][112] = 9'b111111111;
assign micromatrizz[18][113] = 9'b111111111;
assign micromatrizz[18][114] = 9'b111111111;
assign micromatrizz[18][115] = 9'b111111111;
assign micromatrizz[18][116] = 9'b111111111;
assign micromatrizz[18][117] = 9'b111111111;
assign micromatrizz[18][118] = 9'b111111111;
assign micromatrizz[18][119] = 9'b111111111;
assign micromatrizz[18][120] = 9'b111111111;
assign micromatrizz[18][121] = 9'b111111111;
assign micromatrizz[18][122] = 9'b111111111;
assign micromatrizz[18][123] = 9'b111111111;
assign micromatrizz[18][124] = 9'b111111111;
assign micromatrizz[18][125] = 9'b111111111;
assign micromatrizz[18][126] = 9'b111111111;
assign micromatrizz[18][127] = 9'b111111111;
assign micromatrizz[18][128] = 9'b111111111;
assign micromatrizz[18][129] = 9'b111111111;
assign micromatrizz[18][130] = 9'b111111111;
assign micromatrizz[18][131] = 9'b111111111;
assign micromatrizz[18][132] = 9'b111111111;
assign micromatrizz[18][133] = 9'b111111111;
assign micromatrizz[18][134] = 9'b111111111;
assign micromatrizz[18][135] = 9'b111111111;
assign micromatrizz[18][136] = 9'b111111111;
assign micromatrizz[18][137] = 9'b111111111;
assign micromatrizz[18][138] = 9'b111111111;
assign micromatrizz[18][139] = 9'b111111111;
assign micromatrizz[18][140] = 9'b111111111;
assign micromatrizz[18][141] = 9'b111111111;
assign micromatrizz[18][142] = 9'b111111111;
assign micromatrizz[18][143] = 9'b111111111;
assign micromatrizz[18][144] = 9'b111111111;
assign micromatrizz[18][145] = 9'b111111111;
assign micromatrizz[18][146] = 9'b111111111;
assign micromatrizz[18][147] = 9'b111111111;
assign micromatrizz[18][148] = 9'b111111111;
assign micromatrizz[18][149] = 9'b111111111;
assign micromatrizz[18][150] = 9'b111111111;
assign micromatrizz[18][151] = 9'b111111111;
assign micromatrizz[18][152] = 9'b111111111;
assign micromatrizz[18][153] = 9'b111111111;
assign micromatrizz[18][154] = 9'b111111111;
assign micromatrizz[18][155] = 9'b111111111;
assign micromatrizz[18][156] = 9'b111111111;
assign micromatrizz[18][157] = 9'b111111111;
assign micromatrizz[18][158] = 9'b111111111;
assign micromatrizz[18][159] = 9'b111111111;
assign micromatrizz[18][160] = 9'b111111111;
assign micromatrizz[18][161] = 9'b111111111;
assign micromatrizz[18][162] = 9'b111111111;
assign micromatrizz[18][163] = 9'b111111111;
assign micromatrizz[18][164] = 9'b111111111;
assign micromatrizz[18][165] = 9'b111111111;
assign micromatrizz[18][166] = 9'b111111111;
assign micromatrizz[18][167] = 9'b111111111;
assign micromatrizz[18][168] = 9'b111111111;
assign micromatrizz[18][169] = 9'b111111111;
assign micromatrizz[18][170] = 9'b111111111;
assign micromatrizz[18][171] = 9'b111111111;
assign micromatrizz[18][172] = 9'b111111111;
assign micromatrizz[18][173] = 9'b111111111;
assign micromatrizz[18][174] = 9'b111111111;
assign micromatrizz[18][175] = 9'b111111111;
assign micromatrizz[18][176] = 9'b111111111;
assign micromatrizz[18][177] = 9'b111111111;
assign micromatrizz[18][178] = 9'b111111111;
assign micromatrizz[18][179] = 9'b111111111;
assign micromatrizz[18][180] = 9'b111111111;
assign micromatrizz[18][181] = 9'b111111111;
assign micromatrizz[18][182] = 9'b111111111;
assign micromatrizz[18][183] = 9'b111111111;
assign micromatrizz[18][184] = 9'b111111111;
assign micromatrizz[18][185] = 9'b111111111;
assign micromatrizz[18][186] = 9'b111111111;
assign micromatrizz[18][187] = 9'b111111111;
assign micromatrizz[18][188] = 9'b111111111;
assign micromatrizz[18][189] = 9'b111111111;
assign micromatrizz[18][190] = 9'b111111111;
assign micromatrizz[18][191] = 9'b111111111;
assign micromatrizz[18][192] = 9'b111111111;
assign micromatrizz[18][193] = 9'b111111111;
assign micromatrizz[18][194] = 9'b111111111;
assign micromatrizz[18][195] = 9'b111111111;
assign micromatrizz[18][196] = 9'b111111111;
assign micromatrizz[18][197] = 9'b111111111;
assign micromatrizz[18][198] = 9'b111111111;
assign micromatrizz[18][199] = 9'b111111111;
assign micromatrizz[18][200] = 9'b111111111;
assign micromatrizz[18][201] = 9'b111111111;
assign micromatrizz[18][202] = 9'b111111111;
assign micromatrizz[18][203] = 9'b111111111;
assign micromatrizz[18][204] = 9'b111111111;
assign micromatrizz[18][205] = 9'b111111111;
assign micromatrizz[18][206] = 9'b111111111;
assign micromatrizz[18][207] = 9'b111111111;
assign micromatrizz[18][208] = 9'b111111111;
assign micromatrizz[18][209] = 9'b111111111;
assign micromatrizz[18][210] = 9'b111111111;
assign micromatrizz[18][211] = 9'b111111111;
assign micromatrizz[18][212] = 9'b111111111;
assign micromatrizz[18][213] = 9'b111111111;
assign micromatrizz[18][214] = 9'b111111111;
assign micromatrizz[18][215] = 9'b111111111;
assign micromatrizz[18][216] = 9'b111111111;
assign micromatrizz[18][217] = 9'b111111111;
assign micromatrizz[18][218] = 9'b111111111;
assign micromatrizz[18][219] = 9'b111111111;
assign micromatrizz[18][220] = 9'b111111111;
assign micromatrizz[18][221] = 9'b111111111;
assign micromatrizz[18][222] = 9'b111111111;
assign micromatrizz[18][223] = 9'b111111111;
assign micromatrizz[18][224] = 9'b111111111;
assign micromatrizz[18][225] = 9'b111111111;
assign micromatrizz[18][226] = 9'b111111111;
assign micromatrizz[18][227] = 9'b111111111;
assign micromatrizz[18][228] = 9'b111111111;
assign micromatrizz[18][229] = 9'b111111111;
assign micromatrizz[18][230] = 9'b111111111;
assign micromatrizz[18][231] = 9'b111111111;
assign micromatrizz[18][232] = 9'b111111111;
assign micromatrizz[18][233] = 9'b111111111;
assign micromatrizz[18][234] = 9'b111111111;
assign micromatrizz[18][235] = 9'b111111111;
assign micromatrizz[18][236] = 9'b111111111;
assign micromatrizz[18][237] = 9'b111111111;
assign micromatrizz[18][238] = 9'b111111111;
assign micromatrizz[18][239] = 9'b111111111;
assign micromatrizz[18][240] = 9'b111111111;
assign micromatrizz[18][241] = 9'b111111111;
assign micromatrizz[18][242] = 9'b111111111;
assign micromatrizz[18][243] = 9'b111111111;
assign micromatrizz[18][244] = 9'b111111111;
assign micromatrizz[18][245] = 9'b111111111;
assign micromatrizz[18][246] = 9'b111111111;
assign micromatrizz[18][247] = 9'b111111111;
assign micromatrizz[18][248] = 9'b111111111;
assign micromatrizz[18][249] = 9'b111111111;
assign micromatrizz[18][250] = 9'b111111111;
assign micromatrizz[18][251] = 9'b111111111;
assign micromatrizz[18][252] = 9'b111111111;
assign micromatrizz[18][253] = 9'b111111111;
assign micromatrizz[18][254] = 9'b111111111;
assign micromatrizz[18][255] = 9'b111111111;
assign micromatrizz[18][256] = 9'b111111111;
assign micromatrizz[18][257] = 9'b111111111;
assign micromatrizz[18][258] = 9'b111111111;
assign micromatrizz[18][259] = 9'b111111111;
assign micromatrizz[18][260] = 9'b111111111;
assign micromatrizz[18][261] = 9'b111111111;
assign micromatrizz[18][262] = 9'b111111111;
assign micromatrizz[18][263] = 9'b111111111;
assign micromatrizz[18][264] = 9'b111111111;
assign micromatrizz[18][265] = 9'b111111111;
assign micromatrizz[18][266] = 9'b111111111;
assign micromatrizz[18][267] = 9'b111111111;
assign micromatrizz[18][268] = 9'b111111111;
assign micromatrizz[18][269] = 9'b111111111;
assign micromatrizz[18][270] = 9'b111110010;
assign micromatrizz[18][271] = 9'b111110010;
assign micromatrizz[18][272] = 9'b111110010;
assign micromatrizz[18][273] = 9'b111110010;
assign micromatrizz[18][274] = 9'b111110010;
assign micromatrizz[18][275] = 9'b111110010;
assign micromatrizz[18][276] = 9'b111110010;
assign micromatrizz[18][277] = 9'b111110010;
assign micromatrizz[18][278] = 9'b111110010;
assign micromatrizz[18][279] = 9'b111111111;
assign micromatrizz[18][280] = 9'b111111111;
assign micromatrizz[18][281] = 9'b111111111;
assign micromatrizz[18][282] = 9'b111111111;
assign micromatrizz[18][283] = 9'b111111111;
assign micromatrizz[18][284] = 9'b111111111;
assign micromatrizz[18][285] = 9'b111111111;
assign micromatrizz[18][286] = 9'b111111111;
assign micromatrizz[18][287] = 9'b111111111;
assign micromatrizz[18][288] = 9'b111111111;
assign micromatrizz[18][289] = 9'b111111111;
assign micromatrizz[18][290] = 9'b111111111;
assign micromatrizz[18][291] = 9'b111111111;
assign micromatrizz[18][292] = 9'b111111111;
assign micromatrizz[18][293] = 9'b111111111;
assign micromatrizz[18][294] = 9'b111111111;
assign micromatrizz[18][295] = 9'b111111111;
assign micromatrizz[18][296] = 9'b111111111;
assign micromatrizz[18][297] = 9'b111111111;
assign micromatrizz[18][298] = 9'b111111111;
assign micromatrizz[18][299] = 9'b111111111;
assign micromatrizz[18][300] = 9'b111111111;
assign micromatrizz[18][301] = 9'b111111111;
assign micromatrizz[18][302] = 9'b111111111;
assign micromatrizz[18][303] = 9'b111111111;
assign micromatrizz[18][304] = 9'b111111111;
assign micromatrizz[18][305] = 9'b111111111;
assign micromatrizz[18][306] = 9'b111111111;
assign micromatrizz[18][307] = 9'b111111111;
assign micromatrizz[18][308] = 9'b111111111;
assign micromatrizz[18][309] = 9'b111111111;
assign micromatrizz[18][310] = 9'b111111111;
assign micromatrizz[18][311] = 9'b111111111;
assign micromatrizz[18][312] = 9'b111111111;
assign micromatrizz[18][313] = 9'b111111111;
assign micromatrizz[18][314] = 9'b111111111;
assign micromatrizz[18][315] = 9'b111111111;
assign micromatrizz[18][316] = 9'b111111111;
assign micromatrizz[18][317] = 9'b111111111;
assign micromatrizz[18][318] = 9'b111111111;
assign micromatrizz[18][319] = 9'b111111111;
assign micromatrizz[18][320] = 9'b111111111;
assign micromatrizz[18][321] = 9'b111111111;
assign micromatrizz[18][322] = 9'b111111111;
assign micromatrizz[18][323] = 9'b111111111;
assign micromatrizz[18][324] = 9'b111111111;
assign micromatrizz[18][325] = 9'b111111111;
assign micromatrizz[18][326] = 9'b111111111;
assign micromatrizz[18][327] = 9'b111111111;
assign micromatrizz[18][328] = 9'b111111111;
assign micromatrizz[18][329] = 9'b111111111;
assign micromatrizz[18][330] = 9'b111111111;
assign micromatrizz[18][331] = 9'b111111111;
assign micromatrizz[18][332] = 9'b111111111;
assign micromatrizz[18][333] = 9'b111111111;
assign micromatrizz[18][334] = 9'b111111111;
assign micromatrizz[18][335] = 9'b111111111;
assign micromatrizz[18][336] = 9'b111111111;
assign micromatrizz[18][337] = 9'b111111111;
assign micromatrizz[18][338] = 9'b111111111;
assign micromatrizz[18][339] = 9'b111111111;
assign micromatrizz[18][340] = 9'b111111111;
assign micromatrizz[18][341] = 9'b111111111;
assign micromatrizz[18][342] = 9'b111111111;
assign micromatrizz[18][343] = 9'b111111111;
assign micromatrizz[18][344] = 9'b111111111;
assign micromatrizz[18][345] = 9'b111111111;
assign micromatrizz[18][346] = 9'b111111111;
assign micromatrizz[18][347] = 9'b111111111;
assign micromatrizz[18][348] = 9'b111111111;
assign micromatrizz[18][349] = 9'b111111111;
assign micromatrizz[18][350] = 9'b111111111;
assign micromatrizz[18][351] = 9'b111111111;
assign micromatrizz[18][352] = 9'b111111111;
assign micromatrizz[18][353] = 9'b111111111;
assign micromatrizz[18][354] = 9'b111111111;
assign micromatrizz[18][355] = 9'b111111111;
assign micromatrizz[18][356] = 9'b111111111;
assign micromatrizz[18][357] = 9'b111111111;
assign micromatrizz[18][358] = 9'b111111111;
assign micromatrizz[18][359] = 9'b111111111;
assign micromatrizz[18][360] = 9'b111111111;
assign micromatrizz[18][361] = 9'b111111111;
assign micromatrizz[18][362] = 9'b111111111;
assign micromatrizz[18][363] = 9'b111111111;
assign micromatrizz[18][364] = 9'b111111111;
assign micromatrizz[18][365] = 9'b111111111;
assign micromatrizz[18][366] = 9'b111111111;
assign micromatrizz[18][367] = 9'b111111111;
assign micromatrizz[18][368] = 9'b111111111;
assign micromatrizz[18][369] = 9'b111111111;
assign micromatrizz[18][370] = 9'b111111111;
assign micromatrizz[18][371] = 9'b111111111;
assign micromatrizz[18][372] = 9'b111111111;
assign micromatrizz[18][373] = 9'b111111111;
assign micromatrizz[18][374] = 9'b111111111;
assign micromatrizz[18][375] = 9'b111111111;
assign micromatrizz[18][376] = 9'b111111111;
assign micromatrizz[18][377] = 9'b111111111;
assign micromatrizz[18][378] = 9'b111111111;
assign micromatrizz[18][379] = 9'b111111111;
assign micromatrizz[18][380] = 9'b111111111;
assign micromatrizz[18][381] = 9'b111111111;
assign micromatrizz[18][382] = 9'b111111111;
assign micromatrizz[18][383] = 9'b111111111;
assign micromatrizz[18][384] = 9'b111111111;
assign micromatrizz[18][385] = 9'b111111111;
assign micromatrizz[18][386] = 9'b111111111;
assign micromatrizz[18][387] = 9'b111111111;
assign micromatrizz[18][388] = 9'b111111111;
assign micromatrizz[18][389] = 9'b111111111;
assign micromatrizz[18][390] = 9'b111111111;
assign micromatrizz[18][391] = 9'b111111111;
assign micromatrizz[18][392] = 9'b111111111;
assign micromatrizz[18][393] = 9'b111111111;
assign micromatrizz[18][394] = 9'b111111111;
assign micromatrizz[18][395] = 9'b111111111;
assign micromatrizz[18][396] = 9'b111111111;
assign micromatrizz[18][397] = 9'b111111111;
assign micromatrizz[18][398] = 9'b111111111;
assign micromatrizz[18][399] = 9'b111111111;
assign micromatrizz[18][400] = 9'b111111111;
assign micromatrizz[18][401] = 9'b111111111;
assign micromatrizz[18][402] = 9'b111111111;
assign micromatrizz[18][403] = 9'b111111111;
assign micromatrizz[18][404] = 9'b111111111;
assign micromatrizz[18][405] = 9'b111111111;
assign micromatrizz[18][406] = 9'b111111111;
assign micromatrizz[18][407] = 9'b111111111;
assign micromatrizz[18][408] = 9'b111111111;
assign micromatrizz[18][409] = 9'b111111111;
assign micromatrizz[18][410] = 9'b111111111;
assign micromatrizz[18][411] = 9'b111111111;
assign micromatrizz[18][412] = 9'b111111111;
assign micromatrizz[18][413] = 9'b111111111;
assign micromatrizz[18][414] = 9'b111111111;
assign micromatrizz[18][415] = 9'b111111111;
assign micromatrizz[18][416] = 9'b111111111;
assign micromatrizz[18][417] = 9'b111111111;
assign micromatrizz[18][418] = 9'b111111111;
assign micromatrizz[18][419] = 9'b111111111;
assign micromatrizz[18][420] = 9'b111111111;
assign micromatrizz[18][421] = 9'b111111111;
assign micromatrizz[18][422] = 9'b111111111;
assign micromatrizz[18][423] = 9'b111111111;
assign micromatrizz[18][424] = 9'b111111111;
assign micromatrizz[18][425] = 9'b111111111;
assign micromatrizz[18][426] = 9'b111111111;
assign micromatrizz[18][427] = 9'b111111111;
assign micromatrizz[18][428] = 9'b111111111;
assign micromatrizz[18][429] = 9'b111111111;
assign micromatrizz[18][430] = 9'b111111111;
assign micromatrizz[18][431] = 9'b111111111;
assign micromatrizz[18][432] = 9'b111111111;
assign micromatrizz[18][433] = 9'b111111111;
assign micromatrizz[18][434] = 9'b111111111;
assign micromatrizz[18][435] = 9'b111111111;
assign micromatrizz[18][436] = 9'b111111111;
assign micromatrizz[18][437] = 9'b111111111;
assign micromatrizz[18][438] = 9'b111111111;
assign micromatrizz[18][439] = 9'b111111111;
assign micromatrizz[18][440] = 9'b111111111;
assign micromatrizz[18][441] = 9'b111111111;
assign micromatrizz[18][442] = 9'b111111111;
assign micromatrizz[18][443] = 9'b111111111;
assign micromatrizz[18][444] = 9'b111111111;
assign micromatrizz[18][445] = 9'b111111111;
assign micromatrizz[18][446] = 9'b111111111;
assign micromatrizz[18][447] = 9'b111111111;
assign micromatrizz[18][448] = 9'b111111111;
assign micromatrizz[18][449] = 9'b111111111;
assign micromatrizz[18][450] = 9'b111111111;
assign micromatrizz[18][451] = 9'b111111111;
assign micromatrizz[18][452] = 9'b111111111;
assign micromatrizz[18][453] = 9'b111111111;
assign micromatrizz[18][454] = 9'b111111111;
assign micromatrizz[18][455] = 9'b111111111;
assign micromatrizz[18][456] = 9'b111111111;
assign micromatrizz[18][457] = 9'b111111111;
assign micromatrizz[18][458] = 9'b111111111;
assign micromatrizz[18][459] = 9'b111111111;
assign micromatrizz[18][460] = 9'b111111111;
assign micromatrizz[18][461] = 9'b111111111;
assign micromatrizz[18][462] = 9'b111111111;
assign micromatrizz[18][463] = 9'b111111111;
assign micromatrizz[18][464] = 9'b111111111;
assign micromatrizz[18][465] = 9'b111111111;
assign micromatrizz[18][466] = 9'b111111111;
assign micromatrizz[18][467] = 9'b111111111;
assign micromatrizz[18][468] = 9'b111111111;
assign micromatrizz[18][469] = 9'b111111111;
assign micromatrizz[18][470] = 9'b111111111;
assign micromatrizz[18][471] = 9'b111111111;
assign micromatrizz[18][472] = 9'b111111111;
assign micromatrizz[18][473] = 9'b111111111;
assign micromatrizz[18][474] = 9'b111111111;
assign micromatrizz[18][475] = 9'b111111111;
assign micromatrizz[18][476] = 9'b111111111;
assign micromatrizz[18][477] = 9'b111111111;
assign micromatrizz[18][478] = 9'b111111111;
assign micromatrizz[18][479] = 9'b111111111;
assign micromatrizz[18][480] = 9'b111111111;
assign micromatrizz[18][481] = 9'b111111111;
assign micromatrizz[18][482] = 9'b111111111;
assign micromatrizz[18][483] = 9'b111111111;
assign micromatrizz[18][484] = 9'b111111111;
assign micromatrizz[18][485] = 9'b111111111;
assign micromatrizz[18][486] = 9'b111111111;
assign micromatrizz[18][487] = 9'b111111111;
assign micromatrizz[18][488] = 9'b111111111;
assign micromatrizz[18][489] = 9'b111111111;
assign micromatrizz[18][490] = 9'b111111111;
assign micromatrizz[18][491] = 9'b111111111;
assign micromatrizz[18][492] = 9'b111111111;
assign micromatrizz[18][493] = 9'b111111111;
assign micromatrizz[18][494] = 9'b111111111;
assign micromatrizz[18][495] = 9'b111111111;
assign micromatrizz[18][496] = 9'b111111111;
assign micromatrizz[18][497] = 9'b111111111;
assign micromatrizz[18][498] = 9'b111111111;
assign micromatrizz[18][499] = 9'b111111111;
assign micromatrizz[18][500] = 9'b111111111;
assign micromatrizz[18][501] = 9'b111111111;
assign micromatrizz[18][502] = 9'b111111111;
assign micromatrizz[18][503] = 9'b111111111;
assign micromatrizz[18][504] = 9'b111111111;
assign micromatrizz[18][505] = 9'b111111111;
assign micromatrizz[18][506] = 9'b111111111;
assign micromatrizz[18][507] = 9'b111111111;
assign micromatrizz[18][508] = 9'b111111111;
assign micromatrizz[18][509] = 9'b111111111;
assign micromatrizz[18][510] = 9'b111111111;
assign micromatrizz[18][511] = 9'b111111111;
assign micromatrizz[18][512] = 9'b111111111;
assign micromatrizz[18][513] = 9'b111111111;
assign micromatrizz[18][514] = 9'b111111111;
assign micromatrizz[18][515] = 9'b111111111;
assign micromatrizz[18][516] = 9'b111111111;
assign micromatrizz[18][517] = 9'b111111111;
assign micromatrizz[18][518] = 9'b111111111;
assign micromatrizz[18][519] = 9'b111111111;
assign micromatrizz[18][520] = 9'b111111111;
assign micromatrizz[18][521] = 9'b111111111;
assign micromatrizz[18][522] = 9'b111111111;
assign micromatrizz[18][523] = 9'b111111111;
assign micromatrizz[18][524] = 9'b111111111;
assign micromatrizz[18][525] = 9'b111111111;
assign micromatrizz[18][526] = 9'b111111111;
assign micromatrizz[18][527] = 9'b111111111;
assign micromatrizz[18][528] = 9'b111111111;
assign micromatrizz[18][529] = 9'b111111111;
assign micromatrizz[18][530] = 9'b111111111;
assign micromatrizz[18][531] = 9'b111111111;
assign micromatrizz[18][532] = 9'b111111111;
assign micromatrizz[18][533] = 9'b111111111;
assign micromatrizz[18][534] = 9'b111111111;
assign micromatrizz[18][535] = 9'b111111111;
assign micromatrizz[18][536] = 9'b111111111;
assign micromatrizz[18][537] = 9'b111111111;
assign micromatrizz[18][538] = 9'b111111111;
assign micromatrizz[18][539] = 9'b111111111;
assign micromatrizz[18][540] = 9'b111111111;
assign micromatrizz[18][541] = 9'b111111111;
assign micromatrizz[18][542] = 9'b111111111;
assign micromatrizz[18][543] = 9'b111111111;
assign micromatrizz[18][544] = 9'b111111111;
assign micromatrizz[18][545] = 9'b111111111;
assign micromatrizz[18][546] = 9'b111111111;
assign micromatrizz[18][547] = 9'b111111111;
assign micromatrizz[18][548] = 9'b111111111;
assign micromatrizz[18][549] = 9'b111111111;
assign micromatrizz[18][550] = 9'b111111111;
assign micromatrizz[18][551] = 9'b111111111;
assign micromatrizz[18][552] = 9'b111111111;
assign micromatrizz[18][553] = 9'b111111111;
assign micromatrizz[18][554] = 9'b111111111;
assign micromatrizz[18][555] = 9'b111111111;
assign micromatrizz[18][556] = 9'b111111111;
assign micromatrizz[18][557] = 9'b111111111;
assign micromatrizz[18][558] = 9'b111111111;
assign micromatrizz[18][559] = 9'b111111111;
assign micromatrizz[18][560] = 9'b111111111;
assign micromatrizz[18][561] = 9'b111111111;
assign micromatrizz[18][562] = 9'b111111111;
assign micromatrizz[18][563] = 9'b111111111;
assign micromatrizz[18][564] = 9'b111111111;
assign micromatrizz[18][565] = 9'b111111111;
assign micromatrizz[18][566] = 9'b111111111;
assign micromatrizz[18][567] = 9'b111111111;
assign micromatrizz[18][568] = 9'b111111111;
assign micromatrizz[18][569] = 9'b111111111;
assign micromatrizz[18][570] = 9'b111111111;
assign micromatrizz[18][571] = 9'b111111111;
assign micromatrizz[18][572] = 9'b111111111;
assign micromatrizz[18][573] = 9'b111111111;
assign micromatrizz[18][574] = 9'b111111111;
assign micromatrizz[18][575] = 9'b111111111;
assign micromatrizz[18][576] = 9'b111111111;
assign micromatrizz[18][577] = 9'b111111111;
assign micromatrizz[18][578] = 9'b111111111;
assign micromatrizz[18][579] = 9'b111111111;
assign micromatrizz[18][580] = 9'b111111111;
assign micromatrizz[18][581] = 9'b111111111;
assign micromatrizz[18][582] = 9'b111111111;
assign micromatrizz[18][583] = 9'b111111111;
assign micromatrizz[18][584] = 9'b111111111;
assign micromatrizz[18][585] = 9'b111111111;
assign micromatrizz[18][586] = 9'b111111111;
assign micromatrizz[18][587] = 9'b111111111;
assign micromatrizz[18][588] = 9'b111111111;
assign micromatrizz[18][589] = 9'b111111111;
assign micromatrizz[18][590] = 9'b111111111;
assign micromatrizz[18][591] = 9'b111111111;
assign micromatrizz[18][592] = 9'b111111111;
assign micromatrizz[18][593] = 9'b111111111;
assign micromatrizz[18][594] = 9'b111111111;
assign micromatrizz[18][595] = 9'b111111111;
assign micromatrizz[18][596] = 9'b111111111;
assign micromatrizz[18][597] = 9'b111111111;
assign micromatrizz[18][598] = 9'b111111111;
assign micromatrizz[18][599] = 9'b111111111;
assign micromatrizz[18][600] = 9'b111111111;
assign micromatrizz[18][601] = 9'b111111111;
assign micromatrizz[18][602] = 9'b111111111;
assign micromatrizz[18][603] = 9'b111111111;
assign micromatrizz[18][604] = 9'b111111111;
assign micromatrizz[18][605] = 9'b111111111;
assign micromatrizz[18][606] = 9'b111111111;
assign micromatrizz[18][607] = 9'b111111111;
assign micromatrizz[18][608] = 9'b111111111;
assign micromatrizz[18][609] = 9'b111111111;
assign micromatrizz[18][610] = 9'b111111111;
assign micromatrizz[18][611] = 9'b111111111;
assign micromatrizz[18][612] = 9'b111111111;
assign micromatrizz[18][613] = 9'b111111111;
assign micromatrizz[18][614] = 9'b111111111;
assign micromatrizz[18][615] = 9'b111111111;
assign micromatrizz[18][616] = 9'b111111111;
assign micromatrizz[18][617] = 9'b111111111;
assign micromatrizz[18][618] = 9'b111111111;
assign micromatrizz[18][619] = 9'b111111111;
assign micromatrizz[18][620] = 9'b111111111;
assign micromatrizz[18][621] = 9'b111111111;
assign micromatrizz[18][622] = 9'b111111111;
assign micromatrizz[18][623] = 9'b111111111;
assign micromatrizz[18][624] = 9'b111111111;
assign micromatrizz[18][625] = 9'b111111111;
assign micromatrizz[18][626] = 9'b111111111;
assign micromatrizz[18][627] = 9'b111111111;
assign micromatrizz[18][628] = 9'b111111111;
assign micromatrizz[18][629] = 9'b111111111;
assign micromatrizz[18][630] = 9'b111111111;
assign micromatrizz[18][631] = 9'b111111111;
assign micromatrizz[18][632] = 9'b111111111;
assign micromatrizz[18][633] = 9'b111111111;
assign micromatrizz[18][634] = 9'b111111111;
assign micromatrizz[18][635] = 9'b111111111;
assign micromatrizz[18][636] = 9'b111111111;
assign micromatrizz[18][637] = 9'b111111111;
assign micromatrizz[18][638] = 9'b111111111;
assign micromatrizz[18][639] = 9'b111111111;
assign micromatrizz[19][0] = 9'b111111111;
assign micromatrizz[19][1] = 9'b111111111;
assign micromatrizz[19][2] = 9'b111111111;
assign micromatrizz[19][3] = 9'b111111111;
assign micromatrizz[19][4] = 9'b111111111;
assign micromatrizz[19][5] = 9'b111111111;
assign micromatrizz[19][6] = 9'b111111111;
assign micromatrizz[19][7] = 9'b111111111;
assign micromatrizz[19][8] = 9'b111111111;
assign micromatrizz[19][9] = 9'b111111111;
assign micromatrizz[19][10] = 9'b111111111;
assign micromatrizz[19][11] = 9'b111111111;
assign micromatrizz[19][12] = 9'b111111111;
assign micromatrizz[19][13] = 9'b111111111;
assign micromatrizz[19][14] = 9'b111111111;
assign micromatrizz[19][15] = 9'b111111111;
assign micromatrizz[19][16] = 9'b111111111;
assign micromatrizz[19][17] = 9'b111111111;
assign micromatrizz[19][18] = 9'b111111111;
assign micromatrizz[19][19] = 9'b111111111;
assign micromatrizz[19][20] = 9'b111111111;
assign micromatrizz[19][21] = 9'b111111111;
assign micromatrizz[19][22] = 9'b111111111;
assign micromatrizz[19][23] = 9'b111111111;
assign micromatrizz[19][24] = 9'b111111111;
assign micromatrizz[19][25] = 9'b111111111;
assign micromatrizz[19][26] = 9'b111111111;
assign micromatrizz[19][27] = 9'b111111111;
assign micromatrizz[19][28] = 9'b111111111;
assign micromatrizz[19][29] = 9'b111111111;
assign micromatrizz[19][30] = 9'b111111111;
assign micromatrizz[19][31] = 9'b111111111;
assign micromatrizz[19][32] = 9'b111111111;
assign micromatrizz[19][33] = 9'b111111111;
assign micromatrizz[19][34] = 9'b111111111;
assign micromatrizz[19][35] = 9'b111111111;
assign micromatrizz[19][36] = 9'b111111111;
assign micromatrizz[19][37] = 9'b111111111;
assign micromatrizz[19][38] = 9'b111111111;
assign micromatrizz[19][39] = 9'b111111111;
assign micromatrizz[19][40] = 9'b111111111;
assign micromatrizz[19][41] = 9'b111111111;
assign micromatrizz[19][42] = 9'b111111111;
assign micromatrizz[19][43] = 9'b111111111;
assign micromatrizz[19][44] = 9'b111111111;
assign micromatrizz[19][45] = 9'b111111111;
assign micromatrizz[19][46] = 9'b111111111;
assign micromatrizz[19][47] = 9'b111111111;
assign micromatrizz[19][48] = 9'b111111111;
assign micromatrizz[19][49] = 9'b111111111;
assign micromatrizz[19][50] = 9'b111111111;
assign micromatrizz[19][51] = 9'b111111111;
assign micromatrizz[19][52] = 9'b111111111;
assign micromatrizz[19][53] = 9'b111111111;
assign micromatrizz[19][54] = 9'b111111111;
assign micromatrizz[19][55] = 9'b111111111;
assign micromatrizz[19][56] = 9'b111111111;
assign micromatrizz[19][57] = 9'b111111111;
assign micromatrizz[19][58] = 9'b111111111;
assign micromatrizz[19][59] = 9'b111111111;
assign micromatrizz[19][60] = 9'b111111111;
assign micromatrizz[19][61] = 9'b111111111;
assign micromatrizz[19][62] = 9'b111111111;
assign micromatrizz[19][63] = 9'b111111111;
assign micromatrizz[19][64] = 9'b111111111;
assign micromatrizz[19][65] = 9'b111111111;
assign micromatrizz[19][66] = 9'b111111111;
assign micromatrizz[19][67] = 9'b111111111;
assign micromatrizz[19][68] = 9'b111111111;
assign micromatrizz[19][69] = 9'b111111111;
assign micromatrizz[19][70] = 9'b111111111;
assign micromatrizz[19][71] = 9'b111111111;
assign micromatrizz[19][72] = 9'b111111111;
assign micromatrizz[19][73] = 9'b111111111;
assign micromatrizz[19][74] = 9'b111111111;
assign micromatrizz[19][75] = 9'b111111111;
assign micromatrizz[19][76] = 9'b111111111;
assign micromatrizz[19][77] = 9'b111111111;
assign micromatrizz[19][78] = 9'b111111111;
assign micromatrizz[19][79] = 9'b111111111;
assign micromatrizz[19][80] = 9'b111111111;
assign micromatrizz[19][81] = 9'b111111111;
assign micromatrizz[19][82] = 9'b111111111;
assign micromatrizz[19][83] = 9'b111111111;
assign micromatrizz[19][84] = 9'b111111111;
assign micromatrizz[19][85] = 9'b111111111;
assign micromatrizz[19][86] = 9'b111111111;
assign micromatrizz[19][87] = 9'b111111111;
assign micromatrizz[19][88] = 9'b111111111;
assign micromatrizz[19][89] = 9'b111111111;
assign micromatrizz[19][90] = 9'b111111111;
assign micromatrizz[19][91] = 9'b111111111;
assign micromatrizz[19][92] = 9'b111111111;
assign micromatrizz[19][93] = 9'b111111111;
assign micromatrizz[19][94] = 9'b111111111;
assign micromatrizz[19][95] = 9'b111111111;
assign micromatrizz[19][96] = 9'b111111111;
assign micromatrizz[19][97] = 9'b111111111;
assign micromatrizz[19][98] = 9'b111111111;
assign micromatrizz[19][99] = 9'b111111111;
assign micromatrizz[19][100] = 9'b111111111;
assign micromatrizz[19][101] = 9'b111111111;
assign micromatrizz[19][102] = 9'b111111111;
assign micromatrizz[19][103] = 9'b111111111;
assign micromatrizz[19][104] = 9'b111111111;
assign micromatrizz[19][105] = 9'b111111111;
assign micromatrizz[19][106] = 9'b111111111;
assign micromatrizz[19][107] = 9'b111111111;
assign micromatrizz[19][108] = 9'b111111111;
assign micromatrizz[19][109] = 9'b111111111;
assign micromatrizz[19][110] = 9'b111111111;
assign micromatrizz[19][111] = 9'b111111111;
assign micromatrizz[19][112] = 9'b111111111;
assign micromatrizz[19][113] = 9'b111111111;
assign micromatrizz[19][114] = 9'b111111111;
assign micromatrizz[19][115] = 9'b111111111;
assign micromatrizz[19][116] = 9'b111111111;
assign micromatrizz[19][117] = 9'b111111111;
assign micromatrizz[19][118] = 9'b111111111;
assign micromatrizz[19][119] = 9'b111111111;
assign micromatrizz[19][120] = 9'b111111111;
assign micromatrizz[19][121] = 9'b111111111;
assign micromatrizz[19][122] = 9'b111111111;
assign micromatrizz[19][123] = 9'b111111111;
assign micromatrizz[19][124] = 9'b111111111;
assign micromatrizz[19][125] = 9'b111111111;
assign micromatrizz[19][126] = 9'b111111111;
assign micromatrizz[19][127] = 9'b111111111;
assign micromatrizz[19][128] = 9'b111111111;
assign micromatrizz[19][129] = 9'b111111111;
assign micromatrizz[19][130] = 9'b111111111;
assign micromatrizz[19][131] = 9'b111111111;
assign micromatrizz[19][132] = 9'b111111111;
assign micromatrizz[19][133] = 9'b111111111;
assign micromatrizz[19][134] = 9'b111111111;
assign micromatrizz[19][135] = 9'b111111111;
assign micromatrizz[19][136] = 9'b111111111;
assign micromatrizz[19][137] = 9'b111111111;
assign micromatrizz[19][138] = 9'b111111111;
assign micromatrizz[19][139] = 9'b111111111;
assign micromatrizz[19][140] = 9'b111111111;
assign micromatrizz[19][141] = 9'b111111111;
assign micromatrizz[19][142] = 9'b111111111;
assign micromatrizz[19][143] = 9'b111111111;
assign micromatrizz[19][144] = 9'b111111111;
assign micromatrizz[19][145] = 9'b111111111;
assign micromatrizz[19][146] = 9'b111111111;
assign micromatrizz[19][147] = 9'b111111111;
assign micromatrizz[19][148] = 9'b111111111;
assign micromatrizz[19][149] = 9'b111111111;
assign micromatrizz[19][150] = 9'b111111111;
assign micromatrizz[19][151] = 9'b111111111;
assign micromatrizz[19][152] = 9'b111111111;
assign micromatrizz[19][153] = 9'b111111111;
assign micromatrizz[19][154] = 9'b111111111;
assign micromatrizz[19][155] = 9'b111111111;
assign micromatrizz[19][156] = 9'b111111111;
assign micromatrizz[19][157] = 9'b111111111;
assign micromatrizz[19][158] = 9'b111111111;
assign micromatrizz[19][159] = 9'b111111111;
assign micromatrizz[19][160] = 9'b111111111;
assign micromatrizz[19][161] = 9'b111111111;
assign micromatrizz[19][162] = 9'b111111111;
assign micromatrizz[19][163] = 9'b111111111;
assign micromatrizz[19][164] = 9'b111111111;
assign micromatrizz[19][165] = 9'b111111111;
assign micromatrizz[19][166] = 9'b111111111;
assign micromatrizz[19][167] = 9'b111111111;
assign micromatrizz[19][168] = 9'b111111111;
assign micromatrizz[19][169] = 9'b111111111;
assign micromatrizz[19][170] = 9'b111111111;
assign micromatrizz[19][171] = 9'b111111111;
assign micromatrizz[19][172] = 9'b111111111;
assign micromatrizz[19][173] = 9'b111111111;
assign micromatrizz[19][174] = 9'b111111111;
assign micromatrizz[19][175] = 9'b111111111;
assign micromatrizz[19][176] = 9'b111111111;
assign micromatrizz[19][177] = 9'b111111111;
assign micromatrizz[19][178] = 9'b111111111;
assign micromatrizz[19][179] = 9'b111111111;
assign micromatrizz[19][180] = 9'b111111111;
assign micromatrizz[19][181] = 9'b111111111;
assign micromatrizz[19][182] = 9'b111111111;
assign micromatrizz[19][183] = 9'b111111111;
assign micromatrizz[19][184] = 9'b111111111;
assign micromatrizz[19][185] = 9'b111111111;
assign micromatrizz[19][186] = 9'b111111111;
assign micromatrizz[19][187] = 9'b111111111;
assign micromatrizz[19][188] = 9'b111111111;
assign micromatrizz[19][189] = 9'b111111111;
assign micromatrizz[19][190] = 9'b111111111;
assign micromatrizz[19][191] = 9'b111111111;
assign micromatrizz[19][192] = 9'b111111111;
assign micromatrizz[19][193] = 9'b111111111;
assign micromatrizz[19][194] = 9'b111111111;
assign micromatrizz[19][195] = 9'b111111111;
assign micromatrizz[19][196] = 9'b111111111;
assign micromatrizz[19][197] = 9'b111111111;
assign micromatrizz[19][198] = 9'b111111111;
assign micromatrizz[19][199] = 9'b111111111;
assign micromatrizz[19][200] = 9'b111111111;
assign micromatrizz[19][201] = 9'b111111111;
assign micromatrizz[19][202] = 9'b111111111;
assign micromatrizz[19][203] = 9'b111111111;
assign micromatrizz[19][204] = 9'b111111111;
assign micromatrizz[19][205] = 9'b111111111;
assign micromatrizz[19][206] = 9'b111111111;
assign micromatrizz[19][207] = 9'b111111111;
assign micromatrizz[19][208] = 9'b111111111;
assign micromatrizz[19][209] = 9'b111111111;
assign micromatrizz[19][210] = 9'b111111111;
assign micromatrizz[19][211] = 9'b111111111;
assign micromatrizz[19][212] = 9'b111111111;
assign micromatrizz[19][213] = 9'b111111111;
assign micromatrizz[19][214] = 9'b111111111;
assign micromatrizz[19][215] = 9'b111111111;
assign micromatrizz[19][216] = 9'b111111111;
assign micromatrizz[19][217] = 9'b111111111;
assign micromatrizz[19][218] = 9'b111111111;
assign micromatrizz[19][219] = 9'b111111111;
assign micromatrizz[19][220] = 9'b111111111;
assign micromatrizz[19][221] = 9'b111111111;
assign micromatrizz[19][222] = 9'b111111111;
assign micromatrizz[19][223] = 9'b111111111;
assign micromatrizz[19][224] = 9'b111111111;
assign micromatrizz[19][225] = 9'b111111111;
assign micromatrizz[19][226] = 9'b111111111;
assign micromatrizz[19][227] = 9'b111111111;
assign micromatrizz[19][228] = 9'b111111111;
assign micromatrizz[19][229] = 9'b111111111;
assign micromatrizz[19][230] = 9'b111111111;
assign micromatrizz[19][231] = 9'b111111111;
assign micromatrizz[19][232] = 9'b111111111;
assign micromatrizz[19][233] = 9'b111111111;
assign micromatrizz[19][234] = 9'b111111111;
assign micromatrizz[19][235] = 9'b111111111;
assign micromatrizz[19][236] = 9'b111111111;
assign micromatrizz[19][237] = 9'b111111111;
assign micromatrizz[19][238] = 9'b111111111;
assign micromatrizz[19][239] = 9'b111111111;
assign micromatrizz[19][240] = 9'b111111111;
assign micromatrizz[19][241] = 9'b111111111;
assign micromatrizz[19][242] = 9'b111111111;
assign micromatrizz[19][243] = 9'b111111111;
assign micromatrizz[19][244] = 9'b111111111;
assign micromatrizz[19][245] = 9'b111111111;
assign micromatrizz[19][246] = 9'b111111111;
assign micromatrizz[19][247] = 9'b111111111;
assign micromatrizz[19][248] = 9'b111111111;
assign micromatrizz[19][249] = 9'b111111111;
assign micromatrizz[19][250] = 9'b111111111;
assign micromatrizz[19][251] = 9'b111111111;
assign micromatrizz[19][252] = 9'b111111111;
assign micromatrizz[19][253] = 9'b111111111;
assign micromatrizz[19][254] = 9'b111111111;
assign micromatrizz[19][255] = 9'b111111111;
assign micromatrizz[19][256] = 9'b111111111;
assign micromatrizz[19][257] = 9'b111111111;
assign micromatrizz[19][258] = 9'b111111111;
assign micromatrizz[19][259] = 9'b111111111;
assign micromatrizz[19][260] = 9'b111111111;
assign micromatrizz[19][261] = 9'b111111111;
assign micromatrizz[19][262] = 9'b111111111;
assign micromatrizz[19][263] = 9'b111111111;
assign micromatrizz[19][264] = 9'b111111111;
assign micromatrizz[19][265] = 9'b111111111;
assign micromatrizz[19][266] = 9'b111111111;
assign micromatrizz[19][267] = 9'b111111111;
assign micromatrizz[19][268] = 9'b111111111;
assign micromatrizz[19][269] = 9'b111111111;
assign micromatrizz[19][270] = 9'b111110010;
assign micromatrizz[19][271] = 9'b111110010;
assign micromatrizz[19][272] = 9'b111110010;
assign micromatrizz[19][273] = 9'b111110010;
assign micromatrizz[19][274] = 9'b111110011;
assign micromatrizz[19][275] = 9'b111110011;
assign micromatrizz[19][276] = 9'b111110011;
assign micromatrizz[19][277] = 9'b111110010;
assign micromatrizz[19][278] = 9'b111110011;
assign micromatrizz[19][279] = 9'b111111111;
assign micromatrizz[19][280] = 9'b111111111;
assign micromatrizz[19][281] = 9'b111111111;
assign micromatrizz[19][282] = 9'b111111111;
assign micromatrizz[19][283] = 9'b111111111;
assign micromatrizz[19][284] = 9'b111111111;
assign micromatrizz[19][285] = 9'b111111111;
assign micromatrizz[19][286] = 9'b111111111;
assign micromatrizz[19][287] = 9'b111111111;
assign micromatrizz[19][288] = 9'b111111111;
assign micromatrizz[19][289] = 9'b111111111;
assign micromatrizz[19][290] = 9'b111111111;
assign micromatrizz[19][291] = 9'b111111111;
assign micromatrizz[19][292] = 9'b111111111;
assign micromatrizz[19][293] = 9'b111111111;
assign micromatrizz[19][294] = 9'b111111111;
assign micromatrizz[19][295] = 9'b111111111;
assign micromatrizz[19][296] = 9'b111111111;
assign micromatrizz[19][297] = 9'b111111111;
assign micromatrizz[19][298] = 9'b111111111;
assign micromatrizz[19][299] = 9'b111111111;
assign micromatrizz[19][300] = 9'b111111111;
assign micromatrizz[19][301] = 9'b111111111;
assign micromatrizz[19][302] = 9'b111111111;
assign micromatrizz[19][303] = 9'b111111111;
assign micromatrizz[19][304] = 9'b111111111;
assign micromatrizz[19][305] = 9'b111111111;
assign micromatrizz[19][306] = 9'b111111111;
assign micromatrizz[19][307] = 9'b111111111;
assign micromatrizz[19][308] = 9'b111111111;
assign micromatrizz[19][309] = 9'b111111111;
assign micromatrizz[19][310] = 9'b111111111;
assign micromatrizz[19][311] = 9'b111111111;
assign micromatrizz[19][312] = 9'b111111111;
assign micromatrizz[19][313] = 9'b111111111;
assign micromatrizz[19][314] = 9'b111111111;
assign micromatrizz[19][315] = 9'b111111111;
assign micromatrizz[19][316] = 9'b111111111;
assign micromatrizz[19][317] = 9'b111111111;
assign micromatrizz[19][318] = 9'b111111111;
assign micromatrizz[19][319] = 9'b111111111;
assign micromatrizz[19][320] = 9'b111111111;
assign micromatrizz[19][321] = 9'b111111111;
assign micromatrizz[19][322] = 9'b111111111;
assign micromatrizz[19][323] = 9'b111111111;
assign micromatrizz[19][324] = 9'b111111111;
assign micromatrizz[19][325] = 9'b111111111;
assign micromatrizz[19][326] = 9'b111111111;
assign micromatrizz[19][327] = 9'b111111111;
assign micromatrizz[19][328] = 9'b111111111;
assign micromatrizz[19][329] = 9'b111111111;
assign micromatrizz[19][330] = 9'b111111111;
assign micromatrizz[19][331] = 9'b111111111;
assign micromatrizz[19][332] = 9'b111111111;
assign micromatrizz[19][333] = 9'b111111111;
assign micromatrizz[19][334] = 9'b111111111;
assign micromatrizz[19][335] = 9'b111111111;
assign micromatrizz[19][336] = 9'b111111111;
assign micromatrizz[19][337] = 9'b111111111;
assign micromatrizz[19][338] = 9'b111111111;
assign micromatrizz[19][339] = 9'b111111111;
assign micromatrizz[19][340] = 9'b111111111;
assign micromatrizz[19][341] = 9'b111111111;
assign micromatrizz[19][342] = 9'b111111111;
assign micromatrizz[19][343] = 9'b111111111;
assign micromatrizz[19][344] = 9'b111111111;
assign micromatrizz[19][345] = 9'b111111111;
assign micromatrizz[19][346] = 9'b111111111;
assign micromatrizz[19][347] = 9'b111111111;
assign micromatrizz[19][348] = 9'b111111111;
assign micromatrizz[19][349] = 9'b111111111;
assign micromatrizz[19][350] = 9'b111111111;
assign micromatrizz[19][351] = 9'b111111111;
assign micromatrizz[19][352] = 9'b111111111;
assign micromatrizz[19][353] = 9'b111111111;
assign micromatrizz[19][354] = 9'b111111111;
assign micromatrizz[19][355] = 9'b111111111;
assign micromatrizz[19][356] = 9'b111111111;
assign micromatrizz[19][357] = 9'b111111111;
assign micromatrizz[19][358] = 9'b111111111;
assign micromatrizz[19][359] = 9'b111111111;
assign micromatrizz[19][360] = 9'b111111111;
assign micromatrizz[19][361] = 9'b111111111;
assign micromatrizz[19][362] = 9'b111111111;
assign micromatrizz[19][363] = 9'b111111111;
assign micromatrizz[19][364] = 9'b111111111;
assign micromatrizz[19][365] = 9'b111111111;
assign micromatrizz[19][366] = 9'b111111111;
assign micromatrizz[19][367] = 9'b111111111;
assign micromatrizz[19][368] = 9'b111111111;
assign micromatrizz[19][369] = 9'b111111111;
assign micromatrizz[19][370] = 9'b111111111;
assign micromatrizz[19][371] = 9'b111111111;
assign micromatrizz[19][372] = 9'b111111111;
assign micromatrizz[19][373] = 9'b111111111;
assign micromatrizz[19][374] = 9'b111111111;
assign micromatrizz[19][375] = 9'b111111111;
assign micromatrizz[19][376] = 9'b111111111;
assign micromatrizz[19][377] = 9'b111111111;
assign micromatrizz[19][378] = 9'b111111111;
assign micromatrizz[19][379] = 9'b111111111;
assign micromatrizz[19][380] = 9'b111111111;
assign micromatrizz[19][381] = 9'b111111111;
assign micromatrizz[19][382] = 9'b111111111;
assign micromatrizz[19][383] = 9'b111111111;
assign micromatrizz[19][384] = 9'b111111111;
assign micromatrizz[19][385] = 9'b111111111;
assign micromatrizz[19][386] = 9'b111111111;
assign micromatrizz[19][387] = 9'b111111111;
assign micromatrizz[19][388] = 9'b111111111;
assign micromatrizz[19][389] = 9'b111111111;
assign micromatrizz[19][390] = 9'b111111111;
assign micromatrizz[19][391] = 9'b111111111;
assign micromatrizz[19][392] = 9'b111111111;
assign micromatrizz[19][393] = 9'b111111111;
assign micromatrizz[19][394] = 9'b111111111;
assign micromatrizz[19][395] = 9'b111111111;
assign micromatrizz[19][396] = 9'b111111111;
assign micromatrizz[19][397] = 9'b111111111;
assign micromatrizz[19][398] = 9'b111111111;
assign micromatrizz[19][399] = 9'b111111111;
assign micromatrizz[19][400] = 9'b111111111;
assign micromatrizz[19][401] = 9'b111111111;
assign micromatrizz[19][402] = 9'b111111111;
assign micromatrizz[19][403] = 9'b111111111;
assign micromatrizz[19][404] = 9'b111111111;
assign micromatrizz[19][405] = 9'b111111111;
assign micromatrizz[19][406] = 9'b111111111;
assign micromatrizz[19][407] = 9'b111111111;
assign micromatrizz[19][408] = 9'b111111111;
assign micromatrizz[19][409] = 9'b111111111;
assign micromatrizz[19][410] = 9'b111111111;
assign micromatrizz[19][411] = 9'b111111111;
assign micromatrizz[19][412] = 9'b111111111;
assign micromatrizz[19][413] = 9'b111111111;
assign micromatrizz[19][414] = 9'b111111111;
assign micromatrizz[19][415] = 9'b111111111;
assign micromatrizz[19][416] = 9'b111111111;
assign micromatrizz[19][417] = 9'b111111111;
assign micromatrizz[19][418] = 9'b111111111;
assign micromatrizz[19][419] = 9'b111111111;
assign micromatrizz[19][420] = 9'b111111111;
assign micromatrizz[19][421] = 9'b111111111;
assign micromatrizz[19][422] = 9'b111111111;
assign micromatrizz[19][423] = 9'b111111111;
assign micromatrizz[19][424] = 9'b111111111;
assign micromatrizz[19][425] = 9'b111111111;
assign micromatrizz[19][426] = 9'b111111111;
assign micromatrizz[19][427] = 9'b111111111;
assign micromatrizz[19][428] = 9'b111111111;
assign micromatrizz[19][429] = 9'b111111111;
assign micromatrizz[19][430] = 9'b111111111;
assign micromatrizz[19][431] = 9'b111111111;
assign micromatrizz[19][432] = 9'b111111111;
assign micromatrizz[19][433] = 9'b111111111;
assign micromatrizz[19][434] = 9'b111111111;
assign micromatrizz[19][435] = 9'b111111111;
assign micromatrizz[19][436] = 9'b111111111;
assign micromatrizz[19][437] = 9'b111111111;
assign micromatrizz[19][438] = 9'b111111111;
assign micromatrizz[19][439] = 9'b111111111;
assign micromatrizz[19][440] = 9'b111111111;
assign micromatrizz[19][441] = 9'b111111111;
assign micromatrizz[19][442] = 9'b111111111;
assign micromatrizz[19][443] = 9'b111111111;
assign micromatrizz[19][444] = 9'b111111111;
assign micromatrizz[19][445] = 9'b111111111;
assign micromatrizz[19][446] = 9'b111111111;
assign micromatrizz[19][447] = 9'b111111111;
assign micromatrizz[19][448] = 9'b111111111;
assign micromatrizz[19][449] = 9'b111111111;
assign micromatrizz[19][450] = 9'b111111111;
assign micromatrizz[19][451] = 9'b111111111;
assign micromatrizz[19][452] = 9'b111111111;
assign micromatrizz[19][453] = 9'b111111111;
assign micromatrizz[19][454] = 9'b111111111;
assign micromatrizz[19][455] = 9'b111111111;
assign micromatrizz[19][456] = 9'b111111111;
assign micromatrizz[19][457] = 9'b111111111;
assign micromatrizz[19][458] = 9'b111111111;
assign micromatrizz[19][459] = 9'b111111111;
assign micromatrizz[19][460] = 9'b111111111;
assign micromatrizz[19][461] = 9'b111111111;
assign micromatrizz[19][462] = 9'b111111111;
assign micromatrizz[19][463] = 9'b111111111;
assign micromatrizz[19][464] = 9'b111111111;
assign micromatrizz[19][465] = 9'b111111111;
assign micromatrizz[19][466] = 9'b111111111;
assign micromatrizz[19][467] = 9'b111111111;
assign micromatrizz[19][468] = 9'b111111111;
assign micromatrizz[19][469] = 9'b111111111;
assign micromatrizz[19][470] = 9'b111111111;
assign micromatrizz[19][471] = 9'b111111111;
assign micromatrizz[19][472] = 9'b111111111;
assign micromatrizz[19][473] = 9'b111111111;
assign micromatrizz[19][474] = 9'b111111111;
assign micromatrizz[19][475] = 9'b111111111;
assign micromatrizz[19][476] = 9'b111111111;
assign micromatrizz[19][477] = 9'b111111111;
assign micromatrizz[19][478] = 9'b111111111;
assign micromatrizz[19][479] = 9'b111111111;
assign micromatrizz[19][480] = 9'b111111111;
assign micromatrizz[19][481] = 9'b111111111;
assign micromatrizz[19][482] = 9'b111111111;
assign micromatrizz[19][483] = 9'b111111111;
assign micromatrizz[19][484] = 9'b111111111;
assign micromatrizz[19][485] = 9'b111111111;
assign micromatrizz[19][486] = 9'b111111111;
assign micromatrizz[19][487] = 9'b111111111;
assign micromatrizz[19][488] = 9'b111111111;
assign micromatrizz[19][489] = 9'b111111111;
assign micromatrizz[19][490] = 9'b111111111;
assign micromatrizz[19][491] = 9'b111111111;
assign micromatrizz[19][492] = 9'b111111111;
assign micromatrizz[19][493] = 9'b111111111;
assign micromatrizz[19][494] = 9'b111111111;
assign micromatrizz[19][495] = 9'b111111111;
assign micromatrizz[19][496] = 9'b111111111;
assign micromatrizz[19][497] = 9'b111111111;
assign micromatrizz[19][498] = 9'b111111111;
assign micromatrizz[19][499] = 9'b111111111;
assign micromatrizz[19][500] = 9'b111111111;
assign micromatrizz[19][501] = 9'b111111111;
assign micromatrizz[19][502] = 9'b111111111;
assign micromatrizz[19][503] = 9'b111111111;
assign micromatrizz[19][504] = 9'b111111111;
assign micromatrizz[19][505] = 9'b111111111;
assign micromatrizz[19][506] = 9'b111111111;
assign micromatrizz[19][507] = 9'b111111111;
assign micromatrizz[19][508] = 9'b111111111;
assign micromatrizz[19][509] = 9'b111111111;
assign micromatrizz[19][510] = 9'b111111111;
assign micromatrizz[19][511] = 9'b111111111;
assign micromatrizz[19][512] = 9'b111111111;
assign micromatrizz[19][513] = 9'b111111111;
assign micromatrizz[19][514] = 9'b111111111;
assign micromatrizz[19][515] = 9'b111111111;
assign micromatrizz[19][516] = 9'b111111111;
assign micromatrizz[19][517] = 9'b111111111;
assign micromatrizz[19][518] = 9'b111111111;
assign micromatrizz[19][519] = 9'b111111111;
assign micromatrizz[19][520] = 9'b111111111;
assign micromatrizz[19][521] = 9'b111111111;
assign micromatrizz[19][522] = 9'b111111111;
assign micromatrizz[19][523] = 9'b111111111;
assign micromatrizz[19][524] = 9'b111111111;
assign micromatrizz[19][525] = 9'b111111111;
assign micromatrizz[19][526] = 9'b111111111;
assign micromatrizz[19][527] = 9'b111111111;
assign micromatrizz[19][528] = 9'b111111111;
assign micromatrizz[19][529] = 9'b111111111;
assign micromatrizz[19][530] = 9'b111111111;
assign micromatrizz[19][531] = 9'b111111111;
assign micromatrizz[19][532] = 9'b111111111;
assign micromatrizz[19][533] = 9'b111111111;
assign micromatrizz[19][534] = 9'b111111111;
assign micromatrizz[19][535] = 9'b111111111;
assign micromatrizz[19][536] = 9'b111111111;
assign micromatrizz[19][537] = 9'b111111111;
assign micromatrizz[19][538] = 9'b111111111;
assign micromatrizz[19][539] = 9'b111111111;
assign micromatrizz[19][540] = 9'b111111111;
assign micromatrizz[19][541] = 9'b111111111;
assign micromatrizz[19][542] = 9'b111111111;
assign micromatrizz[19][543] = 9'b111111111;
assign micromatrizz[19][544] = 9'b111111111;
assign micromatrizz[19][545] = 9'b111111111;
assign micromatrizz[19][546] = 9'b111111111;
assign micromatrizz[19][547] = 9'b111111111;
assign micromatrizz[19][548] = 9'b111111111;
assign micromatrizz[19][549] = 9'b111111111;
assign micromatrizz[19][550] = 9'b111111111;
assign micromatrizz[19][551] = 9'b111111111;
assign micromatrizz[19][552] = 9'b111111111;
assign micromatrizz[19][553] = 9'b111111111;
assign micromatrizz[19][554] = 9'b111111111;
assign micromatrizz[19][555] = 9'b111111111;
assign micromatrizz[19][556] = 9'b111111111;
assign micromatrizz[19][557] = 9'b111111111;
assign micromatrizz[19][558] = 9'b111111111;
assign micromatrizz[19][559] = 9'b111111111;
assign micromatrizz[19][560] = 9'b111111111;
assign micromatrizz[19][561] = 9'b111111111;
assign micromatrizz[19][562] = 9'b111111111;
assign micromatrizz[19][563] = 9'b111111111;
assign micromatrizz[19][564] = 9'b111111111;
assign micromatrizz[19][565] = 9'b111111111;
assign micromatrizz[19][566] = 9'b111111111;
assign micromatrizz[19][567] = 9'b111111111;
assign micromatrizz[19][568] = 9'b111111111;
assign micromatrizz[19][569] = 9'b111111111;
assign micromatrizz[19][570] = 9'b111111111;
assign micromatrizz[19][571] = 9'b111111111;
assign micromatrizz[19][572] = 9'b111111111;
assign micromatrizz[19][573] = 9'b111111111;
assign micromatrizz[19][574] = 9'b111111111;
assign micromatrizz[19][575] = 9'b111111111;
assign micromatrizz[19][576] = 9'b111111111;
assign micromatrizz[19][577] = 9'b111111111;
assign micromatrizz[19][578] = 9'b111111111;
assign micromatrizz[19][579] = 9'b111111111;
assign micromatrizz[19][580] = 9'b111111111;
assign micromatrizz[19][581] = 9'b111111111;
assign micromatrizz[19][582] = 9'b111111111;
assign micromatrizz[19][583] = 9'b111111111;
assign micromatrizz[19][584] = 9'b111111111;
assign micromatrizz[19][585] = 9'b111111111;
assign micromatrizz[19][586] = 9'b111111111;
assign micromatrizz[19][587] = 9'b111111111;
assign micromatrizz[19][588] = 9'b111111111;
assign micromatrizz[19][589] = 9'b111111111;
assign micromatrizz[19][590] = 9'b111111111;
assign micromatrizz[19][591] = 9'b111111111;
assign micromatrizz[19][592] = 9'b111111111;
assign micromatrizz[19][593] = 9'b111111111;
assign micromatrizz[19][594] = 9'b111111111;
assign micromatrizz[19][595] = 9'b111111111;
assign micromatrizz[19][596] = 9'b111111111;
assign micromatrizz[19][597] = 9'b111111111;
assign micromatrizz[19][598] = 9'b111111111;
assign micromatrizz[19][599] = 9'b111111111;
assign micromatrizz[19][600] = 9'b111111111;
assign micromatrizz[19][601] = 9'b111111111;
assign micromatrizz[19][602] = 9'b111111111;
assign micromatrizz[19][603] = 9'b111111111;
assign micromatrizz[19][604] = 9'b111111111;
assign micromatrizz[19][605] = 9'b111111111;
assign micromatrizz[19][606] = 9'b111111111;
assign micromatrizz[19][607] = 9'b111111111;
assign micromatrizz[19][608] = 9'b111111111;
assign micromatrizz[19][609] = 9'b111111111;
assign micromatrizz[19][610] = 9'b111111111;
assign micromatrizz[19][611] = 9'b111111111;
assign micromatrizz[19][612] = 9'b111111111;
assign micromatrizz[19][613] = 9'b111111111;
assign micromatrizz[19][614] = 9'b111111111;
assign micromatrizz[19][615] = 9'b111111111;
assign micromatrizz[19][616] = 9'b111111111;
assign micromatrizz[19][617] = 9'b111111111;
assign micromatrizz[19][618] = 9'b111111111;
assign micromatrizz[19][619] = 9'b111111111;
assign micromatrizz[19][620] = 9'b111111111;
assign micromatrizz[19][621] = 9'b111111111;
assign micromatrizz[19][622] = 9'b111111111;
assign micromatrizz[19][623] = 9'b111111111;
assign micromatrizz[19][624] = 9'b111111111;
assign micromatrizz[19][625] = 9'b111111111;
assign micromatrizz[19][626] = 9'b111111111;
assign micromatrizz[19][627] = 9'b111111111;
assign micromatrizz[19][628] = 9'b111111111;
assign micromatrizz[19][629] = 9'b111111111;
assign micromatrizz[19][630] = 9'b111111111;
assign micromatrizz[19][631] = 9'b111111111;
assign micromatrizz[19][632] = 9'b111111111;
assign micromatrizz[19][633] = 9'b111111111;
assign micromatrizz[19][634] = 9'b111111111;
assign micromatrizz[19][635] = 9'b111111111;
assign micromatrizz[19][636] = 9'b111111111;
assign micromatrizz[19][637] = 9'b111111111;
assign micromatrizz[19][638] = 9'b111111111;
assign micromatrizz[19][639] = 9'b111111111;
assign micromatrizz[20][0] = 9'b111111111;
assign micromatrizz[20][1] = 9'b111111111;
assign micromatrizz[20][2] = 9'b111111111;
assign micromatrizz[20][3] = 9'b111111111;
assign micromatrizz[20][4] = 9'b111111111;
assign micromatrizz[20][5] = 9'b111111111;
assign micromatrizz[20][6] = 9'b111111111;
assign micromatrizz[20][7] = 9'b111111111;
assign micromatrizz[20][8] = 9'b111111111;
assign micromatrizz[20][9] = 9'b111111111;
assign micromatrizz[20][10] = 9'b111111111;
assign micromatrizz[20][11] = 9'b111111111;
assign micromatrizz[20][12] = 9'b111111111;
assign micromatrizz[20][13] = 9'b111111111;
assign micromatrizz[20][14] = 9'b111111111;
assign micromatrizz[20][15] = 9'b111111111;
assign micromatrizz[20][16] = 9'b111111111;
assign micromatrizz[20][17] = 9'b111111111;
assign micromatrizz[20][18] = 9'b111111111;
assign micromatrizz[20][19] = 9'b111111111;
assign micromatrizz[20][20] = 9'b111111111;
assign micromatrizz[20][21] = 9'b111111111;
assign micromatrizz[20][22] = 9'b111111111;
assign micromatrizz[20][23] = 9'b111111111;
assign micromatrizz[20][24] = 9'b111111111;
assign micromatrizz[20][25] = 9'b111111111;
assign micromatrizz[20][26] = 9'b111111111;
assign micromatrizz[20][27] = 9'b111111111;
assign micromatrizz[20][28] = 9'b111111111;
assign micromatrizz[20][29] = 9'b111111111;
assign micromatrizz[20][30] = 9'b111111111;
assign micromatrizz[20][31] = 9'b111111111;
assign micromatrizz[20][32] = 9'b111111111;
assign micromatrizz[20][33] = 9'b111111111;
assign micromatrizz[20][34] = 9'b111111111;
assign micromatrizz[20][35] = 9'b111111111;
assign micromatrizz[20][36] = 9'b111111111;
assign micromatrizz[20][37] = 9'b111111111;
assign micromatrizz[20][38] = 9'b111111111;
assign micromatrizz[20][39] = 9'b111111111;
assign micromatrizz[20][40] = 9'b111111111;
assign micromatrizz[20][41] = 9'b111111111;
assign micromatrizz[20][42] = 9'b111111111;
assign micromatrizz[20][43] = 9'b111111111;
assign micromatrizz[20][44] = 9'b111111111;
assign micromatrizz[20][45] = 9'b111111111;
assign micromatrizz[20][46] = 9'b111111111;
assign micromatrizz[20][47] = 9'b111111111;
assign micromatrizz[20][48] = 9'b111111111;
assign micromatrizz[20][49] = 9'b111111111;
assign micromatrizz[20][50] = 9'b111111111;
assign micromatrizz[20][51] = 9'b111111111;
assign micromatrizz[20][52] = 9'b111111111;
assign micromatrizz[20][53] = 9'b111111111;
assign micromatrizz[20][54] = 9'b111111111;
assign micromatrizz[20][55] = 9'b111111111;
assign micromatrizz[20][56] = 9'b111111111;
assign micromatrizz[20][57] = 9'b111111111;
assign micromatrizz[20][58] = 9'b111111111;
assign micromatrizz[20][59] = 9'b111111111;
assign micromatrizz[20][60] = 9'b111111111;
assign micromatrizz[20][61] = 9'b111111111;
assign micromatrizz[20][62] = 9'b111111111;
assign micromatrizz[20][63] = 9'b111111111;
assign micromatrizz[20][64] = 9'b111111111;
assign micromatrizz[20][65] = 9'b111111111;
assign micromatrizz[20][66] = 9'b111111111;
assign micromatrizz[20][67] = 9'b111111111;
assign micromatrizz[20][68] = 9'b111111111;
assign micromatrizz[20][69] = 9'b111111111;
assign micromatrizz[20][70] = 9'b111111111;
assign micromatrizz[20][71] = 9'b111111111;
assign micromatrizz[20][72] = 9'b111111111;
assign micromatrizz[20][73] = 9'b111111111;
assign micromatrizz[20][74] = 9'b111111111;
assign micromatrizz[20][75] = 9'b111111111;
assign micromatrizz[20][76] = 9'b111111111;
assign micromatrizz[20][77] = 9'b111111111;
assign micromatrizz[20][78] = 9'b111111111;
assign micromatrizz[20][79] = 9'b111111111;
assign micromatrizz[20][80] = 9'b111111111;
assign micromatrizz[20][81] = 9'b111111111;
assign micromatrizz[20][82] = 9'b111111111;
assign micromatrizz[20][83] = 9'b111111111;
assign micromatrizz[20][84] = 9'b111111111;
assign micromatrizz[20][85] = 9'b111111111;
assign micromatrizz[20][86] = 9'b111111111;
assign micromatrizz[20][87] = 9'b111111111;
assign micromatrizz[20][88] = 9'b111111111;
assign micromatrizz[20][89] = 9'b111111111;
assign micromatrizz[20][90] = 9'b111111111;
assign micromatrizz[20][91] = 9'b111111111;
assign micromatrizz[20][92] = 9'b111111111;
assign micromatrizz[20][93] = 9'b111111111;
assign micromatrizz[20][94] = 9'b111111111;
assign micromatrizz[20][95] = 9'b111111111;
assign micromatrizz[20][96] = 9'b111111111;
assign micromatrizz[20][97] = 9'b111111111;
assign micromatrizz[20][98] = 9'b111111111;
assign micromatrizz[20][99] = 9'b111111111;
assign micromatrizz[20][100] = 9'b111111111;
assign micromatrizz[20][101] = 9'b111111111;
assign micromatrizz[20][102] = 9'b111111111;
assign micromatrizz[20][103] = 9'b111111111;
assign micromatrizz[20][104] = 9'b111111111;
assign micromatrizz[20][105] = 9'b111111111;
assign micromatrizz[20][106] = 9'b111111111;
assign micromatrizz[20][107] = 9'b111111111;
assign micromatrizz[20][108] = 9'b111111111;
assign micromatrizz[20][109] = 9'b111111111;
assign micromatrizz[20][110] = 9'b111111111;
assign micromatrizz[20][111] = 9'b111111111;
assign micromatrizz[20][112] = 9'b111111111;
assign micromatrizz[20][113] = 9'b111111111;
assign micromatrizz[20][114] = 9'b111111111;
assign micromatrizz[20][115] = 9'b111111111;
assign micromatrizz[20][116] = 9'b111111111;
assign micromatrizz[20][117] = 9'b111111111;
assign micromatrizz[20][118] = 9'b111111111;
assign micromatrizz[20][119] = 9'b111111111;
assign micromatrizz[20][120] = 9'b111111111;
assign micromatrizz[20][121] = 9'b111111111;
assign micromatrizz[20][122] = 9'b111111111;
assign micromatrizz[20][123] = 9'b111111111;
assign micromatrizz[20][124] = 9'b111111111;
assign micromatrizz[20][125] = 9'b111111111;
assign micromatrizz[20][126] = 9'b111111111;
assign micromatrizz[20][127] = 9'b111111111;
assign micromatrizz[20][128] = 9'b111111111;
assign micromatrizz[20][129] = 9'b111111111;
assign micromatrizz[20][130] = 9'b111111111;
assign micromatrizz[20][131] = 9'b111111111;
assign micromatrizz[20][132] = 9'b111111111;
assign micromatrizz[20][133] = 9'b111111111;
assign micromatrizz[20][134] = 9'b111111111;
assign micromatrizz[20][135] = 9'b111111111;
assign micromatrizz[20][136] = 9'b111111111;
assign micromatrizz[20][137] = 9'b111111111;
assign micromatrizz[20][138] = 9'b111111111;
assign micromatrizz[20][139] = 9'b111111111;
assign micromatrizz[20][140] = 9'b111111111;
assign micromatrizz[20][141] = 9'b111111111;
assign micromatrizz[20][142] = 9'b111111111;
assign micromatrizz[20][143] = 9'b111111111;
assign micromatrizz[20][144] = 9'b111111111;
assign micromatrizz[20][145] = 9'b111111111;
assign micromatrizz[20][146] = 9'b111111111;
assign micromatrizz[20][147] = 9'b111111111;
assign micromatrizz[20][148] = 9'b111111111;
assign micromatrizz[20][149] = 9'b111111111;
assign micromatrizz[20][150] = 9'b111111111;
assign micromatrizz[20][151] = 9'b111111111;
assign micromatrizz[20][152] = 9'b111111111;
assign micromatrizz[20][153] = 9'b111111111;
assign micromatrizz[20][154] = 9'b111111111;
assign micromatrizz[20][155] = 9'b111111111;
assign micromatrizz[20][156] = 9'b111111111;
assign micromatrizz[20][157] = 9'b111111111;
assign micromatrizz[20][158] = 9'b111111111;
assign micromatrizz[20][159] = 9'b111111111;
assign micromatrizz[20][160] = 9'b111111111;
assign micromatrizz[20][161] = 9'b111111111;
assign micromatrizz[20][162] = 9'b111111111;
assign micromatrizz[20][163] = 9'b111111111;
assign micromatrizz[20][164] = 9'b111111111;
assign micromatrizz[20][165] = 9'b111111111;
assign micromatrizz[20][166] = 9'b111111111;
assign micromatrizz[20][167] = 9'b111111111;
assign micromatrizz[20][168] = 9'b111111111;
assign micromatrizz[20][169] = 9'b111111111;
assign micromatrizz[20][170] = 9'b111111111;
assign micromatrizz[20][171] = 9'b111111111;
assign micromatrizz[20][172] = 9'b111111111;
assign micromatrizz[20][173] = 9'b111111111;
assign micromatrizz[20][174] = 9'b111111111;
assign micromatrizz[20][175] = 9'b111111111;
assign micromatrizz[20][176] = 9'b111111111;
assign micromatrizz[20][177] = 9'b111111111;
assign micromatrizz[20][178] = 9'b111111111;
assign micromatrizz[20][179] = 9'b111111111;
assign micromatrizz[20][180] = 9'b111111111;
assign micromatrizz[20][181] = 9'b111111111;
assign micromatrizz[20][182] = 9'b111111111;
assign micromatrizz[20][183] = 9'b111111111;
assign micromatrizz[20][184] = 9'b111111111;
assign micromatrizz[20][185] = 9'b111111111;
assign micromatrizz[20][186] = 9'b111111111;
assign micromatrizz[20][187] = 9'b111111111;
assign micromatrizz[20][188] = 9'b111111111;
assign micromatrizz[20][189] = 9'b111111111;
assign micromatrizz[20][190] = 9'b111111111;
assign micromatrizz[20][191] = 9'b111111111;
assign micromatrizz[20][192] = 9'b111111111;
assign micromatrizz[20][193] = 9'b111111111;
assign micromatrizz[20][194] = 9'b111111111;
assign micromatrizz[20][195] = 9'b111111111;
assign micromatrizz[20][196] = 9'b111111111;
assign micromatrizz[20][197] = 9'b111111111;
assign micromatrizz[20][198] = 9'b111111111;
assign micromatrizz[20][199] = 9'b111111111;
assign micromatrizz[20][200] = 9'b111111111;
assign micromatrizz[20][201] = 9'b111111111;
assign micromatrizz[20][202] = 9'b111111111;
assign micromatrizz[20][203] = 9'b111111111;
assign micromatrizz[20][204] = 9'b111111111;
assign micromatrizz[20][205] = 9'b111111111;
assign micromatrizz[20][206] = 9'b111111111;
assign micromatrizz[20][207] = 9'b111111111;
assign micromatrizz[20][208] = 9'b111111111;
assign micromatrizz[20][209] = 9'b111111111;
assign micromatrizz[20][210] = 9'b111111111;
assign micromatrizz[20][211] = 9'b111111111;
assign micromatrizz[20][212] = 9'b111111111;
assign micromatrizz[20][213] = 9'b111111111;
assign micromatrizz[20][214] = 9'b111111111;
assign micromatrizz[20][215] = 9'b111111111;
assign micromatrizz[20][216] = 9'b111111111;
assign micromatrizz[20][217] = 9'b111111111;
assign micromatrizz[20][218] = 9'b111111111;
assign micromatrizz[20][219] = 9'b111111111;
assign micromatrizz[20][220] = 9'b111111111;
assign micromatrizz[20][221] = 9'b111111111;
assign micromatrizz[20][222] = 9'b111111111;
assign micromatrizz[20][223] = 9'b111111111;
assign micromatrizz[20][224] = 9'b111111111;
assign micromatrizz[20][225] = 9'b111111111;
assign micromatrizz[20][226] = 9'b111111111;
assign micromatrizz[20][227] = 9'b111111111;
assign micromatrizz[20][228] = 9'b111111111;
assign micromatrizz[20][229] = 9'b111111111;
assign micromatrizz[20][230] = 9'b111111111;
assign micromatrizz[20][231] = 9'b111111111;
assign micromatrizz[20][232] = 9'b111111111;
assign micromatrizz[20][233] = 9'b111111111;
assign micromatrizz[20][234] = 9'b111111111;
assign micromatrizz[20][235] = 9'b111111111;
assign micromatrizz[20][236] = 9'b111111111;
assign micromatrizz[20][237] = 9'b111111111;
assign micromatrizz[20][238] = 9'b111111111;
assign micromatrizz[20][239] = 9'b111111111;
assign micromatrizz[20][240] = 9'b111111111;
assign micromatrizz[20][241] = 9'b111111111;
assign micromatrizz[20][242] = 9'b111111111;
assign micromatrizz[20][243] = 9'b111111111;
assign micromatrizz[20][244] = 9'b111111111;
assign micromatrizz[20][245] = 9'b111111111;
assign micromatrizz[20][246] = 9'b111111111;
assign micromatrizz[20][247] = 9'b111111111;
assign micromatrizz[20][248] = 9'b111111111;
assign micromatrizz[20][249] = 9'b111111111;
assign micromatrizz[20][250] = 9'b111111111;
assign micromatrizz[20][251] = 9'b111111111;
assign micromatrizz[20][252] = 9'b111111111;
assign micromatrizz[20][253] = 9'b111111111;
assign micromatrizz[20][254] = 9'b111111111;
assign micromatrizz[20][255] = 9'b111111111;
assign micromatrizz[20][256] = 9'b111111111;
assign micromatrizz[20][257] = 9'b111111111;
assign micromatrizz[20][258] = 9'b111111111;
assign micromatrizz[20][259] = 9'b111111111;
assign micromatrizz[20][260] = 9'b111111111;
assign micromatrizz[20][261] = 9'b111111111;
assign micromatrizz[20][262] = 9'b111111111;
assign micromatrizz[20][263] = 9'b111111111;
assign micromatrizz[20][264] = 9'b111111111;
assign micromatrizz[20][265] = 9'b111111111;
assign micromatrizz[20][266] = 9'b111111111;
assign micromatrizz[20][267] = 9'b111111111;
assign micromatrizz[20][268] = 9'b111111111;
assign micromatrizz[20][269] = 9'b111111111;
assign micromatrizz[20][270] = 9'b111110010;
assign micromatrizz[20][271] = 9'b111110010;
assign micromatrizz[20][272] = 9'b111110010;
assign micromatrizz[20][273] = 9'b111110010;
assign micromatrizz[20][274] = 9'b111110010;
assign micromatrizz[20][275] = 9'b111110011;
assign micromatrizz[20][276] = 9'b111110011;
assign micromatrizz[20][277] = 9'b111110011;
assign micromatrizz[20][278] = 9'b111110011;
assign micromatrizz[20][279] = 9'b111111111;
assign micromatrizz[20][280] = 9'b111111111;
assign micromatrizz[20][281] = 9'b111111111;
assign micromatrizz[20][282] = 9'b111111111;
assign micromatrizz[20][283] = 9'b111111111;
assign micromatrizz[20][284] = 9'b111111111;
assign micromatrizz[20][285] = 9'b111111111;
assign micromatrizz[20][286] = 9'b111111111;
assign micromatrizz[20][287] = 9'b111111111;
assign micromatrizz[20][288] = 9'b111111111;
assign micromatrizz[20][289] = 9'b111111111;
assign micromatrizz[20][290] = 9'b111111111;
assign micromatrizz[20][291] = 9'b111111111;
assign micromatrizz[20][292] = 9'b111111111;
assign micromatrizz[20][293] = 9'b111111111;
assign micromatrizz[20][294] = 9'b111111111;
assign micromatrizz[20][295] = 9'b111111111;
assign micromatrizz[20][296] = 9'b111111111;
assign micromatrizz[20][297] = 9'b111111111;
assign micromatrizz[20][298] = 9'b111111111;
assign micromatrizz[20][299] = 9'b111111111;
assign micromatrizz[20][300] = 9'b111111111;
assign micromatrizz[20][301] = 9'b111111111;
assign micromatrizz[20][302] = 9'b111111111;
assign micromatrizz[20][303] = 9'b111111111;
assign micromatrizz[20][304] = 9'b111111111;
assign micromatrizz[20][305] = 9'b111111111;
assign micromatrizz[20][306] = 9'b111111111;
assign micromatrizz[20][307] = 9'b111111111;
assign micromatrizz[20][308] = 9'b111111111;
assign micromatrizz[20][309] = 9'b111111111;
assign micromatrizz[20][310] = 9'b111111111;
assign micromatrizz[20][311] = 9'b111111111;
assign micromatrizz[20][312] = 9'b111111111;
assign micromatrizz[20][313] = 9'b111111111;
assign micromatrizz[20][314] = 9'b111111111;
assign micromatrizz[20][315] = 9'b111111111;
assign micromatrizz[20][316] = 9'b111111111;
assign micromatrizz[20][317] = 9'b111111111;
assign micromatrizz[20][318] = 9'b111111111;
assign micromatrizz[20][319] = 9'b111111111;
assign micromatrizz[20][320] = 9'b111111111;
assign micromatrizz[20][321] = 9'b111111111;
assign micromatrizz[20][322] = 9'b111111111;
assign micromatrizz[20][323] = 9'b111111111;
assign micromatrizz[20][324] = 9'b111111111;
assign micromatrizz[20][325] = 9'b111111111;
assign micromatrizz[20][326] = 9'b111111111;
assign micromatrizz[20][327] = 9'b111111111;
assign micromatrizz[20][328] = 9'b111111111;
assign micromatrizz[20][329] = 9'b111111111;
assign micromatrizz[20][330] = 9'b111111111;
assign micromatrizz[20][331] = 9'b111111111;
assign micromatrizz[20][332] = 9'b111111111;
assign micromatrizz[20][333] = 9'b111111111;
assign micromatrizz[20][334] = 9'b111111111;
assign micromatrizz[20][335] = 9'b111111111;
assign micromatrizz[20][336] = 9'b111111111;
assign micromatrizz[20][337] = 9'b111111111;
assign micromatrizz[20][338] = 9'b111111111;
assign micromatrizz[20][339] = 9'b111111111;
assign micromatrizz[20][340] = 9'b111111111;
assign micromatrizz[20][341] = 9'b111111111;
assign micromatrizz[20][342] = 9'b111111111;
assign micromatrizz[20][343] = 9'b111111111;
assign micromatrizz[20][344] = 9'b111111111;
assign micromatrizz[20][345] = 9'b111111111;
assign micromatrizz[20][346] = 9'b111111111;
assign micromatrizz[20][347] = 9'b111111111;
assign micromatrizz[20][348] = 9'b111111111;
assign micromatrizz[20][349] = 9'b111111111;
assign micromatrizz[20][350] = 9'b111111111;
assign micromatrizz[20][351] = 9'b111111111;
assign micromatrizz[20][352] = 9'b111111111;
assign micromatrizz[20][353] = 9'b111111111;
assign micromatrizz[20][354] = 9'b111111111;
assign micromatrizz[20][355] = 9'b111111111;
assign micromatrizz[20][356] = 9'b111111111;
assign micromatrizz[20][357] = 9'b111111111;
assign micromatrizz[20][358] = 9'b111111111;
assign micromatrizz[20][359] = 9'b111111111;
assign micromatrizz[20][360] = 9'b111111111;
assign micromatrizz[20][361] = 9'b111111111;
assign micromatrizz[20][362] = 9'b111111111;
assign micromatrizz[20][363] = 9'b111111111;
assign micromatrizz[20][364] = 9'b111111111;
assign micromatrizz[20][365] = 9'b111111111;
assign micromatrizz[20][366] = 9'b111111111;
assign micromatrizz[20][367] = 9'b111111111;
assign micromatrizz[20][368] = 9'b111111111;
assign micromatrizz[20][369] = 9'b111111111;
assign micromatrizz[20][370] = 9'b111111111;
assign micromatrizz[20][371] = 9'b111111111;
assign micromatrizz[20][372] = 9'b111111111;
assign micromatrizz[20][373] = 9'b111111111;
assign micromatrizz[20][374] = 9'b111111111;
assign micromatrizz[20][375] = 9'b111111111;
assign micromatrizz[20][376] = 9'b111111111;
assign micromatrizz[20][377] = 9'b111111111;
assign micromatrizz[20][378] = 9'b111111111;
assign micromatrizz[20][379] = 9'b111111111;
assign micromatrizz[20][380] = 9'b111111111;
assign micromatrizz[20][381] = 9'b111111111;
assign micromatrizz[20][382] = 9'b111111111;
assign micromatrizz[20][383] = 9'b111111111;
assign micromatrizz[20][384] = 9'b111111111;
assign micromatrizz[20][385] = 9'b111111111;
assign micromatrizz[20][386] = 9'b111111111;
assign micromatrizz[20][387] = 9'b111111111;
assign micromatrizz[20][388] = 9'b111111111;
assign micromatrizz[20][389] = 9'b111111111;
assign micromatrizz[20][390] = 9'b111111111;
assign micromatrizz[20][391] = 9'b111111111;
assign micromatrizz[20][392] = 9'b111111111;
assign micromatrizz[20][393] = 9'b111111111;
assign micromatrizz[20][394] = 9'b111111111;
assign micromatrizz[20][395] = 9'b111111111;
assign micromatrizz[20][396] = 9'b111111111;
assign micromatrizz[20][397] = 9'b111111111;
assign micromatrizz[20][398] = 9'b111111111;
assign micromatrizz[20][399] = 9'b111111111;
assign micromatrizz[20][400] = 9'b111111111;
assign micromatrizz[20][401] = 9'b111111111;
assign micromatrizz[20][402] = 9'b111111111;
assign micromatrizz[20][403] = 9'b111111111;
assign micromatrizz[20][404] = 9'b111111111;
assign micromatrizz[20][405] = 9'b111111111;
assign micromatrizz[20][406] = 9'b111111111;
assign micromatrizz[20][407] = 9'b111111111;
assign micromatrizz[20][408] = 9'b111111111;
assign micromatrizz[20][409] = 9'b111111111;
assign micromatrizz[20][410] = 9'b111111111;
assign micromatrizz[20][411] = 9'b111111111;
assign micromatrizz[20][412] = 9'b111111111;
assign micromatrizz[20][413] = 9'b111111111;
assign micromatrizz[20][414] = 9'b111111111;
assign micromatrizz[20][415] = 9'b111111111;
assign micromatrizz[20][416] = 9'b111111111;
assign micromatrizz[20][417] = 9'b111111111;
assign micromatrizz[20][418] = 9'b111111111;
assign micromatrizz[20][419] = 9'b111111111;
assign micromatrizz[20][420] = 9'b111111111;
assign micromatrizz[20][421] = 9'b111111111;
assign micromatrizz[20][422] = 9'b111111111;
assign micromatrizz[20][423] = 9'b111111111;
assign micromatrizz[20][424] = 9'b111111111;
assign micromatrizz[20][425] = 9'b111111111;
assign micromatrizz[20][426] = 9'b111111111;
assign micromatrizz[20][427] = 9'b111111111;
assign micromatrizz[20][428] = 9'b111111111;
assign micromatrizz[20][429] = 9'b111111111;
assign micromatrizz[20][430] = 9'b111111111;
assign micromatrizz[20][431] = 9'b111111111;
assign micromatrizz[20][432] = 9'b111111111;
assign micromatrizz[20][433] = 9'b111111111;
assign micromatrizz[20][434] = 9'b111111111;
assign micromatrizz[20][435] = 9'b111111111;
assign micromatrizz[20][436] = 9'b111111111;
assign micromatrizz[20][437] = 9'b111111111;
assign micromatrizz[20][438] = 9'b111111111;
assign micromatrizz[20][439] = 9'b111111111;
assign micromatrizz[20][440] = 9'b111111111;
assign micromatrizz[20][441] = 9'b111111111;
assign micromatrizz[20][442] = 9'b111111111;
assign micromatrizz[20][443] = 9'b111111111;
assign micromatrizz[20][444] = 9'b111111111;
assign micromatrizz[20][445] = 9'b111111111;
assign micromatrizz[20][446] = 9'b111111111;
assign micromatrizz[20][447] = 9'b111111111;
assign micromatrizz[20][448] = 9'b111111111;
assign micromatrizz[20][449] = 9'b111111111;
assign micromatrizz[20][450] = 9'b111111111;
assign micromatrizz[20][451] = 9'b111111111;
assign micromatrizz[20][452] = 9'b111111111;
assign micromatrizz[20][453] = 9'b111111111;
assign micromatrizz[20][454] = 9'b111111111;
assign micromatrizz[20][455] = 9'b111111111;
assign micromatrizz[20][456] = 9'b111111111;
assign micromatrizz[20][457] = 9'b111111111;
assign micromatrizz[20][458] = 9'b111111111;
assign micromatrizz[20][459] = 9'b111111111;
assign micromatrizz[20][460] = 9'b111111111;
assign micromatrizz[20][461] = 9'b111111111;
assign micromatrizz[20][462] = 9'b111111111;
assign micromatrizz[20][463] = 9'b111111111;
assign micromatrizz[20][464] = 9'b111111111;
assign micromatrizz[20][465] = 9'b111111111;
assign micromatrizz[20][466] = 9'b111111111;
assign micromatrizz[20][467] = 9'b111111111;
assign micromatrizz[20][468] = 9'b111111111;
assign micromatrizz[20][469] = 9'b111111111;
assign micromatrizz[20][470] = 9'b111111111;
assign micromatrizz[20][471] = 9'b111111111;
assign micromatrizz[20][472] = 9'b111111111;
assign micromatrizz[20][473] = 9'b111111111;
assign micromatrizz[20][474] = 9'b111111111;
assign micromatrizz[20][475] = 9'b111111111;
assign micromatrizz[20][476] = 9'b111111111;
assign micromatrizz[20][477] = 9'b111111111;
assign micromatrizz[20][478] = 9'b111111111;
assign micromatrizz[20][479] = 9'b111111111;
assign micromatrizz[20][480] = 9'b111111111;
assign micromatrizz[20][481] = 9'b111111111;
assign micromatrizz[20][482] = 9'b111111111;
assign micromatrizz[20][483] = 9'b111111111;
assign micromatrizz[20][484] = 9'b111111111;
assign micromatrizz[20][485] = 9'b111111111;
assign micromatrizz[20][486] = 9'b111111111;
assign micromatrizz[20][487] = 9'b111111111;
assign micromatrizz[20][488] = 9'b111111111;
assign micromatrizz[20][489] = 9'b111111111;
assign micromatrizz[20][490] = 9'b111111111;
assign micromatrizz[20][491] = 9'b111111111;
assign micromatrizz[20][492] = 9'b111111111;
assign micromatrizz[20][493] = 9'b111111111;
assign micromatrizz[20][494] = 9'b111111111;
assign micromatrizz[20][495] = 9'b111111111;
assign micromatrizz[20][496] = 9'b111111111;
assign micromatrizz[20][497] = 9'b111111111;
assign micromatrizz[20][498] = 9'b111111111;
assign micromatrizz[20][499] = 9'b111111111;
assign micromatrizz[20][500] = 9'b111111111;
assign micromatrizz[20][501] = 9'b111111111;
assign micromatrizz[20][502] = 9'b111111111;
assign micromatrizz[20][503] = 9'b111111111;
assign micromatrizz[20][504] = 9'b111111111;
assign micromatrizz[20][505] = 9'b111111111;
assign micromatrizz[20][506] = 9'b111111111;
assign micromatrizz[20][507] = 9'b111111111;
assign micromatrizz[20][508] = 9'b111111111;
assign micromatrizz[20][509] = 9'b111111111;
assign micromatrizz[20][510] = 9'b111111111;
assign micromatrizz[20][511] = 9'b111111111;
assign micromatrizz[20][512] = 9'b111111111;
assign micromatrizz[20][513] = 9'b111111111;
assign micromatrizz[20][514] = 9'b111111111;
assign micromatrizz[20][515] = 9'b111111111;
assign micromatrizz[20][516] = 9'b111111111;
assign micromatrizz[20][517] = 9'b111111111;
assign micromatrizz[20][518] = 9'b111111111;
assign micromatrizz[20][519] = 9'b111111111;
assign micromatrizz[20][520] = 9'b111111111;
assign micromatrizz[20][521] = 9'b111111111;
assign micromatrizz[20][522] = 9'b111111111;
assign micromatrizz[20][523] = 9'b111111111;
assign micromatrizz[20][524] = 9'b111111111;
assign micromatrizz[20][525] = 9'b111111111;
assign micromatrizz[20][526] = 9'b111111111;
assign micromatrizz[20][527] = 9'b111111111;
assign micromatrizz[20][528] = 9'b111111111;
assign micromatrizz[20][529] = 9'b111111111;
assign micromatrizz[20][530] = 9'b111111111;
assign micromatrizz[20][531] = 9'b111111111;
assign micromatrizz[20][532] = 9'b111111111;
assign micromatrizz[20][533] = 9'b111111111;
assign micromatrizz[20][534] = 9'b111111111;
assign micromatrizz[20][535] = 9'b111111111;
assign micromatrizz[20][536] = 9'b111111111;
assign micromatrizz[20][537] = 9'b111111111;
assign micromatrizz[20][538] = 9'b111111111;
assign micromatrizz[20][539] = 9'b111111111;
assign micromatrizz[20][540] = 9'b111111111;
assign micromatrizz[20][541] = 9'b111111111;
assign micromatrizz[20][542] = 9'b111111111;
assign micromatrizz[20][543] = 9'b111111111;
assign micromatrizz[20][544] = 9'b111111111;
assign micromatrizz[20][545] = 9'b111111111;
assign micromatrizz[20][546] = 9'b111111111;
assign micromatrizz[20][547] = 9'b111111111;
assign micromatrizz[20][548] = 9'b111111111;
assign micromatrizz[20][549] = 9'b111111111;
assign micromatrizz[20][550] = 9'b111111111;
assign micromatrizz[20][551] = 9'b111111111;
assign micromatrizz[20][552] = 9'b111111111;
assign micromatrizz[20][553] = 9'b111111111;
assign micromatrizz[20][554] = 9'b111111111;
assign micromatrizz[20][555] = 9'b111111111;
assign micromatrizz[20][556] = 9'b111111111;
assign micromatrizz[20][557] = 9'b111111111;
assign micromatrizz[20][558] = 9'b111111111;
assign micromatrizz[20][559] = 9'b111111111;
assign micromatrizz[20][560] = 9'b111111111;
assign micromatrizz[20][561] = 9'b111111111;
assign micromatrizz[20][562] = 9'b111111111;
assign micromatrizz[20][563] = 9'b111111111;
assign micromatrizz[20][564] = 9'b111111111;
assign micromatrizz[20][565] = 9'b111111111;
assign micromatrizz[20][566] = 9'b111111111;
assign micromatrizz[20][567] = 9'b111111111;
assign micromatrizz[20][568] = 9'b111111111;
assign micromatrizz[20][569] = 9'b111111111;
assign micromatrizz[20][570] = 9'b111111111;
assign micromatrizz[20][571] = 9'b111111111;
assign micromatrizz[20][572] = 9'b111111111;
assign micromatrizz[20][573] = 9'b111111111;
assign micromatrizz[20][574] = 9'b111111111;
assign micromatrizz[20][575] = 9'b111111111;
assign micromatrizz[20][576] = 9'b111111111;
assign micromatrizz[20][577] = 9'b111111111;
assign micromatrizz[20][578] = 9'b111111111;
assign micromatrizz[20][579] = 9'b111111111;
assign micromatrizz[20][580] = 9'b111111111;
assign micromatrizz[20][581] = 9'b111111111;
assign micromatrizz[20][582] = 9'b111111111;
assign micromatrizz[20][583] = 9'b111111111;
assign micromatrizz[20][584] = 9'b111111111;
assign micromatrizz[20][585] = 9'b111111111;
assign micromatrizz[20][586] = 9'b111111111;
assign micromatrizz[20][587] = 9'b111111111;
assign micromatrizz[20][588] = 9'b111111111;
assign micromatrizz[20][589] = 9'b111111111;
assign micromatrizz[20][590] = 9'b111111111;
assign micromatrizz[20][591] = 9'b111111111;
assign micromatrizz[20][592] = 9'b111111111;
assign micromatrizz[20][593] = 9'b111111111;
assign micromatrizz[20][594] = 9'b111111111;
assign micromatrizz[20][595] = 9'b111111111;
assign micromatrizz[20][596] = 9'b111111111;
assign micromatrizz[20][597] = 9'b111111111;
assign micromatrizz[20][598] = 9'b111111111;
assign micromatrizz[20][599] = 9'b111111111;
assign micromatrizz[20][600] = 9'b111111111;
assign micromatrizz[20][601] = 9'b111111111;
assign micromatrizz[20][602] = 9'b111111111;
assign micromatrizz[20][603] = 9'b111111111;
assign micromatrizz[20][604] = 9'b111111111;
assign micromatrizz[20][605] = 9'b111111111;
assign micromatrizz[20][606] = 9'b111111111;
assign micromatrizz[20][607] = 9'b111111111;
assign micromatrizz[20][608] = 9'b111111111;
assign micromatrizz[20][609] = 9'b111111111;
assign micromatrizz[20][610] = 9'b111111111;
assign micromatrizz[20][611] = 9'b111111111;
assign micromatrizz[20][612] = 9'b111111111;
assign micromatrizz[20][613] = 9'b111111111;
assign micromatrizz[20][614] = 9'b111111111;
assign micromatrizz[20][615] = 9'b111111111;
assign micromatrizz[20][616] = 9'b111111111;
assign micromatrizz[20][617] = 9'b111111111;
assign micromatrizz[20][618] = 9'b111111111;
assign micromatrizz[20][619] = 9'b111111111;
assign micromatrizz[20][620] = 9'b111111111;
assign micromatrizz[20][621] = 9'b111111111;
assign micromatrizz[20][622] = 9'b111111111;
assign micromatrizz[20][623] = 9'b111111111;
assign micromatrizz[20][624] = 9'b111111111;
assign micromatrizz[20][625] = 9'b111111111;
assign micromatrizz[20][626] = 9'b111111111;
assign micromatrizz[20][627] = 9'b111111111;
assign micromatrizz[20][628] = 9'b111111111;
assign micromatrizz[20][629] = 9'b111111111;
assign micromatrizz[20][630] = 9'b111111111;
assign micromatrizz[20][631] = 9'b111111111;
assign micromatrizz[20][632] = 9'b111111111;
assign micromatrizz[20][633] = 9'b111111111;
assign micromatrizz[20][634] = 9'b111111111;
assign micromatrizz[20][635] = 9'b111111111;
assign micromatrizz[20][636] = 9'b111111111;
assign micromatrizz[20][637] = 9'b111111111;
assign micromatrizz[20][638] = 9'b111111111;
assign micromatrizz[20][639] = 9'b111111111;
assign micromatrizz[21][0] = 9'b111111111;
assign micromatrizz[21][1] = 9'b111111111;
assign micromatrizz[21][2] = 9'b111111111;
assign micromatrizz[21][3] = 9'b111111111;
assign micromatrizz[21][4] = 9'b111111111;
assign micromatrizz[21][5] = 9'b111111111;
assign micromatrizz[21][6] = 9'b111111111;
assign micromatrizz[21][7] = 9'b111111111;
assign micromatrizz[21][8] = 9'b111111111;
assign micromatrizz[21][9] = 9'b111111111;
assign micromatrizz[21][10] = 9'b111111111;
assign micromatrizz[21][11] = 9'b111111111;
assign micromatrizz[21][12] = 9'b111111111;
assign micromatrizz[21][13] = 9'b111111111;
assign micromatrizz[21][14] = 9'b111111111;
assign micromatrizz[21][15] = 9'b111111111;
assign micromatrizz[21][16] = 9'b111111111;
assign micromatrizz[21][17] = 9'b111111111;
assign micromatrizz[21][18] = 9'b111111111;
assign micromatrizz[21][19] = 9'b111111111;
assign micromatrizz[21][20] = 9'b111111111;
assign micromatrizz[21][21] = 9'b111111111;
assign micromatrizz[21][22] = 9'b111111111;
assign micromatrizz[21][23] = 9'b111111111;
assign micromatrizz[21][24] = 9'b111111111;
assign micromatrizz[21][25] = 9'b111111111;
assign micromatrizz[21][26] = 9'b111111111;
assign micromatrizz[21][27] = 9'b111111111;
assign micromatrizz[21][28] = 9'b111111111;
assign micromatrizz[21][29] = 9'b111111111;
assign micromatrizz[21][30] = 9'b111111111;
assign micromatrizz[21][31] = 9'b111111111;
assign micromatrizz[21][32] = 9'b111111111;
assign micromatrizz[21][33] = 9'b111111111;
assign micromatrizz[21][34] = 9'b111111111;
assign micromatrizz[21][35] = 9'b111111111;
assign micromatrizz[21][36] = 9'b111111111;
assign micromatrizz[21][37] = 9'b111111111;
assign micromatrizz[21][38] = 9'b111111111;
assign micromatrizz[21][39] = 9'b111111111;
assign micromatrizz[21][40] = 9'b111111111;
assign micromatrizz[21][41] = 9'b111111111;
assign micromatrizz[21][42] = 9'b111111111;
assign micromatrizz[21][43] = 9'b111111111;
assign micromatrizz[21][44] = 9'b111111111;
assign micromatrizz[21][45] = 9'b111111111;
assign micromatrizz[21][46] = 9'b111111111;
assign micromatrizz[21][47] = 9'b111111111;
assign micromatrizz[21][48] = 9'b111111111;
assign micromatrizz[21][49] = 9'b111111111;
assign micromatrizz[21][50] = 9'b111111111;
assign micromatrizz[21][51] = 9'b111111111;
assign micromatrizz[21][52] = 9'b111111111;
assign micromatrizz[21][53] = 9'b111111111;
assign micromatrizz[21][54] = 9'b111111111;
assign micromatrizz[21][55] = 9'b111111111;
assign micromatrizz[21][56] = 9'b111111111;
assign micromatrizz[21][57] = 9'b111111111;
assign micromatrizz[21][58] = 9'b111111111;
assign micromatrizz[21][59] = 9'b111111111;
assign micromatrizz[21][60] = 9'b111111111;
assign micromatrizz[21][61] = 9'b111111111;
assign micromatrizz[21][62] = 9'b111111111;
assign micromatrizz[21][63] = 9'b111111111;
assign micromatrizz[21][64] = 9'b111111111;
assign micromatrizz[21][65] = 9'b111111111;
assign micromatrizz[21][66] = 9'b111111111;
assign micromatrizz[21][67] = 9'b111111111;
assign micromatrizz[21][68] = 9'b111111111;
assign micromatrizz[21][69] = 9'b111111111;
assign micromatrizz[21][70] = 9'b111111111;
assign micromatrizz[21][71] = 9'b111111111;
assign micromatrizz[21][72] = 9'b111111111;
assign micromatrizz[21][73] = 9'b111111111;
assign micromatrizz[21][74] = 9'b111111111;
assign micromatrizz[21][75] = 9'b111111111;
assign micromatrizz[21][76] = 9'b111111111;
assign micromatrizz[21][77] = 9'b111111111;
assign micromatrizz[21][78] = 9'b111111111;
assign micromatrizz[21][79] = 9'b111111111;
assign micromatrizz[21][80] = 9'b111111111;
assign micromatrizz[21][81] = 9'b111111111;
assign micromatrizz[21][82] = 9'b111111111;
assign micromatrizz[21][83] = 9'b111111111;
assign micromatrizz[21][84] = 9'b111111111;
assign micromatrizz[21][85] = 9'b111111111;
assign micromatrizz[21][86] = 9'b111111111;
assign micromatrizz[21][87] = 9'b111111111;
assign micromatrizz[21][88] = 9'b111111111;
assign micromatrizz[21][89] = 9'b111111111;
assign micromatrizz[21][90] = 9'b111111111;
assign micromatrizz[21][91] = 9'b111111111;
assign micromatrizz[21][92] = 9'b111111111;
assign micromatrizz[21][93] = 9'b111111111;
assign micromatrizz[21][94] = 9'b111111111;
assign micromatrizz[21][95] = 9'b111111111;
assign micromatrizz[21][96] = 9'b111111111;
assign micromatrizz[21][97] = 9'b111111111;
assign micromatrizz[21][98] = 9'b111111111;
assign micromatrizz[21][99] = 9'b111111111;
assign micromatrizz[21][100] = 9'b111111111;
assign micromatrizz[21][101] = 9'b111111111;
assign micromatrizz[21][102] = 9'b111111111;
assign micromatrizz[21][103] = 9'b111111111;
assign micromatrizz[21][104] = 9'b111111111;
assign micromatrizz[21][105] = 9'b111111111;
assign micromatrizz[21][106] = 9'b111111111;
assign micromatrizz[21][107] = 9'b111111111;
assign micromatrizz[21][108] = 9'b111111111;
assign micromatrizz[21][109] = 9'b111111111;
assign micromatrizz[21][110] = 9'b111111111;
assign micromatrizz[21][111] = 9'b111111111;
assign micromatrizz[21][112] = 9'b111111111;
assign micromatrizz[21][113] = 9'b111111111;
assign micromatrizz[21][114] = 9'b111111111;
assign micromatrizz[21][115] = 9'b111111111;
assign micromatrizz[21][116] = 9'b111111111;
assign micromatrizz[21][117] = 9'b111111111;
assign micromatrizz[21][118] = 9'b111111111;
assign micromatrizz[21][119] = 9'b111111111;
assign micromatrizz[21][120] = 9'b111111111;
assign micromatrizz[21][121] = 9'b111111111;
assign micromatrizz[21][122] = 9'b111111111;
assign micromatrizz[21][123] = 9'b111111111;
assign micromatrizz[21][124] = 9'b111111111;
assign micromatrizz[21][125] = 9'b111111111;
assign micromatrizz[21][126] = 9'b111111111;
assign micromatrizz[21][127] = 9'b111111111;
assign micromatrizz[21][128] = 9'b111111111;
assign micromatrizz[21][129] = 9'b111111111;
assign micromatrizz[21][130] = 9'b111111111;
assign micromatrizz[21][131] = 9'b111111111;
assign micromatrizz[21][132] = 9'b111111111;
assign micromatrizz[21][133] = 9'b111111111;
assign micromatrizz[21][134] = 9'b111111111;
assign micromatrizz[21][135] = 9'b111111111;
assign micromatrizz[21][136] = 9'b111111111;
assign micromatrizz[21][137] = 9'b111111111;
assign micromatrizz[21][138] = 9'b111111111;
assign micromatrizz[21][139] = 9'b111111111;
assign micromatrizz[21][140] = 9'b111111111;
assign micromatrizz[21][141] = 9'b111111111;
assign micromatrizz[21][142] = 9'b111111111;
assign micromatrizz[21][143] = 9'b111111111;
assign micromatrizz[21][144] = 9'b111111111;
assign micromatrizz[21][145] = 9'b111111111;
assign micromatrizz[21][146] = 9'b111111111;
assign micromatrizz[21][147] = 9'b111111111;
assign micromatrizz[21][148] = 9'b111111111;
assign micromatrizz[21][149] = 9'b111111111;
assign micromatrizz[21][150] = 9'b111111111;
assign micromatrizz[21][151] = 9'b111111111;
assign micromatrizz[21][152] = 9'b111111111;
assign micromatrizz[21][153] = 9'b111111111;
assign micromatrizz[21][154] = 9'b111111111;
assign micromatrizz[21][155] = 9'b111111111;
assign micromatrizz[21][156] = 9'b111111111;
assign micromatrizz[21][157] = 9'b111111111;
assign micromatrizz[21][158] = 9'b111111111;
assign micromatrizz[21][159] = 9'b111111111;
assign micromatrizz[21][160] = 9'b111111111;
assign micromatrizz[21][161] = 9'b111111111;
assign micromatrizz[21][162] = 9'b111111111;
assign micromatrizz[21][163] = 9'b111111111;
assign micromatrizz[21][164] = 9'b111111111;
assign micromatrizz[21][165] = 9'b111111111;
assign micromatrizz[21][166] = 9'b111111111;
assign micromatrizz[21][167] = 9'b111111111;
assign micromatrizz[21][168] = 9'b111111111;
assign micromatrizz[21][169] = 9'b111111111;
assign micromatrizz[21][170] = 9'b111111111;
assign micromatrizz[21][171] = 9'b111111111;
assign micromatrizz[21][172] = 9'b111111111;
assign micromatrizz[21][173] = 9'b111111111;
assign micromatrizz[21][174] = 9'b111111111;
assign micromatrizz[21][175] = 9'b111111111;
assign micromatrizz[21][176] = 9'b111111111;
assign micromatrizz[21][177] = 9'b111111111;
assign micromatrizz[21][178] = 9'b111111111;
assign micromatrizz[21][179] = 9'b111111111;
assign micromatrizz[21][180] = 9'b111111111;
assign micromatrizz[21][181] = 9'b111111111;
assign micromatrizz[21][182] = 9'b111111111;
assign micromatrizz[21][183] = 9'b111111111;
assign micromatrizz[21][184] = 9'b111111111;
assign micromatrizz[21][185] = 9'b111111111;
assign micromatrizz[21][186] = 9'b111111111;
assign micromatrizz[21][187] = 9'b111111111;
assign micromatrizz[21][188] = 9'b111111111;
assign micromatrizz[21][189] = 9'b111111111;
assign micromatrizz[21][190] = 9'b111111111;
assign micromatrizz[21][191] = 9'b111111111;
assign micromatrizz[21][192] = 9'b111111111;
assign micromatrizz[21][193] = 9'b111111111;
assign micromatrizz[21][194] = 9'b111111111;
assign micromatrizz[21][195] = 9'b111111111;
assign micromatrizz[21][196] = 9'b111111111;
assign micromatrizz[21][197] = 9'b111111111;
assign micromatrizz[21][198] = 9'b111111111;
assign micromatrizz[21][199] = 9'b111111111;
assign micromatrizz[21][200] = 9'b111111111;
assign micromatrizz[21][201] = 9'b111111111;
assign micromatrizz[21][202] = 9'b111111111;
assign micromatrizz[21][203] = 9'b111111111;
assign micromatrizz[21][204] = 9'b111111111;
assign micromatrizz[21][205] = 9'b111111111;
assign micromatrizz[21][206] = 9'b111111111;
assign micromatrizz[21][207] = 9'b111111111;
assign micromatrizz[21][208] = 9'b111111111;
assign micromatrizz[21][209] = 9'b111111111;
assign micromatrizz[21][210] = 9'b111111111;
assign micromatrizz[21][211] = 9'b111111111;
assign micromatrizz[21][212] = 9'b111111111;
assign micromatrizz[21][213] = 9'b111111111;
assign micromatrizz[21][214] = 9'b111111111;
assign micromatrizz[21][215] = 9'b111111111;
assign micromatrizz[21][216] = 9'b111111111;
assign micromatrizz[21][217] = 9'b111111111;
assign micromatrizz[21][218] = 9'b111111111;
assign micromatrizz[21][219] = 9'b111111111;
assign micromatrizz[21][220] = 9'b111111111;
assign micromatrizz[21][221] = 9'b111111111;
assign micromatrizz[21][222] = 9'b111111111;
assign micromatrizz[21][223] = 9'b111111111;
assign micromatrizz[21][224] = 9'b111111111;
assign micromatrizz[21][225] = 9'b111111111;
assign micromatrizz[21][226] = 9'b111111111;
assign micromatrizz[21][227] = 9'b111111111;
assign micromatrizz[21][228] = 9'b111111111;
assign micromatrizz[21][229] = 9'b111111111;
assign micromatrizz[21][230] = 9'b111111111;
assign micromatrizz[21][231] = 9'b111111111;
assign micromatrizz[21][232] = 9'b111111111;
assign micromatrizz[21][233] = 9'b111111111;
assign micromatrizz[21][234] = 9'b111111111;
assign micromatrizz[21][235] = 9'b111111111;
assign micromatrizz[21][236] = 9'b111111111;
assign micromatrizz[21][237] = 9'b111111111;
assign micromatrizz[21][238] = 9'b111111111;
assign micromatrizz[21][239] = 9'b111111111;
assign micromatrizz[21][240] = 9'b111111111;
assign micromatrizz[21][241] = 9'b111111111;
assign micromatrizz[21][242] = 9'b111111111;
assign micromatrizz[21][243] = 9'b111111111;
assign micromatrizz[21][244] = 9'b111111111;
assign micromatrizz[21][245] = 9'b111111111;
assign micromatrizz[21][246] = 9'b111111111;
assign micromatrizz[21][247] = 9'b111111111;
assign micromatrizz[21][248] = 9'b111111111;
assign micromatrizz[21][249] = 9'b111111111;
assign micromatrizz[21][250] = 9'b111111111;
assign micromatrizz[21][251] = 9'b111111111;
assign micromatrizz[21][252] = 9'b111111111;
assign micromatrizz[21][253] = 9'b111111111;
assign micromatrizz[21][254] = 9'b111111111;
assign micromatrizz[21][255] = 9'b111111111;
assign micromatrizz[21][256] = 9'b111111111;
assign micromatrizz[21][257] = 9'b111111111;
assign micromatrizz[21][258] = 9'b111111111;
assign micromatrizz[21][259] = 9'b111111111;
assign micromatrizz[21][260] = 9'b111111111;
assign micromatrizz[21][261] = 9'b111111111;
assign micromatrizz[21][262] = 9'b111111111;
assign micromatrizz[21][263] = 9'b111111111;
assign micromatrizz[21][264] = 9'b111111111;
assign micromatrizz[21][265] = 9'b111111111;
assign micromatrizz[21][266] = 9'b111111111;
assign micromatrizz[21][267] = 9'b111111111;
assign micromatrizz[21][268] = 9'b111111111;
assign micromatrizz[21][269] = 9'b111111111;
assign micromatrizz[21][270] = 9'b111110010;
assign micromatrizz[21][271] = 9'b111110010;
assign micromatrizz[21][272] = 9'b111110010;
assign micromatrizz[21][273] = 9'b111110010;
assign micromatrizz[21][274] = 9'b111110010;
assign micromatrizz[21][275] = 9'b111110011;
assign micromatrizz[21][276] = 9'b111110011;
assign micromatrizz[21][277] = 9'b111110011;
assign micromatrizz[21][278] = 9'b111110011;
assign micromatrizz[21][279] = 9'b111111111;
assign micromatrizz[21][280] = 9'b111111111;
assign micromatrizz[21][281] = 9'b111111111;
assign micromatrizz[21][282] = 9'b111111111;
assign micromatrizz[21][283] = 9'b111111111;
assign micromatrizz[21][284] = 9'b111111111;
assign micromatrizz[21][285] = 9'b111111111;
assign micromatrizz[21][286] = 9'b111111111;
assign micromatrizz[21][287] = 9'b111111111;
assign micromatrizz[21][288] = 9'b111111111;
assign micromatrizz[21][289] = 9'b111111111;
assign micromatrizz[21][290] = 9'b111111111;
assign micromatrizz[21][291] = 9'b111111111;
assign micromatrizz[21][292] = 9'b111111111;
assign micromatrizz[21][293] = 9'b111111111;
assign micromatrizz[21][294] = 9'b111111111;
assign micromatrizz[21][295] = 9'b111111111;
assign micromatrizz[21][296] = 9'b111111111;
assign micromatrizz[21][297] = 9'b111111111;
assign micromatrizz[21][298] = 9'b111111111;
assign micromatrizz[21][299] = 9'b111111111;
assign micromatrizz[21][300] = 9'b111111111;
assign micromatrizz[21][301] = 9'b111111111;
assign micromatrizz[21][302] = 9'b111111111;
assign micromatrizz[21][303] = 9'b111111111;
assign micromatrizz[21][304] = 9'b111111111;
assign micromatrizz[21][305] = 9'b111111111;
assign micromatrizz[21][306] = 9'b111111111;
assign micromatrizz[21][307] = 9'b111111111;
assign micromatrizz[21][308] = 9'b111111111;
assign micromatrizz[21][309] = 9'b111111111;
assign micromatrizz[21][310] = 9'b111111111;
assign micromatrizz[21][311] = 9'b111111111;
assign micromatrizz[21][312] = 9'b111111111;
assign micromatrizz[21][313] = 9'b111111111;
assign micromatrizz[21][314] = 9'b111111111;
assign micromatrizz[21][315] = 9'b111111111;
assign micromatrizz[21][316] = 9'b111111111;
assign micromatrizz[21][317] = 9'b111111111;
assign micromatrizz[21][318] = 9'b111111111;
assign micromatrizz[21][319] = 9'b111111111;
assign micromatrizz[21][320] = 9'b111111111;
assign micromatrizz[21][321] = 9'b111111111;
assign micromatrizz[21][322] = 9'b111111111;
assign micromatrizz[21][323] = 9'b111111111;
assign micromatrizz[21][324] = 9'b111111111;
assign micromatrizz[21][325] = 9'b111111111;
assign micromatrizz[21][326] = 9'b111111111;
assign micromatrizz[21][327] = 9'b111111111;
assign micromatrizz[21][328] = 9'b111111111;
assign micromatrizz[21][329] = 9'b111111111;
assign micromatrizz[21][330] = 9'b111111111;
assign micromatrizz[21][331] = 9'b111111111;
assign micromatrizz[21][332] = 9'b111111111;
assign micromatrizz[21][333] = 9'b111111111;
assign micromatrizz[21][334] = 9'b111111111;
assign micromatrizz[21][335] = 9'b111111111;
assign micromatrizz[21][336] = 9'b111111111;
assign micromatrizz[21][337] = 9'b111111111;
assign micromatrizz[21][338] = 9'b111111111;
assign micromatrizz[21][339] = 9'b111111111;
assign micromatrizz[21][340] = 9'b111111111;
assign micromatrizz[21][341] = 9'b111111111;
assign micromatrizz[21][342] = 9'b111111111;
assign micromatrizz[21][343] = 9'b111111111;
assign micromatrizz[21][344] = 9'b111111111;
assign micromatrizz[21][345] = 9'b111111111;
assign micromatrizz[21][346] = 9'b111111111;
assign micromatrizz[21][347] = 9'b111111111;
assign micromatrizz[21][348] = 9'b111111111;
assign micromatrizz[21][349] = 9'b111111111;
assign micromatrizz[21][350] = 9'b111111111;
assign micromatrizz[21][351] = 9'b111111111;
assign micromatrizz[21][352] = 9'b111111111;
assign micromatrizz[21][353] = 9'b111111111;
assign micromatrizz[21][354] = 9'b111111111;
assign micromatrizz[21][355] = 9'b111111111;
assign micromatrizz[21][356] = 9'b111111111;
assign micromatrizz[21][357] = 9'b111111111;
assign micromatrizz[21][358] = 9'b111111111;
assign micromatrizz[21][359] = 9'b111111111;
assign micromatrizz[21][360] = 9'b111111111;
assign micromatrizz[21][361] = 9'b111111111;
assign micromatrizz[21][362] = 9'b111111111;
assign micromatrizz[21][363] = 9'b111111111;
assign micromatrizz[21][364] = 9'b111111111;
assign micromatrizz[21][365] = 9'b111111111;
assign micromatrizz[21][366] = 9'b111111111;
assign micromatrizz[21][367] = 9'b111111111;
assign micromatrizz[21][368] = 9'b111111111;
assign micromatrizz[21][369] = 9'b111111111;
assign micromatrizz[21][370] = 9'b111111111;
assign micromatrizz[21][371] = 9'b111111111;
assign micromatrizz[21][372] = 9'b111111111;
assign micromatrizz[21][373] = 9'b111111111;
assign micromatrizz[21][374] = 9'b111111111;
assign micromatrizz[21][375] = 9'b111111111;
assign micromatrizz[21][376] = 9'b111111111;
assign micromatrizz[21][377] = 9'b111111111;
assign micromatrizz[21][378] = 9'b111111111;
assign micromatrizz[21][379] = 9'b111111111;
assign micromatrizz[21][380] = 9'b111111111;
assign micromatrizz[21][381] = 9'b111111111;
assign micromatrizz[21][382] = 9'b111111111;
assign micromatrizz[21][383] = 9'b111111111;
assign micromatrizz[21][384] = 9'b111111111;
assign micromatrizz[21][385] = 9'b111111111;
assign micromatrizz[21][386] = 9'b111111111;
assign micromatrizz[21][387] = 9'b111111111;
assign micromatrizz[21][388] = 9'b111111111;
assign micromatrizz[21][389] = 9'b111111111;
assign micromatrizz[21][390] = 9'b111111111;
assign micromatrizz[21][391] = 9'b111111111;
assign micromatrizz[21][392] = 9'b111111111;
assign micromatrizz[21][393] = 9'b111111111;
assign micromatrizz[21][394] = 9'b111111111;
assign micromatrizz[21][395] = 9'b111111111;
assign micromatrizz[21][396] = 9'b111111111;
assign micromatrizz[21][397] = 9'b111111111;
assign micromatrizz[21][398] = 9'b111111111;
assign micromatrizz[21][399] = 9'b111111111;
assign micromatrizz[21][400] = 9'b111111111;
assign micromatrizz[21][401] = 9'b111111111;
assign micromatrizz[21][402] = 9'b111111111;
assign micromatrizz[21][403] = 9'b111111111;
assign micromatrizz[21][404] = 9'b111111111;
assign micromatrizz[21][405] = 9'b111111111;
assign micromatrizz[21][406] = 9'b111111111;
assign micromatrizz[21][407] = 9'b111111111;
assign micromatrizz[21][408] = 9'b111111111;
assign micromatrizz[21][409] = 9'b111111111;
assign micromatrizz[21][410] = 9'b111111111;
assign micromatrizz[21][411] = 9'b111111111;
assign micromatrizz[21][412] = 9'b111111111;
assign micromatrizz[21][413] = 9'b111111111;
assign micromatrizz[21][414] = 9'b111111111;
assign micromatrizz[21][415] = 9'b111111111;
assign micromatrizz[21][416] = 9'b111111111;
assign micromatrizz[21][417] = 9'b111111111;
assign micromatrizz[21][418] = 9'b111111111;
assign micromatrizz[21][419] = 9'b111111111;
assign micromatrizz[21][420] = 9'b111111111;
assign micromatrizz[21][421] = 9'b111111111;
assign micromatrizz[21][422] = 9'b111111111;
assign micromatrizz[21][423] = 9'b111111111;
assign micromatrizz[21][424] = 9'b111111111;
assign micromatrizz[21][425] = 9'b111111111;
assign micromatrizz[21][426] = 9'b111111111;
assign micromatrizz[21][427] = 9'b111111111;
assign micromatrizz[21][428] = 9'b111111111;
assign micromatrizz[21][429] = 9'b111111111;
assign micromatrizz[21][430] = 9'b111111111;
assign micromatrizz[21][431] = 9'b111111111;
assign micromatrizz[21][432] = 9'b111111111;
assign micromatrizz[21][433] = 9'b111111111;
assign micromatrizz[21][434] = 9'b111111111;
assign micromatrizz[21][435] = 9'b111111111;
assign micromatrizz[21][436] = 9'b111111111;
assign micromatrizz[21][437] = 9'b111111111;
assign micromatrizz[21][438] = 9'b111111111;
assign micromatrizz[21][439] = 9'b111111111;
assign micromatrizz[21][440] = 9'b111111111;
assign micromatrizz[21][441] = 9'b111111111;
assign micromatrizz[21][442] = 9'b111111111;
assign micromatrizz[21][443] = 9'b111111111;
assign micromatrizz[21][444] = 9'b111111111;
assign micromatrizz[21][445] = 9'b111111111;
assign micromatrizz[21][446] = 9'b111111111;
assign micromatrizz[21][447] = 9'b111111111;
assign micromatrizz[21][448] = 9'b111111111;
assign micromatrizz[21][449] = 9'b111111111;
assign micromatrizz[21][450] = 9'b111111111;
assign micromatrizz[21][451] = 9'b111111111;
assign micromatrizz[21][452] = 9'b111111111;
assign micromatrizz[21][453] = 9'b111111111;
assign micromatrizz[21][454] = 9'b111111111;
assign micromatrizz[21][455] = 9'b111111111;
assign micromatrizz[21][456] = 9'b111111111;
assign micromatrizz[21][457] = 9'b111111111;
assign micromatrizz[21][458] = 9'b111111111;
assign micromatrizz[21][459] = 9'b111111111;
assign micromatrizz[21][460] = 9'b111111111;
assign micromatrizz[21][461] = 9'b111111111;
assign micromatrizz[21][462] = 9'b111111111;
assign micromatrizz[21][463] = 9'b111111111;
assign micromatrizz[21][464] = 9'b111111111;
assign micromatrizz[21][465] = 9'b111111111;
assign micromatrizz[21][466] = 9'b111111111;
assign micromatrizz[21][467] = 9'b111111111;
assign micromatrizz[21][468] = 9'b111111111;
assign micromatrizz[21][469] = 9'b111111111;
assign micromatrizz[21][470] = 9'b111111111;
assign micromatrizz[21][471] = 9'b111111111;
assign micromatrizz[21][472] = 9'b111111111;
assign micromatrizz[21][473] = 9'b111111111;
assign micromatrizz[21][474] = 9'b111111111;
assign micromatrizz[21][475] = 9'b111111111;
assign micromatrizz[21][476] = 9'b111111111;
assign micromatrizz[21][477] = 9'b111111111;
assign micromatrizz[21][478] = 9'b111111111;
assign micromatrizz[21][479] = 9'b111111111;
assign micromatrizz[21][480] = 9'b111111111;
assign micromatrizz[21][481] = 9'b111111111;
assign micromatrizz[21][482] = 9'b111111111;
assign micromatrizz[21][483] = 9'b111111111;
assign micromatrizz[21][484] = 9'b111111111;
assign micromatrizz[21][485] = 9'b111111111;
assign micromatrizz[21][486] = 9'b111111111;
assign micromatrizz[21][487] = 9'b111111111;
assign micromatrizz[21][488] = 9'b111111111;
assign micromatrizz[21][489] = 9'b111111111;
assign micromatrizz[21][490] = 9'b111111111;
assign micromatrizz[21][491] = 9'b111111111;
assign micromatrizz[21][492] = 9'b111111111;
assign micromatrizz[21][493] = 9'b111111111;
assign micromatrizz[21][494] = 9'b111111111;
assign micromatrizz[21][495] = 9'b111111111;
assign micromatrizz[21][496] = 9'b111111111;
assign micromatrizz[21][497] = 9'b111111111;
assign micromatrizz[21][498] = 9'b111111111;
assign micromatrizz[21][499] = 9'b111111111;
assign micromatrizz[21][500] = 9'b111111111;
assign micromatrizz[21][501] = 9'b111111111;
assign micromatrizz[21][502] = 9'b111111111;
assign micromatrizz[21][503] = 9'b111111111;
assign micromatrizz[21][504] = 9'b111111111;
assign micromatrizz[21][505] = 9'b111111111;
assign micromatrizz[21][506] = 9'b111111111;
assign micromatrizz[21][507] = 9'b111111111;
assign micromatrizz[21][508] = 9'b111111111;
assign micromatrizz[21][509] = 9'b111111111;
assign micromatrizz[21][510] = 9'b111111111;
assign micromatrizz[21][511] = 9'b111111111;
assign micromatrizz[21][512] = 9'b111111111;
assign micromatrizz[21][513] = 9'b111111111;
assign micromatrizz[21][514] = 9'b111111111;
assign micromatrizz[21][515] = 9'b111111111;
assign micromatrizz[21][516] = 9'b111111111;
assign micromatrizz[21][517] = 9'b111111111;
assign micromatrizz[21][518] = 9'b111111111;
assign micromatrizz[21][519] = 9'b111111111;
assign micromatrizz[21][520] = 9'b111111111;
assign micromatrizz[21][521] = 9'b111111111;
assign micromatrizz[21][522] = 9'b111111111;
assign micromatrizz[21][523] = 9'b111111111;
assign micromatrizz[21][524] = 9'b111111111;
assign micromatrizz[21][525] = 9'b111111111;
assign micromatrizz[21][526] = 9'b111111111;
assign micromatrizz[21][527] = 9'b111111111;
assign micromatrizz[21][528] = 9'b111111111;
assign micromatrizz[21][529] = 9'b111111111;
assign micromatrizz[21][530] = 9'b111111111;
assign micromatrizz[21][531] = 9'b111111111;
assign micromatrizz[21][532] = 9'b111111111;
assign micromatrizz[21][533] = 9'b111111111;
assign micromatrizz[21][534] = 9'b111111111;
assign micromatrizz[21][535] = 9'b111111111;
assign micromatrizz[21][536] = 9'b111111111;
assign micromatrizz[21][537] = 9'b111111111;
assign micromatrizz[21][538] = 9'b111111111;
assign micromatrizz[21][539] = 9'b111111111;
assign micromatrizz[21][540] = 9'b111111111;
assign micromatrizz[21][541] = 9'b111111111;
assign micromatrizz[21][542] = 9'b111111111;
assign micromatrizz[21][543] = 9'b111111111;
assign micromatrizz[21][544] = 9'b111111111;
assign micromatrizz[21][545] = 9'b111111111;
assign micromatrizz[21][546] = 9'b111111111;
assign micromatrizz[21][547] = 9'b111111111;
assign micromatrizz[21][548] = 9'b111111111;
assign micromatrizz[21][549] = 9'b111111111;
assign micromatrizz[21][550] = 9'b111111111;
assign micromatrizz[21][551] = 9'b111111111;
assign micromatrizz[21][552] = 9'b111111111;
assign micromatrizz[21][553] = 9'b111111111;
assign micromatrizz[21][554] = 9'b111111111;
assign micromatrizz[21][555] = 9'b111111111;
assign micromatrizz[21][556] = 9'b111111111;
assign micromatrizz[21][557] = 9'b111111111;
assign micromatrizz[21][558] = 9'b111111111;
assign micromatrizz[21][559] = 9'b111111111;
assign micromatrizz[21][560] = 9'b111111111;
assign micromatrizz[21][561] = 9'b111111111;
assign micromatrizz[21][562] = 9'b111111111;
assign micromatrizz[21][563] = 9'b111111111;
assign micromatrizz[21][564] = 9'b111111111;
assign micromatrizz[21][565] = 9'b111111111;
assign micromatrizz[21][566] = 9'b111111111;
assign micromatrizz[21][567] = 9'b111111111;
assign micromatrizz[21][568] = 9'b111111111;
assign micromatrizz[21][569] = 9'b111111111;
assign micromatrizz[21][570] = 9'b111111111;
assign micromatrizz[21][571] = 9'b111111111;
assign micromatrizz[21][572] = 9'b111111111;
assign micromatrizz[21][573] = 9'b111111111;
assign micromatrizz[21][574] = 9'b111111111;
assign micromatrizz[21][575] = 9'b111111111;
assign micromatrizz[21][576] = 9'b111111111;
assign micromatrizz[21][577] = 9'b111111111;
assign micromatrizz[21][578] = 9'b111111111;
assign micromatrizz[21][579] = 9'b111111111;
assign micromatrizz[21][580] = 9'b111111111;
assign micromatrizz[21][581] = 9'b111111111;
assign micromatrizz[21][582] = 9'b111111111;
assign micromatrizz[21][583] = 9'b111111111;
assign micromatrizz[21][584] = 9'b111111111;
assign micromatrizz[21][585] = 9'b111111111;
assign micromatrizz[21][586] = 9'b111111111;
assign micromatrizz[21][587] = 9'b111111111;
assign micromatrizz[21][588] = 9'b111111111;
assign micromatrizz[21][589] = 9'b111111111;
assign micromatrizz[21][590] = 9'b111111111;
assign micromatrizz[21][591] = 9'b111111111;
assign micromatrizz[21][592] = 9'b111111111;
assign micromatrizz[21][593] = 9'b111111111;
assign micromatrizz[21][594] = 9'b111111111;
assign micromatrizz[21][595] = 9'b111111111;
assign micromatrizz[21][596] = 9'b111111111;
assign micromatrizz[21][597] = 9'b111111111;
assign micromatrizz[21][598] = 9'b111111111;
assign micromatrizz[21][599] = 9'b111111111;
assign micromatrizz[21][600] = 9'b111111111;
assign micromatrizz[21][601] = 9'b111111111;
assign micromatrizz[21][602] = 9'b111111111;
assign micromatrizz[21][603] = 9'b111111111;
assign micromatrizz[21][604] = 9'b111111111;
assign micromatrizz[21][605] = 9'b111111111;
assign micromatrizz[21][606] = 9'b111111111;
assign micromatrizz[21][607] = 9'b111111111;
assign micromatrizz[21][608] = 9'b111111111;
assign micromatrizz[21][609] = 9'b111111111;
assign micromatrizz[21][610] = 9'b111111111;
assign micromatrizz[21][611] = 9'b111111111;
assign micromatrizz[21][612] = 9'b111111111;
assign micromatrizz[21][613] = 9'b111111111;
assign micromatrizz[21][614] = 9'b111111111;
assign micromatrizz[21][615] = 9'b111111111;
assign micromatrizz[21][616] = 9'b111111111;
assign micromatrizz[21][617] = 9'b111111111;
assign micromatrizz[21][618] = 9'b111111111;
assign micromatrizz[21][619] = 9'b111111111;
assign micromatrizz[21][620] = 9'b111111111;
assign micromatrizz[21][621] = 9'b111111111;
assign micromatrizz[21][622] = 9'b111111111;
assign micromatrizz[21][623] = 9'b111111111;
assign micromatrizz[21][624] = 9'b111111111;
assign micromatrizz[21][625] = 9'b111111111;
assign micromatrizz[21][626] = 9'b111111111;
assign micromatrizz[21][627] = 9'b111111111;
assign micromatrizz[21][628] = 9'b111111111;
assign micromatrizz[21][629] = 9'b111111111;
assign micromatrizz[21][630] = 9'b111111111;
assign micromatrizz[21][631] = 9'b111111111;
assign micromatrizz[21][632] = 9'b111111111;
assign micromatrizz[21][633] = 9'b111111111;
assign micromatrizz[21][634] = 9'b111111111;
assign micromatrizz[21][635] = 9'b111111111;
assign micromatrizz[21][636] = 9'b111111111;
assign micromatrizz[21][637] = 9'b111111111;
assign micromatrizz[21][638] = 9'b111111111;
assign micromatrizz[21][639] = 9'b111111111;
assign micromatrizz[22][0] = 9'b111111111;
assign micromatrizz[22][1] = 9'b111111111;
assign micromatrizz[22][2] = 9'b111111111;
assign micromatrizz[22][3] = 9'b111111111;
assign micromatrizz[22][4] = 9'b111111111;
assign micromatrizz[22][5] = 9'b111111111;
assign micromatrizz[22][6] = 9'b111111111;
assign micromatrizz[22][7] = 9'b111111111;
assign micromatrizz[22][8] = 9'b111111111;
assign micromatrizz[22][9] = 9'b111111111;
assign micromatrizz[22][10] = 9'b111111111;
assign micromatrizz[22][11] = 9'b111111111;
assign micromatrizz[22][12] = 9'b111111111;
assign micromatrizz[22][13] = 9'b111111111;
assign micromatrizz[22][14] = 9'b111111111;
assign micromatrizz[22][15] = 9'b111111111;
assign micromatrizz[22][16] = 9'b111111111;
assign micromatrizz[22][17] = 9'b111111111;
assign micromatrizz[22][18] = 9'b111111111;
assign micromatrizz[22][19] = 9'b111111111;
assign micromatrizz[22][20] = 9'b111111111;
assign micromatrizz[22][21] = 9'b111111111;
assign micromatrizz[22][22] = 9'b111111111;
assign micromatrizz[22][23] = 9'b111111111;
assign micromatrizz[22][24] = 9'b111111111;
assign micromatrizz[22][25] = 9'b111111111;
assign micromatrizz[22][26] = 9'b111111111;
assign micromatrizz[22][27] = 9'b111111111;
assign micromatrizz[22][28] = 9'b111111111;
assign micromatrizz[22][29] = 9'b111111111;
assign micromatrizz[22][30] = 9'b111111111;
assign micromatrizz[22][31] = 9'b111111111;
assign micromatrizz[22][32] = 9'b111111111;
assign micromatrizz[22][33] = 9'b111111111;
assign micromatrizz[22][34] = 9'b111111111;
assign micromatrizz[22][35] = 9'b111111111;
assign micromatrizz[22][36] = 9'b111111111;
assign micromatrizz[22][37] = 9'b111111111;
assign micromatrizz[22][38] = 9'b111111111;
assign micromatrizz[22][39] = 9'b111111111;
assign micromatrizz[22][40] = 9'b111111111;
assign micromatrizz[22][41] = 9'b111111111;
assign micromatrizz[22][42] = 9'b111111111;
assign micromatrizz[22][43] = 9'b111111111;
assign micromatrizz[22][44] = 9'b111111111;
assign micromatrizz[22][45] = 9'b111111111;
assign micromatrizz[22][46] = 9'b111111111;
assign micromatrizz[22][47] = 9'b111111111;
assign micromatrizz[22][48] = 9'b111111111;
assign micromatrizz[22][49] = 9'b111111111;
assign micromatrizz[22][50] = 9'b111111111;
assign micromatrizz[22][51] = 9'b111111111;
assign micromatrizz[22][52] = 9'b111111111;
assign micromatrizz[22][53] = 9'b111111111;
assign micromatrizz[22][54] = 9'b111111111;
assign micromatrizz[22][55] = 9'b111111111;
assign micromatrizz[22][56] = 9'b111111111;
assign micromatrizz[22][57] = 9'b111111111;
assign micromatrizz[22][58] = 9'b111111111;
assign micromatrizz[22][59] = 9'b111111111;
assign micromatrizz[22][60] = 9'b111111111;
assign micromatrizz[22][61] = 9'b111111111;
assign micromatrizz[22][62] = 9'b111111111;
assign micromatrizz[22][63] = 9'b111111111;
assign micromatrizz[22][64] = 9'b111111111;
assign micromatrizz[22][65] = 9'b111111111;
assign micromatrizz[22][66] = 9'b111111111;
assign micromatrizz[22][67] = 9'b111111111;
assign micromatrizz[22][68] = 9'b111111111;
assign micromatrizz[22][69] = 9'b111111111;
assign micromatrizz[22][70] = 9'b111111111;
assign micromatrizz[22][71] = 9'b111111111;
assign micromatrizz[22][72] = 9'b111111111;
assign micromatrizz[22][73] = 9'b111111111;
assign micromatrizz[22][74] = 9'b111111111;
assign micromatrizz[22][75] = 9'b111111111;
assign micromatrizz[22][76] = 9'b111111111;
assign micromatrizz[22][77] = 9'b111111111;
assign micromatrizz[22][78] = 9'b111111111;
assign micromatrizz[22][79] = 9'b111111111;
assign micromatrizz[22][80] = 9'b111111111;
assign micromatrizz[22][81] = 9'b111111111;
assign micromatrizz[22][82] = 9'b111111111;
assign micromatrizz[22][83] = 9'b111111111;
assign micromatrizz[22][84] = 9'b111111111;
assign micromatrizz[22][85] = 9'b111111111;
assign micromatrizz[22][86] = 9'b111111111;
assign micromatrizz[22][87] = 9'b111111111;
assign micromatrizz[22][88] = 9'b111111111;
assign micromatrizz[22][89] = 9'b111111111;
assign micromatrizz[22][90] = 9'b111111111;
assign micromatrizz[22][91] = 9'b111111111;
assign micromatrizz[22][92] = 9'b111111111;
assign micromatrizz[22][93] = 9'b111111111;
assign micromatrizz[22][94] = 9'b111111111;
assign micromatrizz[22][95] = 9'b111111111;
assign micromatrizz[22][96] = 9'b111111111;
assign micromatrizz[22][97] = 9'b111111111;
assign micromatrizz[22][98] = 9'b111111111;
assign micromatrizz[22][99] = 9'b111111111;
assign micromatrizz[22][100] = 9'b111111111;
assign micromatrizz[22][101] = 9'b111111111;
assign micromatrizz[22][102] = 9'b111111111;
assign micromatrizz[22][103] = 9'b111111111;
assign micromatrizz[22][104] = 9'b111111111;
assign micromatrizz[22][105] = 9'b111111111;
assign micromatrizz[22][106] = 9'b111111111;
assign micromatrizz[22][107] = 9'b111111111;
assign micromatrizz[22][108] = 9'b111111111;
assign micromatrizz[22][109] = 9'b111111111;
assign micromatrizz[22][110] = 9'b111111111;
assign micromatrizz[22][111] = 9'b111111111;
assign micromatrizz[22][112] = 9'b111111111;
assign micromatrizz[22][113] = 9'b111111111;
assign micromatrizz[22][114] = 9'b111111111;
assign micromatrizz[22][115] = 9'b111111111;
assign micromatrizz[22][116] = 9'b111111111;
assign micromatrizz[22][117] = 9'b111111111;
assign micromatrizz[22][118] = 9'b111111111;
assign micromatrizz[22][119] = 9'b111111111;
assign micromatrizz[22][120] = 9'b111111111;
assign micromatrizz[22][121] = 9'b111111111;
assign micromatrizz[22][122] = 9'b111111111;
assign micromatrizz[22][123] = 9'b111111111;
assign micromatrizz[22][124] = 9'b111111111;
assign micromatrizz[22][125] = 9'b111111111;
assign micromatrizz[22][126] = 9'b111111111;
assign micromatrizz[22][127] = 9'b111111111;
assign micromatrizz[22][128] = 9'b111111111;
assign micromatrizz[22][129] = 9'b111111111;
assign micromatrizz[22][130] = 9'b111111111;
assign micromatrizz[22][131] = 9'b111111111;
assign micromatrizz[22][132] = 9'b111111111;
assign micromatrizz[22][133] = 9'b111111111;
assign micromatrizz[22][134] = 9'b111111111;
assign micromatrizz[22][135] = 9'b111111111;
assign micromatrizz[22][136] = 9'b111111111;
assign micromatrizz[22][137] = 9'b111111111;
assign micromatrizz[22][138] = 9'b111111111;
assign micromatrizz[22][139] = 9'b111111111;
assign micromatrizz[22][140] = 9'b111111111;
assign micromatrizz[22][141] = 9'b111111111;
assign micromatrizz[22][142] = 9'b111111111;
assign micromatrizz[22][143] = 9'b111111111;
assign micromatrizz[22][144] = 9'b111111111;
assign micromatrizz[22][145] = 9'b111111111;
assign micromatrizz[22][146] = 9'b111111111;
assign micromatrizz[22][147] = 9'b111111111;
assign micromatrizz[22][148] = 9'b111111111;
assign micromatrizz[22][149] = 9'b111111111;
assign micromatrizz[22][150] = 9'b111111111;
assign micromatrizz[22][151] = 9'b111111111;
assign micromatrizz[22][152] = 9'b111111111;
assign micromatrizz[22][153] = 9'b111111111;
assign micromatrizz[22][154] = 9'b111111111;
assign micromatrizz[22][155] = 9'b111111111;
assign micromatrizz[22][156] = 9'b111111111;
assign micromatrizz[22][157] = 9'b111111111;
assign micromatrizz[22][158] = 9'b111111111;
assign micromatrizz[22][159] = 9'b111111111;
assign micromatrizz[22][160] = 9'b111111111;
assign micromatrizz[22][161] = 9'b111111111;
assign micromatrizz[22][162] = 9'b111111111;
assign micromatrizz[22][163] = 9'b111111111;
assign micromatrizz[22][164] = 9'b111111111;
assign micromatrizz[22][165] = 9'b111111111;
assign micromatrizz[22][166] = 9'b111111111;
assign micromatrizz[22][167] = 9'b111111111;
assign micromatrizz[22][168] = 9'b111111111;
assign micromatrizz[22][169] = 9'b111111111;
assign micromatrizz[22][170] = 9'b111111111;
assign micromatrizz[22][171] = 9'b111111111;
assign micromatrizz[22][172] = 9'b111111111;
assign micromatrizz[22][173] = 9'b111111111;
assign micromatrizz[22][174] = 9'b111111111;
assign micromatrizz[22][175] = 9'b111111111;
assign micromatrizz[22][176] = 9'b111111111;
assign micromatrizz[22][177] = 9'b111111111;
assign micromatrizz[22][178] = 9'b111111111;
assign micromatrizz[22][179] = 9'b111111111;
assign micromatrizz[22][180] = 9'b111111111;
assign micromatrizz[22][181] = 9'b111111111;
assign micromatrizz[22][182] = 9'b111111111;
assign micromatrizz[22][183] = 9'b111111111;
assign micromatrizz[22][184] = 9'b111111111;
assign micromatrizz[22][185] = 9'b111111111;
assign micromatrizz[22][186] = 9'b111111111;
assign micromatrizz[22][187] = 9'b111111111;
assign micromatrizz[22][188] = 9'b111111111;
assign micromatrizz[22][189] = 9'b111111111;
assign micromatrizz[22][190] = 9'b111111111;
assign micromatrizz[22][191] = 9'b111111111;
assign micromatrizz[22][192] = 9'b111111111;
assign micromatrizz[22][193] = 9'b111111111;
assign micromatrizz[22][194] = 9'b111111111;
assign micromatrizz[22][195] = 9'b111111111;
assign micromatrizz[22][196] = 9'b111111111;
assign micromatrizz[22][197] = 9'b111111111;
assign micromatrizz[22][198] = 9'b111111111;
assign micromatrizz[22][199] = 9'b111111111;
assign micromatrizz[22][200] = 9'b111111111;
assign micromatrizz[22][201] = 9'b111111111;
assign micromatrizz[22][202] = 9'b111111111;
assign micromatrizz[22][203] = 9'b111111111;
assign micromatrizz[22][204] = 9'b111111111;
assign micromatrizz[22][205] = 9'b111111111;
assign micromatrizz[22][206] = 9'b111111111;
assign micromatrizz[22][207] = 9'b111111111;
assign micromatrizz[22][208] = 9'b111111111;
assign micromatrizz[22][209] = 9'b111111111;
assign micromatrizz[22][210] = 9'b111111111;
assign micromatrizz[22][211] = 9'b111111111;
assign micromatrizz[22][212] = 9'b111111111;
assign micromatrizz[22][213] = 9'b111111111;
assign micromatrizz[22][214] = 9'b111111111;
assign micromatrizz[22][215] = 9'b111111111;
assign micromatrizz[22][216] = 9'b111111111;
assign micromatrizz[22][217] = 9'b111111111;
assign micromatrizz[22][218] = 9'b111111111;
assign micromatrizz[22][219] = 9'b111111111;
assign micromatrizz[22][220] = 9'b111111111;
assign micromatrizz[22][221] = 9'b111111111;
assign micromatrizz[22][222] = 9'b111111111;
assign micromatrizz[22][223] = 9'b111111111;
assign micromatrizz[22][224] = 9'b111111111;
assign micromatrizz[22][225] = 9'b111111111;
assign micromatrizz[22][226] = 9'b111111111;
assign micromatrizz[22][227] = 9'b111111111;
assign micromatrizz[22][228] = 9'b111111111;
assign micromatrizz[22][229] = 9'b111111111;
assign micromatrizz[22][230] = 9'b111111111;
assign micromatrizz[22][231] = 9'b111111111;
assign micromatrizz[22][232] = 9'b111111111;
assign micromatrizz[22][233] = 9'b111111111;
assign micromatrizz[22][234] = 9'b111111111;
assign micromatrizz[22][235] = 9'b111111111;
assign micromatrizz[22][236] = 9'b111111111;
assign micromatrizz[22][237] = 9'b111111111;
assign micromatrizz[22][238] = 9'b111111111;
assign micromatrizz[22][239] = 9'b111111111;
assign micromatrizz[22][240] = 9'b111111111;
assign micromatrizz[22][241] = 9'b111111111;
assign micromatrizz[22][242] = 9'b111111111;
assign micromatrizz[22][243] = 9'b111111111;
assign micromatrizz[22][244] = 9'b111111111;
assign micromatrizz[22][245] = 9'b111111111;
assign micromatrizz[22][246] = 9'b111111111;
assign micromatrizz[22][247] = 9'b111111111;
assign micromatrizz[22][248] = 9'b111111111;
assign micromatrizz[22][249] = 9'b111111111;
assign micromatrizz[22][250] = 9'b111111111;
assign micromatrizz[22][251] = 9'b111111111;
assign micromatrizz[22][252] = 9'b111111111;
assign micromatrizz[22][253] = 9'b111111111;
assign micromatrizz[22][254] = 9'b111111111;
assign micromatrizz[22][255] = 9'b111111111;
assign micromatrizz[22][256] = 9'b111111111;
assign micromatrizz[22][257] = 9'b111111111;
assign micromatrizz[22][258] = 9'b111111111;
assign micromatrizz[22][259] = 9'b111111111;
assign micromatrizz[22][260] = 9'b111111111;
assign micromatrizz[22][261] = 9'b111111111;
assign micromatrizz[22][262] = 9'b111111111;
assign micromatrizz[22][263] = 9'b111111111;
assign micromatrizz[22][264] = 9'b111111111;
assign micromatrizz[22][265] = 9'b111111111;
assign micromatrizz[22][266] = 9'b111111111;
assign micromatrizz[22][267] = 9'b111111111;
assign micromatrizz[22][268] = 9'b111111111;
assign micromatrizz[22][269] = 9'b111111111;
assign micromatrizz[22][270] = 9'b111110010;
assign micromatrizz[22][271] = 9'b111110010;
assign micromatrizz[22][272] = 9'b111110010;
assign micromatrizz[22][273] = 9'b111110010;
assign micromatrizz[22][274] = 9'b111110010;
assign micromatrizz[22][275] = 9'b111110011;
assign micromatrizz[22][276] = 9'b111110011;
assign micromatrizz[22][277] = 9'b111110011;
assign micromatrizz[22][278] = 9'b111110011;
assign micromatrizz[22][279] = 9'b111111111;
assign micromatrizz[22][280] = 9'b111111111;
assign micromatrizz[22][281] = 9'b111111111;
assign micromatrizz[22][282] = 9'b111111111;
assign micromatrizz[22][283] = 9'b111111111;
assign micromatrizz[22][284] = 9'b111111111;
assign micromatrizz[22][285] = 9'b111111111;
assign micromatrizz[22][286] = 9'b111111111;
assign micromatrizz[22][287] = 9'b111111111;
assign micromatrizz[22][288] = 9'b111111111;
assign micromatrizz[22][289] = 9'b111111111;
assign micromatrizz[22][290] = 9'b111111111;
assign micromatrizz[22][291] = 9'b111111111;
assign micromatrizz[22][292] = 9'b111111111;
assign micromatrizz[22][293] = 9'b111111111;
assign micromatrizz[22][294] = 9'b111110111;
assign micromatrizz[22][295] = 9'b111110111;
assign micromatrizz[22][296] = 9'b111110111;
assign micromatrizz[22][297] = 9'b111111111;
assign micromatrizz[22][298] = 9'b111111111;
assign micromatrizz[22][299] = 9'b111111111;
assign micromatrizz[22][300] = 9'b111111111;
assign micromatrizz[22][301] = 9'b111110111;
assign micromatrizz[22][302] = 9'b111111111;
assign micromatrizz[22][303] = 9'b111111111;
assign micromatrizz[22][304] = 9'b111111111;
assign micromatrizz[22][305] = 9'b111111111;
assign micromatrizz[22][306] = 9'b111111111;
assign micromatrizz[22][307] = 9'b111111111;
assign micromatrizz[22][308] = 9'b111111111;
assign micromatrizz[22][309] = 9'b111111111;
assign micromatrizz[22][310] = 9'b111111111;
assign micromatrizz[22][311] = 9'b111110111;
assign micromatrizz[22][312] = 9'b111110111;
assign micromatrizz[22][313] = 9'b111110111;
assign micromatrizz[22][314] = 9'b111111111;
assign micromatrizz[22][315] = 9'b111111111;
assign micromatrizz[22][316] = 9'b111111111;
assign micromatrizz[22][317] = 9'b111111111;
assign micromatrizz[22][318] = 9'b111111111;
assign micromatrizz[22][319] = 9'b111110111;
assign micromatrizz[22][320] = 9'b111111111;
assign micromatrizz[22][321] = 9'b111111111;
assign micromatrizz[22][322] = 9'b111111111;
assign micromatrizz[22][323] = 9'b111111111;
assign micromatrizz[22][324] = 9'b111111111;
assign micromatrizz[22][325] = 9'b111111111;
assign micromatrizz[22][326] = 9'b111111111;
assign micromatrizz[22][327] = 9'b111111111;
assign micromatrizz[22][328] = 9'b111111111;
assign micromatrizz[22][329] = 9'b111111111;
assign micromatrizz[22][330] = 9'b111111111;
assign micromatrizz[22][331] = 9'b111111111;
assign micromatrizz[22][332] = 9'b111111111;
assign micromatrizz[22][333] = 9'b111111111;
assign micromatrizz[22][334] = 9'b111111111;
assign micromatrizz[22][335] = 9'b111111111;
assign micromatrizz[22][336] = 9'b111111111;
assign micromatrizz[22][337] = 9'b111111111;
assign micromatrizz[22][338] = 9'b111111111;
assign micromatrizz[22][339] = 9'b111111111;
assign micromatrizz[22][340] = 9'b111111111;
assign micromatrizz[22][341] = 9'b111111111;
assign micromatrizz[22][342] = 9'b111111111;
assign micromatrizz[22][343] = 9'b111111111;
assign micromatrizz[22][344] = 9'b111111111;
assign micromatrizz[22][345] = 9'b111111111;
assign micromatrizz[22][346] = 9'b111111111;
assign micromatrizz[22][347] = 9'b111111111;
assign micromatrizz[22][348] = 9'b111111111;
assign micromatrizz[22][349] = 9'b111111111;
assign micromatrizz[22][350] = 9'b111111111;
assign micromatrizz[22][351] = 9'b111111111;
assign micromatrizz[22][352] = 9'b111111111;
assign micromatrizz[22][353] = 9'b111111111;
assign micromatrizz[22][354] = 9'b111111111;
assign micromatrizz[22][355] = 9'b111111111;
assign micromatrizz[22][356] = 9'b111111111;
assign micromatrizz[22][357] = 9'b111111111;
assign micromatrizz[22][358] = 9'b111111111;
assign micromatrizz[22][359] = 9'b111111111;
assign micromatrizz[22][360] = 9'b111111111;
assign micromatrizz[22][361] = 9'b111111111;
assign micromatrizz[22][362] = 9'b111111111;
assign micromatrizz[22][363] = 9'b111111111;
assign micromatrizz[22][364] = 9'b111111111;
assign micromatrizz[22][365] = 9'b111111111;
assign micromatrizz[22][366] = 9'b111111111;
assign micromatrizz[22][367] = 9'b111111111;
assign micromatrizz[22][368] = 9'b111111111;
assign micromatrizz[22][369] = 9'b111111111;
assign micromatrizz[22][370] = 9'b111111111;
assign micromatrizz[22][371] = 9'b111111111;
assign micromatrizz[22][372] = 9'b111111111;
assign micromatrizz[22][373] = 9'b111111111;
assign micromatrizz[22][374] = 9'b111111111;
assign micromatrizz[22][375] = 9'b111111111;
assign micromatrizz[22][376] = 9'b111111111;
assign micromatrizz[22][377] = 9'b111111111;
assign micromatrizz[22][378] = 9'b111111111;
assign micromatrizz[22][379] = 9'b111111111;
assign micromatrizz[22][380] = 9'b111111111;
assign micromatrizz[22][381] = 9'b111111111;
assign micromatrizz[22][382] = 9'b111111111;
assign micromatrizz[22][383] = 9'b111111111;
assign micromatrizz[22][384] = 9'b111111111;
assign micromatrizz[22][385] = 9'b111111111;
assign micromatrizz[22][386] = 9'b111111111;
assign micromatrizz[22][387] = 9'b111111111;
assign micromatrizz[22][388] = 9'b111111111;
assign micromatrizz[22][389] = 9'b111111111;
assign micromatrizz[22][390] = 9'b111111111;
assign micromatrizz[22][391] = 9'b111111111;
assign micromatrizz[22][392] = 9'b111111111;
assign micromatrizz[22][393] = 9'b111111111;
assign micromatrizz[22][394] = 9'b111111111;
assign micromatrizz[22][395] = 9'b111111111;
assign micromatrizz[22][396] = 9'b111111111;
assign micromatrizz[22][397] = 9'b111111111;
assign micromatrizz[22][398] = 9'b111111111;
assign micromatrizz[22][399] = 9'b111111111;
assign micromatrizz[22][400] = 9'b111111111;
assign micromatrizz[22][401] = 9'b111111111;
assign micromatrizz[22][402] = 9'b111111111;
assign micromatrizz[22][403] = 9'b111111111;
assign micromatrizz[22][404] = 9'b111111111;
assign micromatrizz[22][405] = 9'b111111111;
assign micromatrizz[22][406] = 9'b111111111;
assign micromatrizz[22][407] = 9'b111111111;
assign micromatrizz[22][408] = 9'b111111111;
assign micromatrizz[22][409] = 9'b111111111;
assign micromatrizz[22][410] = 9'b111111111;
assign micromatrizz[22][411] = 9'b111111111;
assign micromatrizz[22][412] = 9'b111111111;
assign micromatrizz[22][413] = 9'b111111111;
assign micromatrizz[22][414] = 9'b111111111;
assign micromatrizz[22][415] = 9'b111111111;
assign micromatrizz[22][416] = 9'b111111111;
assign micromatrizz[22][417] = 9'b111111111;
assign micromatrizz[22][418] = 9'b111111111;
assign micromatrizz[22][419] = 9'b111111111;
assign micromatrizz[22][420] = 9'b111111111;
assign micromatrizz[22][421] = 9'b111111111;
assign micromatrizz[22][422] = 9'b111111111;
assign micromatrizz[22][423] = 9'b111111111;
assign micromatrizz[22][424] = 9'b111111111;
assign micromatrizz[22][425] = 9'b111111111;
assign micromatrizz[22][426] = 9'b111111111;
assign micromatrizz[22][427] = 9'b111111111;
assign micromatrizz[22][428] = 9'b111111111;
assign micromatrizz[22][429] = 9'b111111111;
assign micromatrizz[22][430] = 9'b111111111;
assign micromatrizz[22][431] = 9'b111111111;
assign micromatrizz[22][432] = 9'b111111111;
assign micromatrizz[22][433] = 9'b111111111;
assign micromatrizz[22][434] = 9'b111111111;
assign micromatrizz[22][435] = 9'b111111111;
assign micromatrizz[22][436] = 9'b111111111;
assign micromatrizz[22][437] = 9'b111111111;
assign micromatrizz[22][438] = 9'b111111111;
assign micromatrizz[22][439] = 9'b111111111;
assign micromatrizz[22][440] = 9'b111111111;
assign micromatrizz[22][441] = 9'b111111111;
assign micromatrizz[22][442] = 9'b111111111;
assign micromatrizz[22][443] = 9'b111111111;
assign micromatrizz[22][444] = 9'b111111111;
assign micromatrizz[22][445] = 9'b111111111;
assign micromatrizz[22][446] = 9'b111111111;
assign micromatrizz[22][447] = 9'b111111111;
assign micromatrizz[22][448] = 9'b111111111;
assign micromatrizz[22][449] = 9'b111111111;
assign micromatrizz[22][450] = 9'b111111111;
assign micromatrizz[22][451] = 9'b111111111;
assign micromatrizz[22][452] = 9'b111111111;
assign micromatrizz[22][453] = 9'b111111111;
assign micromatrizz[22][454] = 9'b111111111;
assign micromatrizz[22][455] = 9'b111111111;
assign micromatrizz[22][456] = 9'b111111111;
assign micromatrizz[22][457] = 9'b111111111;
assign micromatrizz[22][458] = 9'b111111111;
assign micromatrizz[22][459] = 9'b111111111;
assign micromatrizz[22][460] = 9'b111111111;
assign micromatrizz[22][461] = 9'b111111111;
assign micromatrizz[22][462] = 9'b111111111;
assign micromatrizz[22][463] = 9'b111111111;
assign micromatrizz[22][464] = 9'b111111111;
assign micromatrizz[22][465] = 9'b111111111;
assign micromatrizz[22][466] = 9'b111111111;
assign micromatrizz[22][467] = 9'b111111111;
assign micromatrizz[22][468] = 9'b111111111;
assign micromatrizz[22][469] = 9'b111111111;
assign micromatrizz[22][470] = 9'b111111111;
assign micromatrizz[22][471] = 9'b111111111;
assign micromatrizz[22][472] = 9'b111111111;
assign micromatrizz[22][473] = 9'b111111111;
assign micromatrizz[22][474] = 9'b111111111;
assign micromatrizz[22][475] = 9'b111111111;
assign micromatrizz[22][476] = 9'b111111111;
assign micromatrizz[22][477] = 9'b111111111;
assign micromatrizz[22][478] = 9'b111111111;
assign micromatrizz[22][479] = 9'b111111111;
assign micromatrizz[22][480] = 9'b111111111;
assign micromatrizz[22][481] = 9'b111111111;
assign micromatrizz[22][482] = 9'b111111111;
assign micromatrizz[22][483] = 9'b111111111;
assign micromatrizz[22][484] = 9'b111111111;
assign micromatrizz[22][485] = 9'b111111111;
assign micromatrizz[22][486] = 9'b111111111;
assign micromatrizz[22][487] = 9'b111111111;
assign micromatrizz[22][488] = 9'b111111111;
assign micromatrizz[22][489] = 9'b111111111;
assign micromatrizz[22][490] = 9'b111111111;
assign micromatrizz[22][491] = 9'b111111111;
assign micromatrizz[22][492] = 9'b111111111;
assign micromatrizz[22][493] = 9'b111111111;
assign micromatrizz[22][494] = 9'b111111111;
assign micromatrizz[22][495] = 9'b111111111;
assign micromatrizz[22][496] = 9'b111111111;
assign micromatrizz[22][497] = 9'b111111111;
assign micromatrizz[22][498] = 9'b111111111;
assign micromatrizz[22][499] = 9'b111111111;
assign micromatrizz[22][500] = 9'b111111111;
assign micromatrizz[22][501] = 9'b111111111;
assign micromatrizz[22][502] = 9'b111111111;
assign micromatrizz[22][503] = 9'b111111111;
assign micromatrizz[22][504] = 9'b111111111;
assign micromatrizz[22][505] = 9'b111111111;
assign micromatrizz[22][506] = 9'b111111111;
assign micromatrizz[22][507] = 9'b111111111;
assign micromatrizz[22][508] = 9'b111111111;
assign micromatrizz[22][509] = 9'b111111111;
assign micromatrizz[22][510] = 9'b111111111;
assign micromatrizz[22][511] = 9'b111111111;
assign micromatrizz[22][512] = 9'b111111111;
assign micromatrizz[22][513] = 9'b111111111;
assign micromatrizz[22][514] = 9'b111111111;
assign micromatrizz[22][515] = 9'b111111111;
assign micromatrizz[22][516] = 9'b111111111;
assign micromatrizz[22][517] = 9'b111111111;
assign micromatrizz[22][518] = 9'b111111111;
assign micromatrizz[22][519] = 9'b111111111;
assign micromatrizz[22][520] = 9'b111111111;
assign micromatrizz[22][521] = 9'b111111111;
assign micromatrizz[22][522] = 9'b111111111;
assign micromatrizz[22][523] = 9'b111111111;
assign micromatrizz[22][524] = 9'b111111111;
assign micromatrizz[22][525] = 9'b111111111;
assign micromatrizz[22][526] = 9'b111111111;
assign micromatrizz[22][527] = 9'b111111111;
assign micromatrizz[22][528] = 9'b111111111;
assign micromatrizz[22][529] = 9'b111111111;
assign micromatrizz[22][530] = 9'b111111111;
assign micromatrizz[22][531] = 9'b111111111;
assign micromatrizz[22][532] = 9'b111111111;
assign micromatrizz[22][533] = 9'b111111111;
assign micromatrizz[22][534] = 9'b111111111;
assign micromatrizz[22][535] = 9'b111111111;
assign micromatrizz[22][536] = 9'b111111111;
assign micromatrizz[22][537] = 9'b111111111;
assign micromatrizz[22][538] = 9'b111111111;
assign micromatrizz[22][539] = 9'b111111111;
assign micromatrizz[22][540] = 9'b111111111;
assign micromatrizz[22][541] = 9'b111111111;
assign micromatrizz[22][542] = 9'b111111111;
assign micromatrizz[22][543] = 9'b111111111;
assign micromatrizz[22][544] = 9'b111111111;
assign micromatrizz[22][545] = 9'b111111111;
assign micromatrizz[22][546] = 9'b111111111;
assign micromatrizz[22][547] = 9'b111111111;
assign micromatrizz[22][548] = 9'b111111111;
assign micromatrizz[22][549] = 9'b111111111;
assign micromatrizz[22][550] = 9'b111111111;
assign micromatrizz[22][551] = 9'b111111111;
assign micromatrizz[22][552] = 9'b111111111;
assign micromatrizz[22][553] = 9'b111111111;
assign micromatrizz[22][554] = 9'b111111111;
assign micromatrizz[22][555] = 9'b111111111;
assign micromatrizz[22][556] = 9'b111111111;
assign micromatrizz[22][557] = 9'b111111111;
assign micromatrizz[22][558] = 9'b111111111;
assign micromatrizz[22][559] = 9'b111111111;
assign micromatrizz[22][560] = 9'b111111111;
assign micromatrizz[22][561] = 9'b111111111;
assign micromatrizz[22][562] = 9'b111111111;
assign micromatrizz[22][563] = 9'b111111111;
assign micromatrizz[22][564] = 9'b111111111;
assign micromatrizz[22][565] = 9'b111111111;
assign micromatrizz[22][566] = 9'b111111111;
assign micromatrizz[22][567] = 9'b111111111;
assign micromatrizz[22][568] = 9'b111111111;
assign micromatrizz[22][569] = 9'b111111111;
assign micromatrizz[22][570] = 9'b111111111;
assign micromatrizz[22][571] = 9'b111111111;
assign micromatrizz[22][572] = 9'b111111111;
assign micromatrizz[22][573] = 9'b111111111;
assign micromatrizz[22][574] = 9'b111111111;
assign micromatrizz[22][575] = 9'b111111111;
assign micromatrizz[22][576] = 9'b111111111;
assign micromatrizz[22][577] = 9'b111111111;
assign micromatrizz[22][578] = 9'b111111111;
assign micromatrizz[22][579] = 9'b111111111;
assign micromatrizz[22][580] = 9'b111111111;
assign micromatrizz[22][581] = 9'b111111111;
assign micromatrizz[22][582] = 9'b111111111;
assign micromatrizz[22][583] = 9'b111111111;
assign micromatrizz[22][584] = 9'b111111111;
assign micromatrizz[22][585] = 9'b111111111;
assign micromatrizz[22][586] = 9'b111111111;
assign micromatrizz[22][587] = 9'b111111111;
assign micromatrizz[22][588] = 9'b111111111;
assign micromatrizz[22][589] = 9'b111111111;
assign micromatrizz[22][590] = 9'b111111111;
assign micromatrizz[22][591] = 9'b111111111;
assign micromatrizz[22][592] = 9'b111111111;
assign micromatrizz[22][593] = 9'b111111111;
assign micromatrizz[22][594] = 9'b111111111;
assign micromatrizz[22][595] = 9'b111111111;
assign micromatrizz[22][596] = 9'b111111111;
assign micromatrizz[22][597] = 9'b111111111;
assign micromatrizz[22][598] = 9'b111111111;
assign micromatrizz[22][599] = 9'b111111111;
assign micromatrizz[22][600] = 9'b111111111;
assign micromatrizz[22][601] = 9'b111111111;
assign micromatrizz[22][602] = 9'b111111111;
assign micromatrizz[22][603] = 9'b111111111;
assign micromatrizz[22][604] = 9'b111111111;
assign micromatrizz[22][605] = 9'b111111111;
assign micromatrizz[22][606] = 9'b111111111;
assign micromatrizz[22][607] = 9'b111111111;
assign micromatrizz[22][608] = 9'b111111111;
assign micromatrizz[22][609] = 9'b111111111;
assign micromatrizz[22][610] = 9'b111111111;
assign micromatrizz[22][611] = 9'b111111111;
assign micromatrizz[22][612] = 9'b111111111;
assign micromatrizz[22][613] = 9'b111111111;
assign micromatrizz[22][614] = 9'b111111111;
assign micromatrizz[22][615] = 9'b111111111;
assign micromatrizz[22][616] = 9'b111111111;
assign micromatrizz[22][617] = 9'b111111111;
assign micromatrizz[22][618] = 9'b111111111;
assign micromatrizz[22][619] = 9'b111111111;
assign micromatrizz[22][620] = 9'b111111111;
assign micromatrizz[22][621] = 9'b111111111;
assign micromatrizz[22][622] = 9'b111111111;
assign micromatrizz[22][623] = 9'b111111111;
assign micromatrizz[22][624] = 9'b111111111;
assign micromatrizz[22][625] = 9'b111111111;
assign micromatrizz[22][626] = 9'b111111111;
assign micromatrizz[22][627] = 9'b111111111;
assign micromatrizz[22][628] = 9'b111111111;
assign micromatrizz[22][629] = 9'b111111111;
assign micromatrizz[22][630] = 9'b111111111;
assign micromatrizz[22][631] = 9'b111111111;
assign micromatrizz[22][632] = 9'b111111111;
assign micromatrizz[22][633] = 9'b111111111;
assign micromatrizz[22][634] = 9'b111111111;
assign micromatrizz[22][635] = 9'b111111111;
assign micromatrizz[22][636] = 9'b111111111;
assign micromatrizz[22][637] = 9'b111111111;
assign micromatrizz[22][638] = 9'b111111111;
assign micromatrizz[22][639] = 9'b111111111;
assign micromatrizz[23][0] = 9'b111111111;
assign micromatrizz[23][1] = 9'b111111111;
assign micromatrizz[23][2] = 9'b111111111;
assign micromatrizz[23][3] = 9'b111111111;
assign micromatrizz[23][4] = 9'b111111111;
assign micromatrizz[23][5] = 9'b111111111;
assign micromatrizz[23][6] = 9'b111111111;
assign micromatrizz[23][7] = 9'b111111111;
assign micromatrizz[23][8] = 9'b111111111;
assign micromatrizz[23][9] = 9'b111111111;
assign micromatrizz[23][10] = 9'b111111111;
assign micromatrizz[23][11] = 9'b111111111;
assign micromatrizz[23][12] = 9'b111111111;
assign micromatrizz[23][13] = 9'b111111111;
assign micromatrizz[23][14] = 9'b111111111;
assign micromatrizz[23][15] = 9'b111111111;
assign micromatrizz[23][16] = 9'b111111111;
assign micromatrizz[23][17] = 9'b111111111;
assign micromatrizz[23][18] = 9'b111111111;
assign micromatrizz[23][19] = 9'b111111111;
assign micromatrizz[23][20] = 9'b111111111;
assign micromatrizz[23][21] = 9'b111111111;
assign micromatrizz[23][22] = 9'b111111111;
assign micromatrizz[23][23] = 9'b111111111;
assign micromatrizz[23][24] = 9'b111111111;
assign micromatrizz[23][25] = 9'b111111111;
assign micromatrizz[23][26] = 9'b111111111;
assign micromatrizz[23][27] = 9'b111111111;
assign micromatrizz[23][28] = 9'b111111111;
assign micromatrizz[23][29] = 9'b111111111;
assign micromatrizz[23][30] = 9'b111111111;
assign micromatrizz[23][31] = 9'b111111111;
assign micromatrizz[23][32] = 9'b111111111;
assign micromatrizz[23][33] = 9'b111111111;
assign micromatrizz[23][34] = 9'b111111111;
assign micromatrizz[23][35] = 9'b111111111;
assign micromatrizz[23][36] = 9'b111111111;
assign micromatrizz[23][37] = 9'b111111111;
assign micromatrizz[23][38] = 9'b111111111;
assign micromatrizz[23][39] = 9'b111111111;
assign micromatrizz[23][40] = 9'b111111111;
assign micromatrizz[23][41] = 9'b111111111;
assign micromatrizz[23][42] = 9'b111111111;
assign micromatrizz[23][43] = 9'b111111111;
assign micromatrizz[23][44] = 9'b111111111;
assign micromatrizz[23][45] = 9'b111111111;
assign micromatrizz[23][46] = 9'b111111111;
assign micromatrizz[23][47] = 9'b111111111;
assign micromatrizz[23][48] = 9'b111111111;
assign micromatrizz[23][49] = 9'b111111111;
assign micromatrizz[23][50] = 9'b111111111;
assign micromatrizz[23][51] = 9'b111111111;
assign micromatrizz[23][52] = 9'b111111111;
assign micromatrizz[23][53] = 9'b111111111;
assign micromatrizz[23][54] = 9'b111111111;
assign micromatrizz[23][55] = 9'b111111111;
assign micromatrizz[23][56] = 9'b111111111;
assign micromatrizz[23][57] = 9'b111111111;
assign micromatrizz[23][58] = 9'b111111111;
assign micromatrizz[23][59] = 9'b111111111;
assign micromatrizz[23][60] = 9'b111111111;
assign micromatrizz[23][61] = 9'b111111111;
assign micromatrizz[23][62] = 9'b111111111;
assign micromatrizz[23][63] = 9'b111111111;
assign micromatrizz[23][64] = 9'b111111111;
assign micromatrizz[23][65] = 9'b111111111;
assign micromatrizz[23][66] = 9'b111111111;
assign micromatrizz[23][67] = 9'b111111111;
assign micromatrizz[23][68] = 9'b111111111;
assign micromatrizz[23][69] = 9'b111111111;
assign micromatrizz[23][70] = 9'b111111111;
assign micromatrizz[23][71] = 9'b111111111;
assign micromatrizz[23][72] = 9'b111111111;
assign micromatrizz[23][73] = 9'b111111111;
assign micromatrizz[23][74] = 9'b111111111;
assign micromatrizz[23][75] = 9'b111111111;
assign micromatrizz[23][76] = 9'b111111111;
assign micromatrizz[23][77] = 9'b111111111;
assign micromatrizz[23][78] = 9'b111111111;
assign micromatrizz[23][79] = 9'b111111111;
assign micromatrizz[23][80] = 9'b111111111;
assign micromatrizz[23][81] = 9'b111111111;
assign micromatrizz[23][82] = 9'b111111111;
assign micromatrizz[23][83] = 9'b111111111;
assign micromatrizz[23][84] = 9'b111111111;
assign micromatrizz[23][85] = 9'b111111111;
assign micromatrizz[23][86] = 9'b111111111;
assign micromatrizz[23][87] = 9'b111111111;
assign micromatrizz[23][88] = 9'b111111111;
assign micromatrizz[23][89] = 9'b111111111;
assign micromatrizz[23][90] = 9'b111111111;
assign micromatrizz[23][91] = 9'b111111111;
assign micromatrizz[23][92] = 9'b111111111;
assign micromatrizz[23][93] = 9'b111111111;
assign micromatrizz[23][94] = 9'b111111111;
assign micromatrizz[23][95] = 9'b111111111;
assign micromatrizz[23][96] = 9'b111111111;
assign micromatrizz[23][97] = 9'b111111111;
assign micromatrizz[23][98] = 9'b111111111;
assign micromatrizz[23][99] = 9'b111111111;
assign micromatrizz[23][100] = 9'b111111111;
assign micromatrizz[23][101] = 9'b111111111;
assign micromatrizz[23][102] = 9'b111111111;
assign micromatrizz[23][103] = 9'b111111111;
assign micromatrizz[23][104] = 9'b111111111;
assign micromatrizz[23][105] = 9'b111111111;
assign micromatrizz[23][106] = 9'b111111111;
assign micromatrizz[23][107] = 9'b111111111;
assign micromatrizz[23][108] = 9'b111111111;
assign micromatrizz[23][109] = 9'b111111111;
assign micromatrizz[23][110] = 9'b111111111;
assign micromatrizz[23][111] = 9'b111111111;
assign micromatrizz[23][112] = 9'b111111111;
assign micromatrizz[23][113] = 9'b111111111;
assign micromatrizz[23][114] = 9'b111111111;
assign micromatrizz[23][115] = 9'b111111111;
assign micromatrizz[23][116] = 9'b111111111;
assign micromatrizz[23][117] = 9'b111111111;
assign micromatrizz[23][118] = 9'b111111111;
assign micromatrizz[23][119] = 9'b111111111;
assign micromatrizz[23][120] = 9'b111111111;
assign micromatrizz[23][121] = 9'b111111111;
assign micromatrizz[23][122] = 9'b111111111;
assign micromatrizz[23][123] = 9'b111111111;
assign micromatrizz[23][124] = 9'b111111111;
assign micromatrizz[23][125] = 9'b111111111;
assign micromatrizz[23][126] = 9'b111111111;
assign micromatrizz[23][127] = 9'b111111111;
assign micromatrizz[23][128] = 9'b111111111;
assign micromatrizz[23][129] = 9'b111111111;
assign micromatrizz[23][130] = 9'b111111111;
assign micromatrizz[23][131] = 9'b111111111;
assign micromatrizz[23][132] = 9'b111111111;
assign micromatrizz[23][133] = 9'b111111111;
assign micromatrizz[23][134] = 9'b111111111;
assign micromatrizz[23][135] = 9'b111111111;
assign micromatrizz[23][136] = 9'b111111111;
assign micromatrizz[23][137] = 9'b111111111;
assign micromatrizz[23][138] = 9'b111111111;
assign micromatrizz[23][139] = 9'b111111111;
assign micromatrizz[23][140] = 9'b111111111;
assign micromatrizz[23][141] = 9'b111111111;
assign micromatrizz[23][142] = 9'b111111111;
assign micromatrizz[23][143] = 9'b111111111;
assign micromatrizz[23][144] = 9'b111111111;
assign micromatrizz[23][145] = 9'b111111111;
assign micromatrizz[23][146] = 9'b111111111;
assign micromatrizz[23][147] = 9'b111111111;
assign micromatrizz[23][148] = 9'b111111111;
assign micromatrizz[23][149] = 9'b111111111;
assign micromatrizz[23][150] = 9'b111111111;
assign micromatrizz[23][151] = 9'b111111111;
assign micromatrizz[23][152] = 9'b111111111;
assign micromatrizz[23][153] = 9'b111111111;
assign micromatrizz[23][154] = 9'b111111111;
assign micromatrizz[23][155] = 9'b111111111;
assign micromatrizz[23][156] = 9'b111111111;
assign micromatrizz[23][157] = 9'b111111111;
assign micromatrizz[23][158] = 9'b111111111;
assign micromatrizz[23][159] = 9'b111111111;
assign micromatrizz[23][160] = 9'b111111111;
assign micromatrizz[23][161] = 9'b111111111;
assign micromatrizz[23][162] = 9'b111111111;
assign micromatrizz[23][163] = 9'b111111111;
assign micromatrizz[23][164] = 9'b111111111;
assign micromatrizz[23][165] = 9'b111111111;
assign micromatrizz[23][166] = 9'b111111111;
assign micromatrizz[23][167] = 9'b111111111;
assign micromatrizz[23][168] = 9'b111111111;
assign micromatrizz[23][169] = 9'b111111111;
assign micromatrizz[23][170] = 9'b111111111;
assign micromatrizz[23][171] = 9'b111111111;
assign micromatrizz[23][172] = 9'b111111111;
assign micromatrizz[23][173] = 9'b111111111;
assign micromatrizz[23][174] = 9'b111111111;
assign micromatrizz[23][175] = 9'b111111111;
assign micromatrizz[23][176] = 9'b111111111;
assign micromatrizz[23][177] = 9'b111111111;
assign micromatrizz[23][178] = 9'b111111111;
assign micromatrizz[23][179] = 9'b111111111;
assign micromatrizz[23][180] = 9'b111111111;
assign micromatrizz[23][181] = 9'b111111111;
assign micromatrizz[23][182] = 9'b111111111;
assign micromatrizz[23][183] = 9'b111111111;
assign micromatrizz[23][184] = 9'b111111111;
assign micromatrizz[23][185] = 9'b111111111;
assign micromatrizz[23][186] = 9'b111111111;
assign micromatrizz[23][187] = 9'b111111111;
assign micromatrizz[23][188] = 9'b111111111;
assign micromatrizz[23][189] = 9'b111111111;
assign micromatrizz[23][190] = 9'b111111111;
assign micromatrizz[23][191] = 9'b111111111;
assign micromatrizz[23][192] = 9'b111111111;
assign micromatrizz[23][193] = 9'b111111111;
assign micromatrizz[23][194] = 9'b111111111;
assign micromatrizz[23][195] = 9'b111111111;
assign micromatrizz[23][196] = 9'b111111111;
assign micromatrizz[23][197] = 9'b111111111;
assign micromatrizz[23][198] = 9'b111111111;
assign micromatrizz[23][199] = 9'b111111111;
assign micromatrizz[23][200] = 9'b111111111;
assign micromatrizz[23][201] = 9'b111111111;
assign micromatrizz[23][202] = 9'b111111111;
assign micromatrizz[23][203] = 9'b111111111;
assign micromatrizz[23][204] = 9'b111111111;
assign micromatrizz[23][205] = 9'b111111111;
assign micromatrizz[23][206] = 9'b111111111;
assign micromatrizz[23][207] = 9'b111111111;
assign micromatrizz[23][208] = 9'b111111111;
assign micromatrizz[23][209] = 9'b111111111;
assign micromatrizz[23][210] = 9'b111111111;
assign micromatrizz[23][211] = 9'b111111111;
assign micromatrizz[23][212] = 9'b111111111;
assign micromatrizz[23][213] = 9'b111111111;
assign micromatrizz[23][214] = 9'b111111111;
assign micromatrizz[23][215] = 9'b111111111;
assign micromatrizz[23][216] = 9'b111111111;
assign micromatrizz[23][217] = 9'b111111111;
assign micromatrizz[23][218] = 9'b111111111;
assign micromatrizz[23][219] = 9'b111111111;
assign micromatrizz[23][220] = 9'b111111111;
assign micromatrizz[23][221] = 9'b111111111;
assign micromatrizz[23][222] = 9'b111111111;
assign micromatrizz[23][223] = 9'b111111111;
assign micromatrizz[23][224] = 9'b111111111;
assign micromatrizz[23][225] = 9'b111111111;
assign micromatrizz[23][226] = 9'b111111111;
assign micromatrizz[23][227] = 9'b111111111;
assign micromatrizz[23][228] = 9'b111111111;
assign micromatrizz[23][229] = 9'b111111111;
assign micromatrizz[23][230] = 9'b111111111;
assign micromatrizz[23][231] = 9'b111111111;
assign micromatrizz[23][232] = 9'b111111111;
assign micromatrizz[23][233] = 9'b111111111;
assign micromatrizz[23][234] = 9'b111111111;
assign micromatrizz[23][235] = 9'b111111111;
assign micromatrizz[23][236] = 9'b111111111;
assign micromatrizz[23][237] = 9'b111111111;
assign micromatrizz[23][238] = 9'b111111111;
assign micromatrizz[23][239] = 9'b111111111;
assign micromatrizz[23][240] = 9'b111111111;
assign micromatrizz[23][241] = 9'b111111111;
assign micromatrizz[23][242] = 9'b111111111;
assign micromatrizz[23][243] = 9'b111111111;
assign micromatrizz[23][244] = 9'b111111111;
assign micromatrizz[23][245] = 9'b111111111;
assign micromatrizz[23][246] = 9'b111111111;
assign micromatrizz[23][247] = 9'b111111111;
assign micromatrizz[23][248] = 9'b111111111;
assign micromatrizz[23][249] = 9'b111111111;
assign micromatrizz[23][250] = 9'b111111111;
assign micromatrizz[23][251] = 9'b111111111;
assign micromatrizz[23][252] = 9'b111111111;
assign micromatrizz[23][253] = 9'b111111111;
assign micromatrizz[23][254] = 9'b111111111;
assign micromatrizz[23][255] = 9'b111111111;
assign micromatrizz[23][256] = 9'b111111111;
assign micromatrizz[23][257] = 9'b111111111;
assign micromatrizz[23][258] = 9'b111111111;
assign micromatrizz[23][259] = 9'b111111111;
assign micromatrizz[23][260] = 9'b111111111;
assign micromatrizz[23][261] = 9'b111111111;
assign micromatrizz[23][262] = 9'b111111111;
assign micromatrizz[23][263] = 9'b111111111;
assign micromatrizz[23][264] = 9'b111111111;
assign micromatrizz[23][265] = 9'b111111111;
assign micromatrizz[23][266] = 9'b111111111;
assign micromatrizz[23][267] = 9'b111111111;
assign micromatrizz[23][268] = 9'b111111111;
assign micromatrizz[23][269] = 9'b111111111;
assign micromatrizz[23][270] = 9'b111110010;
assign micromatrizz[23][271] = 9'b111110010;
assign micromatrizz[23][272] = 9'b111110010;
assign micromatrizz[23][273] = 9'b111110010;
assign micromatrizz[23][274] = 9'b111110010;
assign micromatrizz[23][275] = 9'b111110011;
assign micromatrizz[23][276] = 9'b111110011;
assign micromatrizz[23][277] = 9'b111110011;
assign micromatrizz[23][278] = 9'b111110011;
assign micromatrizz[23][279] = 9'b111111111;
assign micromatrizz[23][280] = 9'b111111111;
assign micromatrizz[23][281] = 9'b111111111;
assign micromatrizz[23][282] = 9'b111111111;
assign micromatrizz[23][283] = 9'b111111111;
assign micromatrizz[23][284] = 9'b111111111;
assign micromatrizz[23][285] = 9'b111111111;
assign micromatrizz[23][286] = 9'b111111111;
assign micromatrizz[23][287] = 9'b111111111;
assign micromatrizz[23][288] = 9'b111111111;
assign micromatrizz[23][289] = 9'b111111111;
assign micromatrizz[23][290] = 9'b111111111;
assign micromatrizz[23][291] = 9'b111111111;
assign micromatrizz[23][292] = 9'b111111111;
assign micromatrizz[23][293] = 9'b111110111;
assign micromatrizz[23][294] = 9'b111110010;
assign micromatrizz[23][295] = 9'b111110011;
assign micromatrizz[23][296] = 9'b111110010;
assign micromatrizz[23][297] = 9'b111110111;
assign micromatrizz[23][298] = 9'b111111111;
assign micromatrizz[23][299] = 9'b111111111;
assign micromatrizz[23][300] = 9'b111111111;
assign micromatrizz[23][301] = 9'b111111111;
assign micromatrizz[23][302] = 9'b111110111;
assign micromatrizz[23][303] = 9'b111111111;
assign micromatrizz[23][304] = 9'b111111111;
assign micromatrizz[23][305] = 9'b111111111;
assign micromatrizz[23][306] = 9'b111111111;
assign micromatrizz[23][307] = 9'b111111111;
assign micromatrizz[23][308] = 9'b111111111;
assign micromatrizz[23][309] = 9'b111111111;
assign micromatrizz[23][310] = 9'b111110110;
assign micromatrizz[23][311] = 9'b111110010;
assign micromatrizz[23][312] = 9'b111110010;
assign micromatrizz[23][313] = 9'b111110010;
assign micromatrizz[23][314] = 9'b111111111;
assign micromatrizz[23][315] = 9'b111111111;
assign micromatrizz[23][316] = 9'b111111111;
assign micromatrizz[23][317] = 9'b111111111;
assign micromatrizz[23][318] = 9'b111111111;
assign micromatrizz[23][319] = 9'b111110111;
assign micromatrizz[23][320] = 9'b111110111;
assign micromatrizz[23][321] = 9'b111111111;
assign micromatrizz[23][322] = 9'b111111111;
assign micromatrizz[23][323] = 9'b111111111;
assign micromatrizz[23][324] = 9'b111111111;
assign micromatrizz[23][325] = 9'b111111111;
assign micromatrizz[23][326] = 9'b111111111;
assign micromatrizz[23][327] = 9'b111111111;
assign micromatrizz[23][328] = 9'b111111111;
assign micromatrizz[23][329] = 9'b111111111;
assign micromatrizz[23][330] = 9'b111111111;
assign micromatrizz[23][331] = 9'b111111111;
assign micromatrizz[23][332] = 9'b111111111;
assign micromatrizz[23][333] = 9'b111111111;
assign micromatrizz[23][334] = 9'b111111111;
assign micromatrizz[23][335] = 9'b111111111;
assign micromatrizz[23][336] = 9'b111111111;
assign micromatrizz[23][337] = 9'b111111111;
assign micromatrizz[23][338] = 9'b111111111;
assign micromatrizz[23][339] = 9'b111111111;
assign micromatrizz[23][340] = 9'b111111111;
assign micromatrizz[23][341] = 9'b111111111;
assign micromatrizz[23][342] = 9'b111111111;
assign micromatrizz[23][343] = 9'b111111111;
assign micromatrizz[23][344] = 9'b111111111;
assign micromatrizz[23][345] = 9'b111111111;
assign micromatrizz[23][346] = 9'b111111111;
assign micromatrizz[23][347] = 9'b111111111;
assign micromatrizz[23][348] = 9'b111111111;
assign micromatrizz[23][349] = 9'b111111111;
assign micromatrizz[23][350] = 9'b111111111;
assign micromatrizz[23][351] = 9'b111111111;
assign micromatrizz[23][352] = 9'b111111111;
assign micromatrizz[23][353] = 9'b111111111;
assign micromatrizz[23][354] = 9'b111111111;
assign micromatrizz[23][355] = 9'b111111111;
assign micromatrizz[23][356] = 9'b111111111;
assign micromatrizz[23][357] = 9'b111111111;
assign micromatrizz[23][358] = 9'b111111111;
assign micromatrizz[23][359] = 9'b111111111;
assign micromatrizz[23][360] = 9'b111111111;
assign micromatrizz[23][361] = 9'b111111111;
assign micromatrizz[23][362] = 9'b111111111;
assign micromatrizz[23][363] = 9'b111111111;
assign micromatrizz[23][364] = 9'b111111111;
assign micromatrizz[23][365] = 9'b111111111;
assign micromatrizz[23][366] = 9'b111111111;
assign micromatrizz[23][367] = 9'b111111111;
assign micromatrizz[23][368] = 9'b111111111;
assign micromatrizz[23][369] = 9'b111111111;
assign micromatrizz[23][370] = 9'b111111111;
assign micromatrizz[23][371] = 9'b111111111;
assign micromatrizz[23][372] = 9'b111111111;
assign micromatrizz[23][373] = 9'b111111111;
assign micromatrizz[23][374] = 9'b111111111;
assign micromatrizz[23][375] = 9'b111111111;
assign micromatrizz[23][376] = 9'b111111111;
assign micromatrizz[23][377] = 9'b111111111;
assign micromatrizz[23][378] = 9'b111111111;
assign micromatrizz[23][379] = 9'b111111111;
assign micromatrizz[23][380] = 9'b111111111;
assign micromatrizz[23][381] = 9'b111111111;
assign micromatrizz[23][382] = 9'b111111111;
assign micromatrizz[23][383] = 9'b111111111;
assign micromatrizz[23][384] = 9'b111111111;
assign micromatrizz[23][385] = 9'b111111111;
assign micromatrizz[23][386] = 9'b111111111;
assign micromatrizz[23][387] = 9'b111111111;
assign micromatrizz[23][388] = 9'b111111111;
assign micromatrizz[23][389] = 9'b111111111;
assign micromatrizz[23][390] = 9'b111111111;
assign micromatrizz[23][391] = 9'b111111111;
assign micromatrizz[23][392] = 9'b111111111;
assign micromatrizz[23][393] = 9'b111111111;
assign micromatrizz[23][394] = 9'b111111111;
assign micromatrizz[23][395] = 9'b111111111;
assign micromatrizz[23][396] = 9'b111111111;
assign micromatrizz[23][397] = 9'b111111111;
assign micromatrizz[23][398] = 9'b111111111;
assign micromatrizz[23][399] = 9'b111111111;
assign micromatrizz[23][400] = 9'b111111111;
assign micromatrizz[23][401] = 9'b111111111;
assign micromatrizz[23][402] = 9'b111111111;
assign micromatrizz[23][403] = 9'b111111111;
assign micromatrizz[23][404] = 9'b111111111;
assign micromatrizz[23][405] = 9'b111111111;
assign micromatrizz[23][406] = 9'b111111111;
assign micromatrizz[23][407] = 9'b111111111;
assign micromatrizz[23][408] = 9'b111111111;
assign micromatrizz[23][409] = 9'b111111111;
assign micromatrizz[23][410] = 9'b111111111;
assign micromatrizz[23][411] = 9'b111111111;
assign micromatrizz[23][412] = 9'b111111111;
assign micromatrizz[23][413] = 9'b111111111;
assign micromatrizz[23][414] = 9'b111111111;
assign micromatrizz[23][415] = 9'b111111111;
assign micromatrizz[23][416] = 9'b111111111;
assign micromatrizz[23][417] = 9'b111111111;
assign micromatrizz[23][418] = 9'b111111111;
assign micromatrizz[23][419] = 9'b111111111;
assign micromatrizz[23][420] = 9'b111111111;
assign micromatrizz[23][421] = 9'b111111111;
assign micromatrizz[23][422] = 9'b111111111;
assign micromatrizz[23][423] = 9'b111111111;
assign micromatrizz[23][424] = 9'b111111111;
assign micromatrizz[23][425] = 9'b111111111;
assign micromatrizz[23][426] = 9'b111111111;
assign micromatrizz[23][427] = 9'b111111111;
assign micromatrizz[23][428] = 9'b111111111;
assign micromatrizz[23][429] = 9'b111111111;
assign micromatrizz[23][430] = 9'b111111111;
assign micromatrizz[23][431] = 9'b111111111;
assign micromatrizz[23][432] = 9'b111111111;
assign micromatrizz[23][433] = 9'b111111111;
assign micromatrizz[23][434] = 9'b111111111;
assign micromatrizz[23][435] = 9'b111111111;
assign micromatrizz[23][436] = 9'b111111111;
assign micromatrizz[23][437] = 9'b111111111;
assign micromatrizz[23][438] = 9'b111111111;
assign micromatrizz[23][439] = 9'b111111111;
assign micromatrizz[23][440] = 9'b111111111;
assign micromatrizz[23][441] = 9'b111111111;
assign micromatrizz[23][442] = 9'b111111111;
assign micromatrizz[23][443] = 9'b111111111;
assign micromatrizz[23][444] = 9'b111111111;
assign micromatrizz[23][445] = 9'b111111111;
assign micromatrizz[23][446] = 9'b111111111;
assign micromatrizz[23][447] = 9'b111111111;
assign micromatrizz[23][448] = 9'b111111111;
assign micromatrizz[23][449] = 9'b111111111;
assign micromatrizz[23][450] = 9'b111111111;
assign micromatrizz[23][451] = 9'b111111111;
assign micromatrizz[23][452] = 9'b111111111;
assign micromatrizz[23][453] = 9'b111111111;
assign micromatrizz[23][454] = 9'b111111111;
assign micromatrizz[23][455] = 9'b111111111;
assign micromatrizz[23][456] = 9'b111111111;
assign micromatrizz[23][457] = 9'b111111111;
assign micromatrizz[23][458] = 9'b111111111;
assign micromatrizz[23][459] = 9'b111111111;
assign micromatrizz[23][460] = 9'b111111111;
assign micromatrizz[23][461] = 9'b111111111;
assign micromatrizz[23][462] = 9'b111111111;
assign micromatrizz[23][463] = 9'b111111111;
assign micromatrizz[23][464] = 9'b111111111;
assign micromatrizz[23][465] = 9'b111111111;
assign micromatrizz[23][466] = 9'b111111111;
assign micromatrizz[23][467] = 9'b111111111;
assign micromatrizz[23][468] = 9'b111111111;
assign micromatrizz[23][469] = 9'b111111111;
assign micromatrizz[23][470] = 9'b111111111;
assign micromatrizz[23][471] = 9'b111111111;
assign micromatrizz[23][472] = 9'b111111111;
assign micromatrizz[23][473] = 9'b111111111;
assign micromatrizz[23][474] = 9'b111111111;
assign micromatrizz[23][475] = 9'b111111111;
assign micromatrizz[23][476] = 9'b111111111;
assign micromatrizz[23][477] = 9'b111111111;
assign micromatrizz[23][478] = 9'b111111111;
assign micromatrizz[23][479] = 9'b111111111;
assign micromatrizz[23][480] = 9'b111111111;
assign micromatrizz[23][481] = 9'b111111111;
assign micromatrizz[23][482] = 9'b111111111;
assign micromatrizz[23][483] = 9'b111111111;
assign micromatrizz[23][484] = 9'b111111111;
assign micromatrizz[23][485] = 9'b111111111;
assign micromatrizz[23][486] = 9'b111111111;
assign micromatrizz[23][487] = 9'b111111111;
assign micromatrizz[23][488] = 9'b111111111;
assign micromatrizz[23][489] = 9'b111111111;
assign micromatrizz[23][490] = 9'b111111111;
assign micromatrizz[23][491] = 9'b111111111;
assign micromatrizz[23][492] = 9'b111111111;
assign micromatrizz[23][493] = 9'b111111111;
assign micromatrizz[23][494] = 9'b111111111;
assign micromatrizz[23][495] = 9'b111111111;
assign micromatrizz[23][496] = 9'b111111111;
assign micromatrizz[23][497] = 9'b111111111;
assign micromatrizz[23][498] = 9'b111111111;
assign micromatrizz[23][499] = 9'b111111111;
assign micromatrizz[23][500] = 9'b111111111;
assign micromatrizz[23][501] = 9'b111111111;
assign micromatrizz[23][502] = 9'b111111111;
assign micromatrizz[23][503] = 9'b111111111;
assign micromatrizz[23][504] = 9'b111111111;
assign micromatrizz[23][505] = 9'b111111111;
assign micromatrizz[23][506] = 9'b111111111;
assign micromatrizz[23][507] = 9'b111111111;
assign micromatrizz[23][508] = 9'b111111111;
assign micromatrizz[23][509] = 9'b111111111;
assign micromatrizz[23][510] = 9'b111111111;
assign micromatrizz[23][511] = 9'b111111111;
assign micromatrizz[23][512] = 9'b111111111;
assign micromatrizz[23][513] = 9'b111111111;
assign micromatrizz[23][514] = 9'b111111111;
assign micromatrizz[23][515] = 9'b111111111;
assign micromatrizz[23][516] = 9'b111111111;
assign micromatrizz[23][517] = 9'b111111111;
assign micromatrizz[23][518] = 9'b111111111;
assign micromatrizz[23][519] = 9'b111111111;
assign micromatrizz[23][520] = 9'b111111111;
assign micromatrizz[23][521] = 9'b111111111;
assign micromatrizz[23][522] = 9'b111111111;
assign micromatrizz[23][523] = 9'b111111111;
assign micromatrizz[23][524] = 9'b111111111;
assign micromatrizz[23][525] = 9'b111111111;
assign micromatrizz[23][526] = 9'b111111111;
assign micromatrizz[23][527] = 9'b111111111;
assign micromatrizz[23][528] = 9'b111111111;
assign micromatrizz[23][529] = 9'b111111111;
assign micromatrizz[23][530] = 9'b111111111;
assign micromatrizz[23][531] = 9'b111111111;
assign micromatrizz[23][532] = 9'b111111111;
assign micromatrizz[23][533] = 9'b111111111;
assign micromatrizz[23][534] = 9'b111111111;
assign micromatrizz[23][535] = 9'b111111111;
assign micromatrizz[23][536] = 9'b111111111;
assign micromatrizz[23][537] = 9'b111111111;
assign micromatrizz[23][538] = 9'b111111111;
assign micromatrizz[23][539] = 9'b111111111;
assign micromatrizz[23][540] = 9'b111111111;
assign micromatrizz[23][541] = 9'b111111111;
assign micromatrizz[23][542] = 9'b111111111;
assign micromatrizz[23][543] = 9'b111111111;
assign micromatrizz[23][544] = 9'b111111111;
assign micromatrizz[23][545] = 9'b111111111;
assign micromatrizz[23][546] = 9'b111111111;
assign micromatrizz[23][547] = 9'b111111111;
assign micromatrizz[23][548] = 9'b111111111;
assign micromatrizz[23][549] = 9'b111111111;
assign micromatrizz[23][550] = 9'b111111111;
assign micromatrizz[23][551] = 9'b111111111;
assign micromatrizz[23][552] = 9'b111111111;
assign micromatrizz[23][553] = 9'b111111111;
assign micromatrizz[23][554] = 9'b111111111;
assign micromatrizz[23][555] = 9'b111111111;
assign micromatrizz[23][556] = 9'b111111111;
assign micromatrizz[23][557] = 9'b111111111;
assign micromatrizz[23][558] = 9'b111111111;
assign micromatrizz[23][559] = 9'b111111111;
assign micromatrizz[23][560] = 9'b111111111;
assign micromatrizz[23][561] = 9'b111111111;
assign micromatrizz[23][562] = 9'b111111111;
assign micromatrizz[23][563] = 9'b111111111;
assign micromatrizz[23][564] = 9'b111111111;
assign micromatrizz[23][565] = 9'b111111111;
assign micromatrizz[23][566] = 9'b111111111;
assign micromatrizz[23][567] = 9'b111111111;
assign micromatrizz[23][568] = 9'b111111111;
assign micromatrizz[23][569] = 9'b111111111;
assign micromatrizz[23][570] = 9'b111111111;
assign micromatrizz[23][571] = 9'b111111111;
assign micromatrizz[23][572] = 9'b111111111;
assign micromatrizz[23][573] = 9'b111111111;
assign micromatrizz[23][574] = 9'b111111111;
assign micromatrizz[23][575] = 9'b111111111;
assign micromatrizz[23][576] = 9'b111111111;
assign micromatrizz[23][577] = 9'b111111111;
assign micromatrizz[23][578] = 9'b111111111;
assign micromatrizz[23][579] = 9'b111111111;
assign micromatrizz[23][580] = 9'b111111111;
assign micromatrizz[23][581] = 9'b111111111;
assign micromatrizz[23][582] = 9'b111111111;
assign micromatrizz[23][583] = 9'b111111111;
assign micromatrizz[23][584] = 9'b111111111;
assign micromatrizz[23][585] = 9'b111111111;
assign micromatrizz[23][586] = 9'b111111111;
assign micromatrizz[23][587] = 9'b111111111;
assign micromatrizz[23][588] = 9'b111111111;
assign micromatrizz[23][589] = 9'b111111111;
assign micromatrizz[23][590] = 9'b111111111;
assign micromatrizz[23][591] = 9'b111111111;
assign micromatrizz[23][592] = 9'b111111111;
assign micromatrizz[23][593] = 9'b111111111;
assign micromatrizz[23][594] = 9'b111111111;
assign micromatrizz[23][595] = 9'b111111111;
assign micromatrizz[23][596] = 9'b111111111;
assign micromatrizz[23][597] = 9'b111111111;
assign micromatrizz[23][598] = 9'b111111111;
assign micromatrizz[23][599] = 9'b111111111;
assign micromatrizz[23][600] = 9'b111111111;
assign micromatrizz[23][601] = 9'b111111111;
assign micromatrizz[23][602] = 9'b111111111;
assign micromatrizz[23][603] = 9'b111111111;
assign micromatrizz[23][604] = 9'b111111111;
assign micromatrizz[23][605] = 9'b111111111;
assign micromatrizz[23][606] = 9'b111111111;
assign micromatrizz[23][607] = 9'b111111111;
assign micromatrizz[23][608] = 9'b111111111;
assign micromatrizz[23][609] = 9'b111111111;
assign micromatrizz[23][610] = 9'b111111111;
assign micromatrizz[23][611] = 9'b111111111;
assign micromatrizz[23][612] = 9'b111111111;
assign micromatrizz[23][613] = 9'b111111111;
assign micromatrizz[23][614] = 9'b111111111;
assign micromatrizz[23][615] = 9'b111111111;
assign micromatrizz[23][616] = 9'b111111111;
assign micromatrizz[23][617] = 9'b111111111;
assign micromatrizz[23][618] = 9'b111111111;
assign micromatrizz[23][619] = 9'b111111111;
assign micromatrizz[23][620] = 9'b111111111;
assign micromatrizz[23][621] = 9'b111111111;
assign micromatrizz[23][622] = 9'b111111111;
assign micromatrizz[23][623] = 9'b111111111;
assign micromatrizz[23][624] = 9'b111111111;
assign micromatrizz[23][625] = 9'b111111111;
assign micromatrizz[23][626] = 9'b111111111;
assign micromatrizz[23][627] = 9'b111111111;
assign micromatrizz[23][628] = 9'b111111111;
assign micromatrizz[23][629] = 9'b111111111;
assign micromatrizz[23][630] = 9'b111111111;
assign micromatrizz[23][631] = 9'b111111111;
assign micromatrizz[23][632] = 9'b111111111;
assign micromatrizz[23][633] = 9'b111111111;
assign micromatrizz[23][634] = 9'b111111111;
assign micromatrizz[23][635] = 9'b111111111;
assign micromatrizz[23][636] = 9'b111111111;
assign micromatrizz[23][637] = 9'b111111111;
assign micromatrizz[23][638] = 9'b111111111;
assign micromatrizz[23][639] = 9'b111111111;
assign micromatrizz[24][0] = 9'b111111111;
assign micromatrizz[24][1] = 9'b111111111;
assign micromatrizz[24][2] = 9'b111111111;
assign micromatrizz[24][3] = 9'b111111111;
assign micromatrizz[24][4] = 9'b111111111;
assign micromatrizz[24][5] = 9'b111111111;
assign micromatrizz[24][6] = 9'b111111111;
assign micromatrizz[24][7] = 9'b111111111;
assign micromatrizz[24][8] = 9'b111111111;
assign micromatrizz[24][9] = 9'b111111111;
assign micromatrizz[24][10] = 9'b111111111;
assign micromatrizz[24][11] = 9'b111111111;
assign micromatrizz[24][12] = 9'b111111111;
assign micromatrizz[24][13] = 9'b111111111;
assign micromatrizz[24][14] = 9'b111111111;
assign micromatrizz[24][15] = 9'b111111111;
assign micromatrizz[24][16] = 9'b111111111;
assign micromatrizz[24][17] = 9'b111111111;
assign micromatrizz[24][18] = 9'b111111111;
assign micromatrizz[24][19] = 9'b111111111;
assign micromatrizz[24][20] = 9'b111111111;
assign micromatrizz[24][21] = 9'b111111111;
assign micromatrizz[24][22] = 9'b111111111;
assign micromatrizz[24][23] = 9'b111111111;
assign micromatrizz[24][24] = 9'b111111111;
assign micromatrizz[24][25] = 9'b111111111;
assign micromatrizz[24][26] = 9'b111111111;
assign micromatrizz[24][27] = 9'b111111111;
assign micromatrizz[24][28] = 9'b111111111;
assign micromatrizz[24][29] = 9'b111111111;
assign micromatrizz[24][30] = 9'b111111111;
assign micromatrizz[24][31] = 9'b111111111;
assign micromatrizz[24][32] = 9'b111111111;
assign micromatrizz[24][33] = 9'b111111111;
assign micromatrizz[24][34] = 9'b111111111;
assign micromatrizz[24][35] = 9'b111111111;
assign micromatrizz[24][36] = 9'b111111111;
assign micromatrizz[24][37] = 9'b111111111;
assign micromatrizz[24][38] = 9'b111111111;
assign micromatrizz[24][39] = 9'b111111111;
assign micromatrizz[24][40] = 9'b111111111;
assign micromatrizz[24][41] = 9'b111111111;
assign micromatrizz[24][42] = 9'b111111111;
assign micromatrizz[24][43] = 9'b111111111;
assign micromatrizz[24][44] = 9'b111111111;
assign micromatrizz[24][45] = 9'b111111111;
assign micromatrizz[24][46] = 9'b111111111;
assign micromatrizz[24][47] = 9'b111111111;
assign micromatrizz[24][48] = 9'b111111111;
assign micromatrizz[24][49] = 9'b111111111;
assign micromatrizz[24][50] = 9'b111111111;
assign micromatrizz[24][51] = 9'b111111111;
assign micromatrizz[24][52] = 9'b111111111;
assign micromatrizz[24][53] = 9'b111111111;
assign micromatrizz[24][54] = 9'b111111111;
assign micromatrizz[24][55] = 9'b111111111;
assign micromatrizz[24][56] = 9'b111111111;
assign micromatrizz[24][57] = 9'b111111111;
assign micromatrizz[24][58] = 9'b111111111;
assign micromatrizz[24][59] = 9'b111111111;
assign micromatrizz[24][60] = 9'b111111111;
assign micromatrizz[24][61] = 9'b111111111;
assign micromatrizz[24][62] = 9'b111111111;
assign micromatrizz[24][63] = 9'b111111111;
assign micromatrizz[24][64] = 9'b111111111;
assign micromatrizz[24][65] = 9'b111111111;
assign micromatrizz[24][66] = 9'b111111111;
assign micromatrizz[24][67] = 9'b111111111;
assign micromatrizz[24][68] = 9'b111111111;
assign micromatrizz[24][69] = 9'b111111111;
assign micromatrizz[24][70] = 9'b111111111;
assign micromatrizz[24][71] = 9'b111111111;
assign micromatrizz[24][72] = 9'b111111111;
assign micromatrizz[24][73] = 9'b111111111;
assign micromatrizz[24][74] = 9'b111111111;
assign micromatrizz[24][75] = 9'b111111111;
assign micromatrizz[24][76] = 9'b111111111;
assign micromatrizz[24][77] = 9'b111111111;
assign micromatrizz[24][78] = 9'b111111111;
assign micromatrizz[24][79] = 9'b111111111;
assign micromatrizz[24][80] = 9'b111111111;
assign micromatrizz[24][81] = 9'b111111111;
assign micromatrizz[24][82] = 9'b111111111;
assign micromatrizz[24][83] = 9'b111111111;
assign micromatrizz[24][84] = 9'b111111111;
assign micromatrizz[24][85] = 9'b111111111;
assign micromatrizz[24][86] = 9'b111111111;
assign micromatrizz[24][87] = 9'b111111111;
assign micromatrizz[24][88] = 9'b111111111;
assign micromatrizz[24][89] = 9'b111111111;
assign micromatrizz[24][90] = 9'b111111111;
assign micromatrizz[24][91] = 9'b111111111;
assign micromatrizz[24][92] = 9'b111111111;
assign micromatrizz[24][93] = 9'b111111111;
assign micromatrizz[24][94] = 9'b111111111;
assign micromatrizz[24][95] = 9'b111111111;
assign micromatrizz[24][96] = 9'b111111111;
assign micromatrizz[24][97] = 9'b111111111;
assign micromatrizz[24][98] = 9'b111111111;
assign micromatrizz[24][99] = 9'b111111111;
assign micromatrizz[24][100] = 9'b111111111;
assign micromatrizz[24][101] = 9'b111111111;
assign micromatrizz[24][102] = 9'b111111111;
assign micromatrizz[24][103] = 9'b111111111;
assign micromatrizz[24][104] = 9'b111111111;
assign micromatrizz[24][105] = 9'b111111111;
assign micromatrizz[24][106] = 9'b111111111;
assign micromatrizz[24][107] = 9'b111111111;
assign micromatrizz[24][108] = 9'b111111111;
assign micromatrizz[24][109] = 9'b111111111;
assign micromatrizz[24][110] = 9'b111111111;
assign micromatrizz[24][111] = 9'b111111111;
assign micromatrizz[24][112] = 9'b111111111;
assign micromatrizz[24][113] = 9'b111111111;
assign micromatrizz[24][114] = 9'b111111111;
assign micromatrizz[24][115] = 9'b111111111;
assign micromatrizz[24][116] = 9'b111111111;
assign micromatrizz[24][117] = 9'b111111111;
assign micromatrizz[24][118] = 9'b111111111;
assign micromatrizz[24][119] = 9'b111111111;
assign micromatrizz[24][120] = 9'b111111111;
assign micromatrizz[24][121] = 9'b111111111;
assign micromatrizz[24][122] = 9'b111111111;
assign micromatrizz[24][123] = 9'b111111111;
assign micromatrizz[24][124] = 9'b111111111;
assign micromatrizz[24][125] = 9'b111111111;
assign micromatrizz[24][126] = 9'b111111111;
assign micromatrizz[24][127] = 9'b111111111;
assign micromatrizz[24][128] = 9'b111111111;
assign micromatrizz[24][129] = 9'b111111111;
assign micromatrizz[24][130] = 9'b111111111;
assign micromatrizz[24][131] = 9'b111111111;
assign micromatrizz[24][132] = 9'b111111111;
assign micromatrizz[24][133] = 9'b111111111;
assign micromatrizz[24][134] = 9'b111111111;
assign micromatrizz[24][135] = 9'b111111111;
assign micromatrizz[24][136] = 9'b111111111;
assign micromatrizz[24][137] = 9'b111111111;
assign micromatrizz[24][138] = 9'b111111111;
assign micromatrizz[24][139] = 9'b111111111;
assign micromatrizz[24][140] = 9'b111111111;
assign micromatrizz[24][141] = 9'b111111111;
assign micromatrizz[24][142] = 9'b111111111;
assign micromatrizz[24][143] = 9'b111111111;
assign micromatrizz[24][144] = 9'b111111111;
assign micromatrizz[24][145] = 9'b111111111;
assign micromatrizz[24][146] = 9'b111111111;
assign micromatrizz[24][147] = 9'b111111111;
assign micromatrizz[24][148] = 9'b111111111;
assign micromatrizz[24][149] = 9'b111111111;
assign micromatrizz[24][150] = 9'b111111111;
assign micromatrizz[24][151] = 9'b111111111;
assign micromatrizz[24][152] = 9'b111111111;
assign micromatrizz[24][153] = 9'b111111111;
assign micromatrizz[24][154] = 9'b111111111;
assign micromatrizz[24][155] = 9'b111111111;
assign micromatrizz[24][156] = 9'b111111111;
assign micromatrizz[24][157] = 9'b111111111;
assign micromatrizz[24][158] = 9'b111111111;
assign micromatrizz[24][159] = 9'b111111111;
assign micromatrizz[24][160] = 9'b111111111;
assign micromatrizz[24][161] = 9'b111111111;
assign micromatrizz[24][162] = 9'b111111111;
assign micromatrizz[24][163] = 9'b111111111;
assign micromatrizz[24][164] = 9'b111111111;
assign micromatrizz[24][165] = 9'b111111111;
assign micromatrizz[24][166] = 9'b111111111;
assign micromatrizz[24][167] = 9'b111111111;
assign micromatrizz[24][168] = 9'b111111111;
assign micromatrizz[24][169] = 9'b111111111;
assign micromatrizz[24][170] = 9'b111111111;
assign micromatrizz[24][171] = 9'b111111111;
assign micromatrizz[24][172] = 9'b111111111;
assign micromatrizz[24][173] = 9'b111111111;
assign micromatrizz[24][174] = 9'b111111111;
assign micromatrizz[24][175] = 9'b111111111;
assign micromatrizz[24][176] = 9'b111111111;
assign micromatrizz[24][177] = 9'b111111111;
assign micromatrizz[24][178] = 9'b111111111;
assign micromatrizz[24][179] = 9'b111111111;
assign micromatrizz[24][180] = 9'b111111111;
assign micromatrizz[24][181] = 9'b111111111;
assign micromatrizz[24][182] = 9'b111111111;
assign micromatrizz[24][183] = 9'b111111111;
assign micromatrizz[24][184] = 9'b111111111;
assign micromatrizz[24][185] = 9'b111111111;
assign micromatrizz[24][186] = 9'b111111111;
assign micromatrizz[24][187] = 9'b111111111;
assign micromatrizz[24][188] = 9'b111111111;
assign micromatrizz[24][189] = 9'b111111111;
assign micromatrizz[24][190] = 9'b111111111;
assign micromatrizz[24][191] = 9'b111111111;
assign micromatrizz[24][192] = 9'b111111111;
assign micromatrizz[24][193] = 9'b111111111;
assign micromatrizz[24][194] = 9'b111111111;
assign micromatrizz[24][195] = 9'b111111111;
assign micromatrizz[24][196] = 9'b111111111;
assign micromatrizz[24][197] = 9'b111111111;
assign micromatrizz[24][198] = 9'b111111111;
assign micromatrizz[24][199] = 9'b111111111;
assign micromatrizz[24][200] = 9'b111111111;
assign micromatrizz[24][201] = 9'b111111111;
assign micromatrizz[24][202] = 9'b111111111;
assign micromatrizz[24][203] = 9'b111111111;
assign micromatrizz[24][204] = 9'b111111111;
assign micromatrizz[24][205] = 9'b111111111;
assign micromatrizz[24][206] = 9'b111111111;
assign micromatrizz[24][207] = 9'b111111111;
assign micromatrizz[24][208] = 9'b111111111;
assign micromatrizz[24][209] = 9'b111111111;
assign micromatrizz[24][210] = 9'b111111111;
assign micromatrizz[24][211] = 9'b111111111;
assign micromatrizz[24][212] = 9'b111111111;
assign micromatrizz[24][213] = 9'b111111111;
assign micromatrizz[24][214] = 9'b111111111;
assign micromatrizz[24][215] = 9'b111111111;
assign micromatrizz[24][216] = 9'b111111111;
assign micromatrizz[24][217] = 9'b111111111;
assign micromatrizz[24][218] = 9'b111111111;
assign micromatrizz[24][219] = 9'b111111111;
assign micromatrizz[24][220] = 9'b111111111;
assign micromatrizz[24][221] = 9'b111111111;
assign micromatrizz[24][222] = 9'b111111111;
assign micromatrizz[24][223] = 9'b111111111;
assign micromatrizz[24][224] = 9'b111111111;
assign micromatrizz[24][225] = 9'b111111111;
assign micromatrizz[24][226] = 9'b111111111;
assign micromatrizz[24][227] = 9'b111111111;
assign micromatrizz[24][228] = 9'b111111111;
assign micromatrizz[24][229] = 9'b111111111;
assign micromatrizz[24][230] = 9'b111111111;
assign micromatrizz[24][231] = 9'b111111111;
assign micromatrizz[24][232] = 9'b111111111;
assign micromatrizz[24][233] = 9'b111111111;
assign micromatrizz[24][234] = 9'b111111111;
assign micromatrizz[24][235] = 9'b111111111;
assign micromatrizz[24][236] = 9'b111111111;
assign micromatrizz[24][237] = 9'b111111111;
assign micromatrizz[24][238] = 9'b111111111;
assign micromatrizz[24][239] = 9'b111111111;
assign micromatrizz[24][240] = 9'b111111111;
assign micromatrizz[24][241] = 9'b111111111;
assign micromatrizz[24][242] = 9'b111111111;
assign micromatrizz[24][243] = 9'b111111111;
assign micromatrizz[24][244] = 9'b111111111;
assign micromatrizz[24][245] = 9'b111111111;
assign micromatrizz[24][246] = 9'b111111111;
assign micromatrizz[24][247] = 9'b111111111;
assign micromatrizz[24][248] = 9'b111111111;
assign micromatrizz[24][249] = 9'b111111111;
assign micromatrizz[24][250] = 9'b111111111;
assign micromatrizz[24][251] = 9'b111111111;
assign micromatrizz[24][252] = 9'b111111111;
assign micromatrizz[24][253] = 9'b111111111;
assign micromatrizz[24][254] = 9'b111111111;
assign micromatrizz[24][255] = 9'b111111111;
assign micromatrizz[24][256] = 9'b111111111;
assign micromatrizz[24][257] = 9'b111111111;
assign micromatrizz[24][258] = 9'b111111111;
assign micromatrizz[24][259] = 9'b111111111;
assign micromatrizz[24][260] = 9'b111111111;
assign micromatrizz[24][261] = 9'b111111111;
assign micromatrizz[24][262] = 9'b111111111;
assign micromatrizz[24][263] = 9'b111111111;
assign micromatrizz[24][264] = 9'b111111111;
assign micromatrizz[24][265] = 9'b111111111;
assign micromatrizz[24][266] = 9'b111111111;
assign micromatrizz[24][267] = 9'b111111111;
assign micromatrizz[24][268] = 9'b111111111;
assign micromatrizz[24][269] = 9'b111111111;
assign micromatrizz[24][270] = 9'b111110010;
assign micromatrizz[24][271] = 9'b111110010;
assign micromatrizz[24][272] = 9'b111110010;
assign micromatrizz[24][273] = 9'b111110010;
assign micromatrizz[24][274] = 9'b111110010;
assign micromatrizz[24][275] = 9'b111110011;
assign micromatrizz[24][276] = 9'b111110011;
assign micromatrizz[24][277] = 9'b111110011;
assign micromatrizz[24][278] = 9'b111110011;
assign micromatrizz[24][279] = 9'b111111111;
assign micromatrizz[24][280] = 9'b111111111;
assign micromatrizz[24][281] = 9'b111111111;
assign micromatrizz[24][282] = 9'b111111111;
assign micromatrizz[24][283] = 9'b111111111;
assign micromatrizz[24][284] = 9'b111111111;
assign micromatrizz[24][285] = 9'b111111111;
assign micromatrizz[24][286] = 9'b111111111;
assign micromatrizz[24][287] = 9'b111111111;
assign micromatrizz[24][288] = 9'b111111111;
assign micromatrizz[24][289] = 9'b111111111;
assign micromatrizz[24][290] = 9'b111111111;
assign micromatrizz[24][291] = 9'b111111111;
assign micromatrizz[24][292] = 9'b111110111;
assign micromatrizz[24][293] = 9'b111110010;
assign micromatrizz[24][294] = 9'b111110011;
assign micromatrizz[24][295] = 9'b111110011;
assign micromatrizz[24][296] = 9'b111110011;
assign micromatrizz[24][297] = 9'b111110111;
assign micromatrizz[24][298] = 9'b111111111;
assign micromatrizz[24][299] = 9'b111111111;
assign micromatrizz[24][300] = 9'b111111111;
assign micromatrizz[24][301] = 9'b111111111;
assign micromatrizz[24][302] = 9'b111111111;
assign micromatrizz[24][303] = 9'b111110111;
assign micromatrizz[24][304] = 9'b111111111;
assign micromatrizz[24][305] = 9'b111111111;
assign micromatrizz[24][306] = 9'b111111111;
assign micromatrizz[24][307] = 9'b111111111;
assign micromatrizz[24][308] = 9'b111111111;
assign micromatrizz[24][309] = 9'b111110010;
assign micromatrizz[24][310] = 9'b111110010;
assign micromatrizz[24][311] = 9'b111110011;
assign micromatrizz[24][312] = 9'b111110011;
assign micromatrizz[24][313] = 9'b111110011;
assign micromatrizz[24][314] = 9'b111110111;
assign micromatrizz[24][315] = 9'b111111111;
assign micromatrizz[24][316] = 9'b111111111;
assign micromatrizz[24][317] = 9'b111111111;
assign micromatrizz[24][318] = 9'b111111111;
assign micromatrizz[24][319] = 9'b111111111;
assign micromatrizz[24][320] = 9'b111111111;
assign micromatrizz[24][321] = 9'b111111111;
assign micromatrizz[24][322] = 9'b111111111;
assign micromatrizz[24][323] = 9'b111111111;
assign micromatrizz[24][324] = 9'b111111111;
assign micromatrizz[24][325] = 9'b111111111;
assign micromatrizz[24][326] = 9'b111111111;
assign micromatrizz[24][327] = 9'b111111111;
assign micromatrizz[24][328] = 9'b111111111;
assign micromatrizz[24][329] = 9'b111111111;
assign micromatrizz[24][330] = 9'b111111111;
assign micromatrizz[24][331] = 9'b111111111;
assign micromatrizz[24][332] = 9'b111111111;
assign micromatrizz[24][333] = 9'b111111111;
assign micromatrizz[24][334] = 9'b111111111;
assign micromatrizz[24][335] = 9'b111111111;
assign micromatrizz[24][336] = 9'b111111111;
assign micromatrizz[24][337] = 9'b111111111;
assign micromatrizz[24][338] = 9'b111111111;
assign micromatrizz[24][339] = 9'b111111111;
assign micromatrizz[24][340] = 9'b111111111;
assign micromatrizz[24][341] = 9'b111111111;
assign micromatrizz[24][342] = 9'b111111111;
assign micromatrizz[24][343] = 9'b111111111;
assign micromatrizz[24][344] = 9'b111111111;
assign micromatrizz[24][345] = 9'b111111111;
assign micromatrizz[24][346] = 9'b111111111;
assign micromatrizz[24][347] = 9'b111111111;
assign micromatrizz[24][348] = 9'b111111111;
assign micromatrizz[24][349] = 9'b111111111;
assign micromatrizz[24][350] = 9'b111111111;
assign micromatrizz[24][351] = 9'b111111111;
assign micromatrizz[24][352] = 9'b111111111;
assign micromatrizz[24][353] = 9'b111111111;
assign micromatrizz[24][354] = 9'b111111111;
assign micromatrizz[24][355] = 9'b111111111;
assign micromatrizz[24][356] = 9'b111111111;
assign micromatrizz[24][357] = 9'b111111111;
assign micromatrizz[24][358] = 9'b111111111;
assign micromatrizz[24][359] = 9'b111111111;
assign micromatrizz[24][360] = 9'b111111111;
assign micromatrizz[24][361] = 9'b111111111;
assign micromatrizz[24][362] = 9'b111111111;
assign micromatrizz[24][363] = 9'b111111111;
assign micromatrizz[24][364] = 9'b111111111;
assign micromatrizz[24][365] = 9'b111111111;
assign micromatrizz[24][366] = 9'b111111111;
assign micromatrizz[24][367] = 9'b111111111;
assign micromatrizz[24][368] = 9'b111111111;
assign micromatrizz[24][369] = 9'b111111111;
assign micromatrizz[24][370] = 9'b111111111;
assign micromatrizz[24][371] = 9'b111111111;
assign micromatrizz[24][372] = 9'b111111111;
assign micromatrizz[24][373] = 9'b111111111;
assign micromatrizz[24][374] = 9'b111111111;
assign micromatrizz[24][375] = 9'b111111111;
assign micromatrizz[24][376] = 9'b111111111;
assign micromatrizz[24][377] = 9'b111111111;
assign micromatrizz[24][378] = 9'b111111111;
assign micromatrizz[24][379] = 9'b111111111;
assign micromatrizz[24][380] = 9'b111111111;
assign micromatrizz[24][381] = 9'b111111111;
assign micromatrizz[24][382] = 9'b111111111;
assign micromatrizz[24][383] = 9'b111111111;
assign micromatrizz[24][384] = 9'b111111111;
assign micromatrizz[24][385] = 9'b111111111;
assign micromatrizz[24][386] = 9'b111111111;
assign micromatrizz[24][387] = 9'b111111111;
assign micromatrizz[24][388] = 9'b111111111;
assign micromatrizz[24][389] = 9'b111111111;
assign micromatrizz[24][390] = 9'b111111111;
assign micromatrizz[24][391] = 9'b111111111;
assign micromatrizz[24][392] = 9'b111111111;
assign micromatrizz[24][393] = 9'b111111111;
assign micromatrizz[24][394] = 9'b111111111;
assign micromatrizz[24][395] = 9'b111111111;
assign micromatrizz[24][396] = 9'b111111111;
assign micromatrizz[24][397] = 9'b111111111;
assign micromatrizz[24][398] = 9'b111111111;
assign micromatrizz[24][399] = 9'b111111111;
assign micromatrizz[24][400] = 9'b111111111;
assign micromatrizz[24][401] = 9'b111111111;
assign micromatrizz[24][402] = 9'b111111111;
assign micromatrizz[24][403] = 9'b111111111;
assign micromatrizz[24][404] = 9'b111111111;
assign micromatrizz[24][405] = 9'b111111111;
assign micromatrizz[24][406] = 9'b111111111;
assign micromatrizz[24][407] = 9'b111111111;
assign micromatrizz[24][408] = 9'b111111111;
assign micromatrizz[24][409] = 9'b111111111;
assign micromatrizz[24][410] = 9'b111111111;
assign micromatrizz[24][411] = 9'b111111111;
assign micromatrizz[24][412] = 9'b111111111;
assign micromatrizz[24][413] = 9'b111111111;
assign micromatrizz[24][414] = 9'b111111111;
assign micromatrizz[24][415] = 9'b111111111;
assign micromatrizz[24][416] = 9'b111111111;
assign micromatrizz[24][417] = 9'b111111111;
assign micromatrizz[24][418] = 9'b111111111;
assign micromatrizz[24][419] = 9'b111111111;
assign micromatrizz[24][420] = 9'b111111111;
assign micromatrizz[24][421] = 9'b111111111;
assign micromatrizz[24][422] = 9'b111111111;
assign micromatrizz[24][423] = 9'b111111111;
assign micromatrizz[24][424] = 9'b111111111;
assign micromatrizz[24][425] = 9'b111111111;
assign micromatrizz[24][426] = 9'b111111111;
assign micromatrizz[24][427] = 9'b111111111;
assign micromatrizz[24][428] = 9'b111111111;
assign micromatrizz[24][429] = 9'b111111111;
assign micromatrizz[24][430] = 9'b111111111;
assign micromatrizz[24][431] = 9'b111111111;
assign micromatrizz[24][432] = 9'b111111111;
assign micromatrizz[24][433] = 9'b111111111;
assign micromatrizz[24][434] = 9'b111111111;
assign micromatrizz[24][435] = 9'b111111111;
assign micromatrizz[24][436] = 9'b111111111;
assign micromatrizz[24][437] = 9'b111111111;
assign micromatrizz[24][438] = 9'b111111111;
assign micromatrizz[24][439] = 9'b111111111;
assign micromatrizz[24][440] = 9'b111111111;
assign micromatrizz[24][441] = 9'b111111111;
assign micromatrizz[24][442] = 9'b111111111;
assign micromatrizz[24][443] = 9'b111111111;
assign micromatrizz[24][444] = 9'b111111111;
assign micromatrizz[24][445] = 9'b111111111;
assign micromatrizz[24][446] = 9'b111111111;
assign micromatrizz[24][447] = 9'b111111111;
assign micromatrizz[24][448] = 9'b111111111;
assign micromatrizz[24][449] = 9'b111111111;
assign micromatrizz[24][450] = 9'b111111111;
assign micromatrizz[24][451] = 9'b111111111;
assign micromatrizz[24][452] = 9'b111111111;
assign micromatrizz[24][453] = 9'b111111111;
assign micromatrizz[24][454] = 9'b111111111;
assign micromatrizz[24][455] = 9'b111111111;
assign micromatrizz[24][456] = 9'b111111111;
assign micromatrizz[24][457] = 9'b111111111;
assign micromatrizz[24][458] = 9'b111111111;
assign micromatrizz[24][459] = 9'b111111111;
assign micromatrizz[24][460] = 9'b111111111;
assign micromatrizz[24][461] = 9'b111111111;
assign micromatrizz[24][462] = 9'b111111111;
assign micromatrizz[24][463] = 9'b111111111;
assign micromatrizz[24][464] = 9'b111111111;
assign micromatrizz[24][465] = 9'b111111111;
assign micromatrizz[24][466] = 9'b111111111;
assign micromatrizz[24][467] = 9'b111111111;
assign micromatrizz[24][468] = 9'b111111111;
assign micromatrizz[24][469] = 9'b111111111;
assign micromatrizz[24][470] = 9'b111111111;
assign micromatrizz[24][471] = 9'b111111111;
assign micromatrizz[24][472] = 9'b111111111;
assign micromatrizz[24][473] = 9'b111111111;
assign micromatrizz[24][474] = 9'b111111111;
assign micromatrizz[24][475] = 9'b111111111;
assign micromatrizz[24][476] = 9'b111111111;
assign micromatrizz[24][477] = 9'b111111111;
assign micromatrizz[24][478] = 9'b111111111;
assign micromatrizz[24][479] = 9'b111111111;
assign micromatrizz[24][480] = 9'b111111111;
assign micromatrizz[24][481] = 9'b111111111;
assign micromatrizz[24][482] = 9'b111111111;
assign micromatrizz[24][483] = 9'b111111111;
assign micromatrizz[24][484] = 9'b111111111;
assign micromatrizz[24][485] = 9'b111111111;
assign micromatrizz[24][486] = 9'b111111111;
assign micromatrizz[24][487] = 9'b111111111;
assign micromatrizz[24][488] = 9'b111111111;
assign micromatrizz[24][489] = 9'b111111111;
assign micromatrizz[24][490] = 9'b111111111;
assign micromatrizz[24][491] = 9'b111111111;
assign micromatrizz[24][492] = 9'b111111111;
assign micromatrizz[24][493] = 9'b111111111;
assign micromatrizz[24][494] = 9'b111111111;
assign micromatrizz[24][495] = 9'b111111111;
assign micromatrizz[24][496] = 9'b111111111;
assign micromatrizz[24][497] = 9'b111111111;
assign micromatrizz[24][498] = 9'b111111111;
assign micromatrizz[24][499] = 9'b111111111;
assign micromatrizz[24][500] = 9'b111111111;
assign micromatrizz[24][501] = 9'b111111111;
assign micromatrizz[24][502] = 9'b111111111;
assign micromatrizz[24][503] = 9'b111111111;
assign micromatrizz[24][504] = 9'b111111111;
assign micromatrizz[24][505] = 9'b111111111;
assign micromatrizz[24][506] = 9'b111111111;
assign micromatrizz[24][507] = 9'b111111111;
assign micromatrizz[24][508] = 9'b111111111;
assign micromatrizz[24][509] = 9'b111111111;
assign micromatrizz[24][510] = 9'b111111111;
assign micromatrizz[24][511] = 9'b111111111;
assign micromatrizz[24][512] = 9'b111111111;
assign micromatrizz[24][513] = 9'b111111111;
assign micromatrizz[24][514] = 9'b111111111;
assign micromatrizz[24][515] = 9'b111111111;
assign micromatrizz[24][516] = 9'b111111111;
assign micromatrizz[24][517] = 9'b111111111;
assign micromatrizz[24][518] = 9'b111111111;
assign micromatrizz[24][519] = 9'b111111111;
assign micromatrizz[24][520] = 9'b111111111;
assign micromatrizz[24][521] = 9'b111111111;
assign micromatrizz[24][522] = 9'b111111111;
assign micromatrizz[24][523] = 9'b111111111;
assign micromatrizz[24][524] = 9'b111111111;
assign micromatrizz[24][525] = 9'b111111111;
assign micromatrizz[24][526] = 9'b111111111;
assign micromatrizz[24][527] = 9'b111111111;
assign micromatrizz[24][528] = 9'b111111111;
assign micromatrizz[24][529] = 9'b111111111;
assign micromatrizz[24][530] = 9'b111111111;
assign micromatrizz[24][531] = 9'b111111111;
assign micromatrizz[24][532] = 9'b111111111;
assign micromatrizz[24][533] = 9'b111111111;
assign micromatrizz[24][534] = 9'b111111111;
assign micromatrizz[24][535] = 9'b111111111;
assign micromatrizz[24][536] = 9'b111111111;
assign micromatrizz[24][537] = 9'b111111111;
assign micromatrizz[24][538] = 9'b111111111;
assign micromatrizz[24][539] = 9'b111111111;
assign micromatrizz[24][540] = 9'b111111111;
assign micromatrizz[24][541] = 9'b111111111;
assign micromatrizz[24][542] = 9'b111111111;
assign micromatrizz[24][543] = 9'b111111111;
assign micromatrizz[24][544] = 9'b111111111;
assign micromatrizz[24][545] = 9'b111111111;
assign micromatrizz[24][546] = 9'b111111111;
assign micromatrizz[24][547] = 9'b111111111;
assign micromatrizz[24][548] = 9'b111111111;
assign micromatrizz[24][549] = 9'b111111111;
assign micromatrizz[24][550] = 9'b111111111;
assign micromatrizz[24][551] = 9'b111111111;
assign micromatrizz[24][552] = 9'b111111111;
assign micromatrizz[24][553] = 9'b111111111;
assign micromatrizz[24][554] = 9'b111111111;
assign micromatrizz[24][555] = 9'b111111111;
assign micromatrizz[24][556] = 9'b111111111;
assign micromatrizz[24][557] = 9'b111111111;
assign micromatrizz[24][558] = 9'b111111111;
assign micromatrizz[24][559] = 9'b111111111;
assign micromatrizz[24][560] = 9'b111111111;
assign micromatrizz[24][561] = 9'b111111111;
assign micromatrizz[24][562] = 9'b111111111;
assign micromatrizz[24][563] = 9'b111111111;
assign micromatrizz[24][564] = 9'b111111111;
assign micromatrizz[24][565] = 9'b111111111;
assign micromatrizz[24][566] = 9'b111111111;
assign micromatrizz[24][567] = 9'b111111111;
assign micromatrizz[24][568] = 9'b111111111;
assign micromatrizz[24][569] = 9'b111111111;
assign micromatrizz[24][570] = 9'b111111111;
assign micromatrizz[24][571] = 9'b111111111;
assign micromatrizz[24][572] = 9'b111111111;
assign micromatrizz[24][573] = 9'b111111111;
assign micromatrizz[24][574] = 9'b111111111;
assign micromatrizz[24][575] = 9'b111111111;
assign micromatrizz[24][576] = 9'b111111111;
assign micromatrizz[24][577] = 9'b111111111;
assign micromatrizz[24][578] = 9'b111111111;
assign micromatrizz[24][579] = 9'b111111111;
assign micromatrizz[24][580] = 9'b111111111;
assign micromatrizz[24][581] = 9'b111111111;
assign micromatrizz[24][582] = 9'b111111111;
assign micromatrizz[24][583] = 9'b111111111;
assign micromatrizz[24][584] = 9'b111111111;
assign micromatrizz[24][585] = 9'b111111111;
assign micromatrizz[24][586] = 9'b111111111;
assign micromatrizz[24][587] = 9'b111111111;
assign micromatrizz[24][588] = 9'b111111111;
assign micromatrizz[24][589] = 9'b111111111;
assign micromatrizz[24][590] = 9'b111111111;
assign micromatrizz[24][591] = 9'b111111111;
assign micromatrizz[24][592] = 9'b111111111;
assign micromatrizz[24][593] = 9'b111111111;
assign micromatrizz[24][594] = 9'b111111111;
assign micromatrizz[24][595] = 9'b111111111;
assign micromatrizz[24][596] = 9'b111111111;
assign micromatrizz[24][597] = 9'b111111111;
assign micromatrizz[24][598] = 9'b111111111;
assign micromatrizz[24][599] = 9'b111111111;
assign micromatrizz[24][600] = 9'b111111111;
assign micromatrizz[24][601] = 9'b111111111;
assign micromatrizz[24][602] = 9'b111111111;
assign micromatrizz[24][603] = 9'b111111111;
assign micromatrizz[24][604] = 9'b111111111;
assign micromatrizz[24][605] = 9'b111111111;
assign micromatrizz[24][606] = 9'b111111111;
assign micromatrizz[24][607] = 9'b111111111;
assign micromatrizz[24][608] = 9'b111111111;
assign micromatrizz[24][609] = 9'b111111111;
assign micromatrizz[24][610] = 9'b111111111;
assign micromatrizz[24][611] = 9'b111111111;
assign micromatrizz[24][612] = 9'b111111111;
assign micromatrizz[24][613] = 9'b111111111;
assign micromatrizz[24][614] = 9'b111111111;
assign micromatrizz[24][615] = 9'b111111111;
assign micromatrizz[24][616] = 9'b111111111;
assign micromatrizz[24][617] = 9'b111111111;
assign micromatrizz[24][618] = 9'b111111111;
assign micromatrizz[24][619] = 9'b111111111;
assign micromatrizz[24][620] = 9'b111111111;
assign micromatrizz[24][621] = 9'b111111111;
assign micromatrizz[24][622] = 9'b111111111;
assign micromatrizz[24][623] = 9'b111111111;
assign micromatrizz[24][624] = 9'b111111111;
assign micromatrizz[24][625] = 9'b111111111;
assign micromatrizz[24][626] = 9'b111111111;
assign micromatrizz[24][627] = 9'b111111111;
assign micromatrizz[24][628] = 9'b111111111;
assign micromatrizz[24][629] = 9'b111111111;
assign micromatrizz[24][630] = 9'b111111111;
assign micromatrizz[24][631] = 9'b111111111;
assign micromatrizz[24][632] = 9'b111111111;
assign micromatrizz[24][633] = 9'b111111111;
assign micromatrizz[24][634] = 9'b111111111;
assign micromatrizz[24][635] = 9'b111111111;
assign micromatrizz[24][636] = 9'b111111111;
assign micromatrizz[24][637] = 9'b111111111;
assign micromatrizz[24][638] = 9'b111111111;
assign micromatrizz[24][639] = 9'b111111111;
assign micromatrizz[25][0] = 9'b111111111;
assign micromatrizz[25][1] = 9'b111111111;
assign micromatrizz[25][2] = 9'b111111111;
assign micromatrizz[25][3] = 9'b111111111;
assign micromatrizz[25][4] = 9'b111111111;
assign micromatrizz[25][5] = 9'b111111111;
assign micromatrizz[25][6] = 9'b111111111;
assign micromatrizz[25][7] = 9'b111111111;
assign micromatrizz[25][8] = 9'b111111111;
assign micromatrizz[25][9] = 9'b111111111;
assign micromatrizz[25][10] = 9'b111111111;
assign micromatrizz[25][11] = 9'b111111111;
assign micromatrizz[25][12] = 9'b111111111;
assign micromatrizz[25][13] = 9'b111111111;
assign micromatrizz[25][14] = 9'b111111111;
assign micromatrizz[25][15] = 9'b111111111;
assign micromatrizz[25][16] = 9'b111111111;
assign micromatrizz[25][17] = 9'b111111111;
assign micromatrizz[25][18] = 9'b111111111;
assign micromatrizz[25][19] = 9'b111111111;
assign micromatrizz[25][20] = 9'b111111111;
assign micromatrizz[25][21] = 9'b111111111;
assign micromatrizz[25][22] = 9'b111111111;
assign micromatrizz[25][23] = 9'b111111111;
assign micromatrizz[25][24] = 9'b111111111;
assign micromatrizz[25][25] = 9'b111111111;
assign micromatrizz[25][26] = 9'b111111111;
assign micromatrizz[25][27] = 9'b111111111;
assign micromatrizz[25][28] = 9'b111111111;
assign micromatrizz[25][29] = 9'b111111111;
assign micromatrizz[25][30] = 9'b111111111;
assign micromatrizz[25][31] = 9'b111111111;
assign micromatrizz[25][32] = 9'b111111111;
assign micromatrizz[25][33] = 9'b111111111;
assign micromatrizz[25][34] = 9'b111111111;
assign micromatrizz[25][35] = 9'b111111111;
assign micromatrizz[25][36] = 9'b111111111;
assign micromatrizz[25][37] = 9'b111111111;
assign micromatrizz[25][38] = 9'b111111111;
assign micromatrizz[25][39] = 9'b111111111;
assign micromatrizz[25][40] = 9'b111111111;
assign micromatrizz[25][41] = 9'b111111111;
assign micromatrizz[25][42] = 9'b111111111;
assign micromatrizz[25][43] = 9'b111111111;
assign micromatrizz[25][44] = 9'b111111111;
assign micromatrizz[25][45] = 9'b111111111;
assign micromatrizz[25][46] = 9'b111111111;
assign micromatrizz[25][47] = 9'b111111111;
assign micromatrizz[25][48] = 9'b111111111;
assign micromatrizz[25][49] = 9'b111111111;
assign micromatrizz[25][50] = 9'b111111111;
assign micromatrizz[25][51] = 9'b111111111;
assign micromatrizz[25][52] = 9'b111111111;
assign micromatrizz[25][53] = 9'b111111111;
assign micromatrizz[25][54] = 9'b111111111;
assign micromatrizz[25][55] = 9'b111111111;
assign micromatrizz[25][56] = 9'b111111111;
assign micromatrizz[25][57] = 9'b111111111;
assign micromatrizz[25][58] = 9'b111111111;
assign micromatrizz[25][59] = 9'b111111111;
assign micromatrizz[25][60] = 9'b111111111;
assign micromatrizz[25][61] = 9'b111111111;
assign micromatrizz[25][62] = 9'b111111111;
assign micromatrizz[25][63] = 9'b111111111;
assign micromatrizz[25][64] = 9'b111111111;
assign micromatrizz[25][65] = 9'b111111111;
assign micromatrizz[25][66] = 9'b111111111;
assign micromatrizz[25][67] = 9'b111111111;
assign micromatrizz[25][68] = 9'b111111111;
assign micromatrizz[25][69] = 9'b111111111;
assign micromatrizz[25][70] = 9'b111111111;
assign micromatrizz[25][71] = 9'b111111111;
assign micromatrizz[25][72] = 9'b111111111;
assign micromatrizz[25][73] = 9'b111111111;
assign micromatrizz[25][74] = 9'b111111111;
assign micromatrizz[25][75] = 9'b111111111;
assign micromatrizz[25][76] = 9'b111111111;
assign micromatrizz[25][77] = 9'b111111111;
assign micromatrizz[25][78] = 9'b111111111;
assign micromatrizz[25][79] = 9'b111111111;
assign micromatrizz[25][80] = 9'b111111111;
assign micromatrizz[25][81] = 9'b111111111;
assign micromatrizz[25][82] = 9'b111111111;
assign micromatrizz[25][83] = 9'b111111111;
assign micromatrizz[25][84] = 9'b111111111;
assign micromatrizz[25][85] = 9'b111111111;
assign micromatrizz[25][86] = 9'b111111111;
assign micromatrizz[25][87] = 9'b111111111;
assign micromatrizz[25][88] = 9'b111111111;
assign micromatrizz[25][89] = 9'b111111111;
assign micromatrizz[25][90] = 9'b111111111;
assign micromatrizz[25][91] = 9'b111111111;
assign micromatrizz[25][92] = 9'b111111111;
assign micromatrizz[25][93] = 9'b111111111;
assign micromatrizz[25][94] = 9'b111111111;
assign micromatrizz[25][95] = 9'b111111111;
assign micromatrizz[25][96] = 9'b111111111;
assign micromatrizz[25][97] = 9'b111111111;
assign micromatrizz[25][98] = 9'b111111111;
assign micromatrizz[25][99] = 9'b111111111;
assign micromatrizz[25][100] = 9'b111111111;
assign micromatrizz[25][101] = 9'b111111111;
assign micromatrizz[25][102] = 9'b111111111;
assign micromatrizz[25][103] = 9'b111111111;
assign micromatrizz[25][104] = 9'b111111111;
assign micromatrizz[25][105] = 9'b111111111;
assign micromatrizz[25][106] = 9'b111111111;
assign micromatrizz[25][107] = 9'b111111111;
assign micromatrizz[25][108] = 9'b111111111;
assign micromatrizz[25][109] = 9'b111111111;
assign micromatrizz[25][110] = 9'b111111111;
assign micromatrizz[25][111] = 9'b111111111;
assign micromatrizz[25][112] = 9'b111111111;
assign micromatrizz[25][113] = 9'b111111111;
assign micromatrizz[25][114] = 9'b111111111;
assign micromatrizz[25][115] = 9'b111111111;
assign micromatrizz[25][116] = 9'b111111111;
assign micromatrizz[25][117] = 9'b111111111;
assign micromatrizz[25][118] = 9'b111111111;
assign micromatrizz[25][119] = 9'b111111111;
assign micromatrizz[25][120] = 9'b111111111;
assign micromatrizz[25][121] = 9'b111111111;
assign micromatrizz[25][122] = 9'b111111111;
assign micromatrizz[25][123] = 9'b111111111;
assign micromatrizz[25][124] = 9'b111111111;
assign micromatrizz[25][125] = 9'b111111111;
assign micromatrizz[25][126] = 9'b111111111;
assign micromatrizz[25][127] = 9'b111111111;
assign micromatrizz[25][128] = 9'b111111111;
assign micromatrizz[25][129] = 9'b111111111;
assign micromatrizz[25][130] = 9'b111111111;
assign micromatrizz[25][131] = 9'b111111111;
assign micromatrizz[25][132] = 9'b111111111;
assign micromatrizz[25][133] = 9'b111111111;
assign micromatrizz[25][134] = 9'b111111111;
assign micromatrizz[25][135] = 9'b111111111;
assign micromatrizz[25][136] = 9'b111111111;
assign micromatrizz[25][137] = 9'b111111111;
assign micromatrizz[25][138] = 9'b111111111;
assign micromatrizz[25][139] = 9'b111111111;
assign micromatrizz[25][140] = 9'b111111111;
assign micromatrizz[25][141] = 9'b111111111;
assign micromatrizz[25][142] = 9'b111111111;
assign micromatrizz[25][143] = 9'b111111111;
assign micromatrizz[25][144] = 9'b111111111;
assign micromatrizz[25][145] = 9'b111111111;
assign micromatrizz[25][146] = 9'b111111111;
assign micromatrizz[25][147] = 9'b111111111;
assign micromatrizz[25][148] = 9'b111111111;
assign micromatrizz[25][149] = 9'b111111111;
assign micromatrizz[25][150] = 9'b111111111;
assign micromatrizz[25][151] = 9'b111111111;
assign micromatrizz[25][152] = 9'b111111111;
assign micromatrizz[25][153] = 9'b111111111;
assign micromatrizz[25][154] = 9'b111111111;
assign micromatrizz[25][155] = 9'b111111111;
assign micromatrizz[25][156] = 9'b111111111;
assign micromatrizz[25][157] = 9'b111111111;
assign micromatrizz[25][158] = 9'b111111111;
assign micromatrizz[25][159] = 9'b111111111;
assign micromatrizz[25][160] = 9'b111111111;
assign micromatrizz[25][161] = 9'b111111111;
assign micromatrizz[25][162] = 9'b111111111;
assign micromatrizz[25][163] = 9'b111111111;
assign micromatrizz[25][164] = 9'b111111111;
assign micromatrizz[25][165] = 9'b111111111;
assign micromatrizz[25][166] = 9'b111111111;
assign micromatrizz[25][167] = 9'b111111111;
assign micromatrizz[25][168] = 9'b111111111;
assign micromatrizz[25][169] = 9'b111111111;
assign micromatrizz[25][170] = 9'b111111111;
assign micromatrizz[25][171] = 9'b111111111;
assign micromatrizz[25][172] = 9'b111111111;
assign micromatrizz[25][173] = 9'b111111111;
assign micromatrizz[25][174] = 9'b111111111;
assign micromatrizz[25][175] = 9'b111111111;
assign micromatrizz[25][176] = 9'b111111111;
assign micromatrizz[25][177] = 9'b111111111;
assign micromatrizz[25][178] = 9'b111111111;
assign micromatrizz[25][179] = 9'b111111111;
assign micromatrizz[25][180] = 9'b111111111;
assign micromatrizz[25][181] = 9'b111111111;
assign micromatrizz[25][182] = 9'b111111111;
assign micromatrizz[25][183] = 9'b111111111;
assign micromatrizz[25][184] = 9'b111111111;
assign micromatrizz[25][185] = 9'b111111111;
assign micromatrizz[25][186] = 9'b111111111;
assign micromatrizz[25][187] = 9'b111111111;
assign micromatrizz[25][188] = 9'b111111111;
assign micromatrizz[25][189] = 9'b111111111;
assign micromatrizz[25][190] = 9'b111111111;
assign micromatrizz[25][191] = 9'b111111111;
assign micromatrizz[25][192] = 9'b111111111;
assign micromatrizz[25][193] = 9'b111111111;
assign micromatrizz[25][194] = 9'b111111111;
assign micromatrizz[25][195] = 9'b111111111;
assign micromatrizz[25][196] = 9'b111111111;
assign micromatrizz[25][197] = 9'b111111111;
assign micromatrizz[25][198] = 9'b111111111;
assign micromatrizz[25][199] = 9'b111111111;
assign micromatrizz[25][200] = 9'b111111111;
assign micromatrizz[25][201] = 9'b111111111;
assign micromatrizz[25][202] = 9'b111111111;
assign micromatrizz[25][203] = 9'b111111111;
assign micromatrizz[25][204] = 9'b111111111;
assign micromatrizz[25][205] = 9'b111111111;
assign micromatrizz[25][206] = 9'b111111111;
assign micromatrizz[25][207] = 9'b111111111;
assign micromatrizz[25][208] = 9'b111111111;
assign micromatrizz[25][209] = 9'b111111111;
assign micromatrizz[25][210] = 9'b111111111;
assign micromatrizz[25][211] = 9'b111111111;
assign micromatrizz[25][212] = 9'b111111111;
assign micromatrizz[25][213] = 9'b111111111;
assign micromatrizz[25][214] = 9'b111111111;
assign micromatrizz[25][215] = 9'b111111111;
assign micromatrizz[25][216] = 9'b111111111;
assign micromatrizz[25][217] = 9'b111111111;
assign micromatrizz[25][218] = 9'b111111111;
assign micromatrizz[25][219] = 9'b111111111;
assign micromatrizz[25][220] = 9'b111111111;
assign micromatrizz[25][221] = 9'b111111111;
assign micromatrizz[25][222] = 9'b111111111;
assign micromatrizz[25][223] = 9'b111111111;
assign micromatrizz[25][224] = 9'b111111111;
assign micromatrizz[25][225] = 9'b111111111;
assign micromatrizz[25][226] = 9'b111111111;
assign micromatrizz[25][227] = 9'b111111111;
assign micromatrizz[25][228] = 9'b111111111;
assign micromatrizz[25][229] = 9'b111111111;
assign micromatrizz[25][230] = 9'b111111111;
assign micromatrizz[25][231] = 9'b111111111;
assign micromatrizz[25][232] = 9'b111111111;
assign micromatrizz[25][233] = 9'b111111111;
assign micromatrizz[25][234] = 9'b111111111;
assign micromatrizz[25][235] = 9'b111111111;
assign micromatrizz[25][236] = 9'b111111111;
assign micromatrizz[25][237] = 9'b111111111;
assign micromatrizz[25][238] = 9'b111111111;
assign micromatrizz[25][239] = 9'b111111111;
assign micromatrizz[25][240] = 9'b111111111;
assign micromatrizz[25][241] = 9'b111111111;
assign micromatrizz[25][242] = 9'b111111111;
assign micromatrizz[25][243] = 9'b111111111;
assign micromatrizz[25][244] = 9'b111111111;
assign micromatrizz[25][245] = 9'b111111111;
assign micromatrizz[25][246] = 9'b111111111;
assign micromatrizz[25][247] = 9'b111111111;
assign micromatrizz[25][248] = 9'b111111111;
assign micromatrizz[25][249] = 9'b111111111;
assign micromatrizz[25][250] = 9'b111111111;
assign micromatrizz[25][251] = 9'b111111111;
assign micromatrizz[25][252] = 9'b111111111;
assign micromatrizz[25][253] = 9'b111111111;
assign micromatrizz[25][254] = 9'b111111111;
assign micromatrizz[25][255] = 9'b111111111;
assign micromatrizz[25][256] = 9'b111111111;
assign micromatrizz[25][257] = 9'b111111111;
assign micromatrizz[25][258] = 9'b111111111;
assign micromatrizz[25][259] = 9'b111111111;
assign micromatrizz[25][260] = 9'b111111111;
assign micromatrizz[25][261] = 9'b111111111;
assign micromatrizz[25][262] = 9'b111111111;
assign micromatrizz[25][263] = 9'b111111111;
assign micromatrizz[25][264] = 9'b111111111;
assign micromatrizz[25][265] = 9'b111111111;
assign micromatrizz[25][266] = 9'b111111111;
assign micromatrizz[25][267] = 9'b111111111;
assign micromatrizz[25][268] = 9'b111111111;
assign micromatrizz[25][269] = 9'b111111111;
assign micromatrizz[25][270] = 9'b111110010;
assign micromatrizz[25][271] = 9'b111110010;
assign micromatrizz[25][272] = 9'b111110010;
assign micromatrizz[25][273] = 9'b111110010;
assign micromatrizz[25][274] = 9'b111110011;
assign micromatrizz[25][275] = 9'b111110011;
assign micromatrizz[25][276] = 9'b111110011;
assign micromatrizz[25][277] = 9'b111110011;
assign micromatrizz[25][278] = 9'b111110011;
assign micromatrizz[25][279] = 9'b111111111;
assign micromatrizz[25][280] = 9'b111111111;
assign micromatrizz[25][281] = 9'b111111111;
assign micromatrizz[25][282] = 9'b111111111;
assign micromatrizz[25][283] = 9'b111111111;
assign micromatrizz[25][284] = 9'b111111111;
assign micromatrizz[25][285] = 9'b111111111;
assign micromatrizz[25][286] = 9'b111111111;
assign micromatrizz[25][287] = 9'b111111111;
assign micromatrizz[25][288] = 9'b111111111;
assign micromatrizz[25][289] = 9'b111111111;
assign micromatrizz[25][290] = 9'b111111111;
assign micromatrizz[25][291] = 9'b111110010;
assign micromatrizz[25][292] = 9'b111110011;
assign micromatrizz[25][293] = 9'b111110011;
assign micromatrizz[25][294] = 9'b111110011;
assign micromatrizz[25][295] = 9'b111110011;
assign micromatrizz[25][296] = 9'b111110011;
assign micromatrizz[25][297] = 9'b111110111;
assign micromatrizz[25][298] = 9'b111111111;
assign micromatrizz[25][299] = 9'b111111111;
assign micromatrizz[25][300] = 9'b111111111;
assign micromatrizz[25][301] = 9'b111111111;
assign micromatrizz[25][302] = 9'b111111111;
assign micromatrizz[25][303] = 9'b111111111;
assign micromatrizz[25][304] = 9'b111110110;
assign micromatrizz[25][305] = 9'b111111111;
assign micromatrizz[25][306] = 9'b111111111;
assign micromatrizz[25][307] = 9'b111111111;
assign micromatrizz[25][308] = 9'b111110111;
assign micromatrizz[25][309] = 9'b111110010;
assign micromatrizz[25][310] = 9'b111110010;
assign micromatrizz[25][311] = 9'b111110010;
assign micromatrizz[25][312] = 9'b111110011;
assign micromatrizz[25][313] = 9'b111110010;
assign micromatrizz[25][314] = 9'b111110010;
assign micromatrizz[25][315] = 9'b111111111;
assign micromatrizz[25][316] = 9'b111111111;
assign micromatrizz[25][317] = 9'b111111111;
assign micromatrizz[25][318] = 9'b111111111;
assign micromatrizz[25][319] = 9'b111111111;
assign micromatrizz[25][320] = 9'b111111111;
assign micromatrizz[25][321] = 9'b111111111;
assign micromatrizz[25][322] = 9'b111111111;
assign micromatrizz[25][323] = 9'b111111111;
assign micromatrizz[25][324] = 9'b111111111;
assign micromatrizz[25][325] = 9'b111111111;
assign micromatrizz[25][326] = 9'b111111111;
assign micromatrizz[25][327] = 9'b111111111;
assign micromatrizz[25][328] = 9'b111111111;
assign micromatrizz[25][329] = 9'b111111111;
assign micromatrizz[25][330] = 9'b111111111;
assign micromatrizz[25][331] = 9'b111111111;
assign micromatrizz[25][332] = 9'b111111111;
assign micromatrizz[25][333] = 9'b111111111;
assign micromatrizz[25][334] = 9'b111111111;
assign micromatrizz[25][335] = 9'b111111111;
assign micromatrizz[25][336] = 9'b111111111;
assign micromatrizz[25][337] = 9'b111111111;
assign micromatrizz[25][338] = 9'b111111111;
assign micromatrizz[25][339] = 9'b111111111;
assign micromatrizz[25][340] = 9'b111111111;
assign micromatrizz[25][341] = 9'b111111111;
assign micromatrizz[25][342] = 9'b111111111;
assign micromatrizz[25][343] = 9'b111111111;
assign micromatrizz[25][344] = 9'b111111111;
assign micromatrizz[25][345] = 9'b111111111;
assign micromatrizz[25][346] = 9'b111111111;
assign micromatrizz[25][347] = 9'b111111111;
assign micromatrizz[25][348] = 9'b111111111;
assign micromatrizz[25][349] = 9'b111111111;
assign micromatrizz[25][350] = 9'b111111111;
assign micromatrizz[25][351] = 9'b111111111;
assign micromatrizz[25][352] = 9'b111111111;
assign micromatrizz[25][353] = 9'b111111111;
assign micromatrizz[25][354] = 9'b111111111;
assign micromatrizz[25][355] = 9'b111111111;
assign micromatrizz[25][356] = 9'b111111111;
assign micromatrizz[25][357] = 9'b111111111;
assign micromatrizz[25][358] = 9'b111111111;
assign micromatrizz[25][359] = 9'b111111111;
assign micromatrizz[25][360] = 9'b111111111;
assign micromatrizz[25][361] = 9'b111111111;
assign micromatrizz[25][362] = 9'b111111111;
assign micromatrizz[25][363] = 9'b111111111;
assign micromatrizz[25][364] = 9'b111111111;
assign micromatrizz[25][365] = 9'b111111111;
assign micromatrizz[25][366] = 9'b111111111;
assign micromatrizz[25][367] = 9'b111111111;
assign micromatrizz[25][368] = 9'b111111111;
assign micromatrizz[25][369] = 9'b111111111;
assign micromatrizz[25][370] = 9'b111111111;
assign micromatrizz[25][371] = 9'b111111111;
assign micromatrizz[25][372] = 9'b111111111;
assign micromatrizz[25][373] = 9'b111111111;
assign micromatrizz[25][374] = 9'b111111111;
assign micromatrizz[25][375] = 9'b111111111;
assign micromatrizz[25][376] = 9'b111111111;
assign micromatrizz[25][377] = 9'b111111111;
assign micromatrizz[25][378] = 9'b111111111;
assign micromatrizz[25][379] = 9'b111111111;
assign micromatrizz[25][380] = 9'b111111111;
assign micromatrizz[25][381] = 9'b111111111;
assign micromatrizz[25][382] = 9'b111111111;
assign micromatrizz[25][383] = 9'b111111111;
assign micromatrizz[25][384] = 9'b111111111;
assign micromatrizz[25][385] = 9'b111111111;
assign micromatrizz[25][386] = 9'b111111111;
assign micromatrizz[25][387] = 9'b111111111;
assign micromatrizz[25][388] = 9'b111111111;
assign micromatrizz[25][389] = 9'b111111111;
assign micromatrizz[25][390] = 9'b111111111;
assign micromatrizz[25][391] = 9'b111111111;
assign micromatrizz[25][392] = 9'b111111111;
assign micromatrizz[25][393] = 9'b111111111;
assign micromatrizz[25][394] = 9'b111111111;
assign micromatrizz[25][395] = 9'b111111111;
assign micromatrizz[25][396] = 9'b111111111;
assign micromatrizz[25][397] = 9'b111111111;
assign micromatrizz[25][398] = 9'b111111111;
assign micromatrizz[25][399] = 9'b111111111;
assign micromatrizz[25][400] = 9'b111111111;
assign micromatrizz[25][401] = 9'b111111111;
assign micromatrizz[25][402] = 9'b111111111;
assign micromatrizz[25][403] = 9'b111111111;
assign micromatrizz[25][404] = 9'b111111111;
assign micromatrizz[25][405] = 9'b111111111;
assign micromatrizz[25][406] = 9'b111111111;
assign micromatrizz[25][407] = 9'b111111111;
assign micromatrizz[25][408] = 9'b111111111;
assign micromatrizz[25][409] = 9'b111111111;
assign micromatrizz[25][410] = 9'b111111111;
assign micromatrizz[25][411] = 9'b111111111;
assign micromatrizz[25][412] = 9'b111111111;
assign micromatrizz[25][413] = 9'b111111111;
assign micromatrizz[25][414] = 9'b111111111;
assign micromatrizz[25][415] = 9'b111111111;
assign micromatrizz[25][416] = 9'b111111111;
assign micromatrizz[25][417] = 9'b111111111;
assign micromatrizz[25][418] = 9'b111111111;
assign micromatrizz[25][419] = 9'b111111111;
assign micromatrizz[25][420] = 9'b111111111;
assign micromatrizz[25][421] = 9'b111111111;
assign micromatrizz[25][422] = 9'b111111111;
assign micromatrizz[25][423] = 9'b111111111;
assign micromatrizz[25][424] = 9'b111111111;
assign micromatrizz[25][425] = 9'b111111111;
assign micromatrizz[25][426] = 9'b111111111;
assign micromatrizz[25][427] = 9'b111111111;
assign micromatrizz[25][428] = 9'b111111111;
assign micromatrizz[25][429] = 9'b111111111;
assign micromatrizz[25][430] = 9'b111111111;
assign micromatrizz[25][431] = 9'b111111111;
assign micromatrizz[25][432] = 9'b111111111;
assign micromatrizz[25][433] = 9'b111111111;
assign micromatrizz[25][434] = 9'b111111111;
assign micromatrizz[25][435] = 9'b111111111;
assign micromatrizz[25][436] = 9'b111111111;
assign micromatrizz[25][437] = 9'b111111111;
assign micromatrizz[25][438] = 9'b111111111;
assign micromatrizz[25][439] = 9'b111111111;
assign micromatrizz[25][440] = 9'b111111111;
assign micromatrizz[25][441] = 9'b111111111;
assign micromatrizz[25][442] = 9'b111111111;
assign micromatrizz[25][443] = 9'b111111111;
assign micromatrizz[25][444] = 9'b111111111;
assign micromatrizz[25][445] = 9'b111111111;
assign micromatrizz[25][446] = 9'b111111111;
assign micromatrizz[25][447] = 9'b111111111;
assign micromatrizz[25][448] = 9'b111111111;
assign micromatrizz[25][449] = 9'b111111111;
assign micromatrizz[25][450] = 9'b111111111;
assign micromatrizz[25][451] = 9'b111111111;
assign micromatrizz[25][452] = 9'b111111111;
assign micromatrizz[25][453] = 9'b111111111;
assign micromatrizz[25][454] = 9'b111111111;
assign micromatrizz[25][455] = 9'b111111111;
assign micromatrizz[25][456] = 9'b111111111;
assign micromatrizz[25][457] = 9'b111111111;
assign micromatrizz[25][458] = 9'b111111111;
assign micromatrizz[25][459] = 9'b111111111;
assign micromatrizz[25][460] = 9'b111111111;
assign micromatrizz[25][461] = 9'b111111111;
assign micromatrizz[25][462] = 9'b111111111;
assign micromatrizz[25][463] = 9'b111111111;
assign micromatrizz[25][464] = 9'b111111111;
assign micromatrizz[25][465] = 9'b111111111;
assign micromatrizz[25][466] = 9'b111111111;
assign micromatrizz[25][467] = 9'b111111111;
assign micromatrizz[25][468] = 9'b111111111;
assign micromatrizz[25][469] = 9'b111111111;
assign micromatrizz[25][470] = 9'b111111111;
assign micromatrizz[25][471] = 9'b111111111;
assign micromatrizz[25][472] = 9'b111111111;
assign micromatrizz[25][473] = 9'b111111111;
assign micromatrizz[25][474] = 9'b111111111;
assign micromatrizz[25][475] = 9'b111111111;
assign micromatrizz[25][476] = 9'b111111111;
assign micromatrizz[25][477] = 9'b111111111;
assign micromatrizz[25][478] = 9'b111111111;
assign micromatrizz[25][479] = 9'b111111111;
assign micromatrizz[25][480] = 9'b111111111;
assign micromatrizz[25][481] = 9'b111111111;
assign micromatrizz[25][482] = 9'b111111111;
assign micromatrizz[25][483] = 9'b111111111;
assign micromatrizz[25][484] = 9'b111111111;
assign micromatrizz[25][485] = 9'b111111111;
assign micromatrizz[25][486] = 9'b111111111;
assign micromatrizz[25][487] = 9'b111111111;
assign micromatrizz[25][488] = 9'b111111111;
assign micromatrizz[25][489] = 9'b111111111;
assign micromatrizz[25][490] = 9'b111111111;
assign micromatrizz[25][491] = 9'b111111111;
assign micromatrizz[25][492] = 9'b111111111;
assign micromatrizz[25][493] = 9'b111111111;
assign micromatrizz[25][494] = 9'b111111111;
assign micromatrizz[25][495] = 9'b111111111;
assign micromatrizz[25][496] = 9'b111111111;
assign micromatrizz[25][497] = 9'b111111111;
assign micromatrizz[25][498] = 9'b111111111;
assign micromatrizz[25][499] = 9'b111111111;
assign micromatrizz[25][500] = 9'b111111111;
assign micromatrizz[25][501] = 9'b111111111;
assign micromatrizz[25][502] = 9'b111111111;
assign micromatrizz[25][503] = 9'b111111111;
assign micromatrizz[25][504] = 9'b111111111;
assign micromatrizz[25][505] = 9'b111111111;
assign micromatrizz[25][506] = 9'b111111111;
assign micromatrizz[25][507] = 9'b111111111;
assign micromatrizz[25][508] = 9'b111111111;
assign micromatrizz[25][509] = 9'b111111111;
assign micromatrizz[25][510] = 9'b111111111;
assign micromatrizz[25][511] = 9'b111111111;
assign micromatrizz[25][512] = 9'b111111111;
assign micromatrizz[25][513] = 9'b111111111;
assign micromatrizz[25][514] = 9'b111111111;
assign micromatrizz[25][515] = 9'b111111111;
assign micromatrizz[25][516] = 9'b111111111;
assign micromatrizz[25][517] = 9'b111111111;
assign micromatrizz[25][518] = 9'b111111111;
assign micromatrizz[25][519] = 9'b111111111;
assign micromatrizz[25][520] = 9'b111111111;
assign micromatrizz[25][521] = 9'b111111111;
assign micromatrizz[25][522] = 9'b111111111;
assign micromatrizz[25][523] = 9'b111111111;
assign micromatrizz[25][524] = 9'b111111111;
assign micromatrizz[25][525] = 9'b111111111;
assign micromatrizz[25][526] = 9'b111111111;
assign micromatrizz[25][527] = 9'b111111111;
assign micromatrizz[25][528] = 9'b111111111;
assign micromatrizz[25][529] = 9'b111111111;
assign micromatrizz[25][530] = 9'b111111111;
assign micromatrizz[25][531] = 9'b111111111;
assign micromatrizz[25][532] = 9'b111111111;
assign micromatrizz[25][533] = 9'b111111111;
assign micromatrizz[25][534] = 9'b111111111;
assign micromatrizz[25][535] = 9'b111111111;
assign micromatrizz[25][536] = 9'b111111111;
assign micromatrizz[25][537] = 9'b111111111;
assign micromatrizz[25][538] = 9'b111111111;
assign micromatrizz[25][539] = 9'b111111111;
assign micromatrizz[25][540] = 9'b111111111;
assign micromatrizz[25][541] = 9'b111111111;
assign micromatrizz[25][542] = 9'b111111111;
assign micromatrizz[25][543] = 9'b111111111;
assign micromatrizz[25][544] = 9'b111111111;
assign micromatrizz[25][545] = 9'b111111111;
assign micromatrizz[25][546] = 9'b111111111;
assign micromatrizz[25][547] = 9'b111111111;
assign micromatrizz[25][548] = 9'b111111111;
assign micromatrizz[25][549] = 9'b111111111;
assign micromatrizz[25][550] = 9'b111111111;
assign micromatrizz[25][551] = 9'b111111111;
assign micromatrizz[25][552] = 9'b111111111;
assign micromatrizz[25][553] = 9'b111111111;
assign micromatrizz[25][554] = 9'b111111111;
assign micromatrizz[25][555] = 9'b111111111;
assign micromatrizz[25][556] = 9'b111111111;
assign micromatrizz[25][557] = 9'b111111111;
assign micromatrizz[25][558] = 9'b111111111;
assign micromatrizz[25][559] = 9'b111111111;
assign micromatrizz[25][560] = 9'b111111111;
assign micromatrizz[25][561] = 9'b111111111;
assign micromatrizz[25][562] = 9'b111111111;
assign micromatrizz[25][563] = 9'b111111111;
assign micromatrizz[25][564] = 9'b111111111;
assign micromatrizz[25][565] = 9'b111111111;
assign micromatrizz[25][566] = 9'b111111111;
assign micromatrizz[25][567] = 9'b111111111;
assign micromatrizz[25][568] = 9'b111111111;
assign micromatrizz[25][569] = 9'b111111111;
assign micromatrizz[25][570] = 9'b111111111;
assign micromatrizz[25][571] = 9'b111111111;
assign micromatrizz[25][572] = 9'b111111111;
assign micromatrizz[25][573] = 9'b111111111;
assign micromatrizz[25][574] = 9'b111111111;
assign micromatrizz[25][575] = 9'b111111111;
assign micromatrizz[25][576] = 9'b111111111;
assign micromatrizz[25][577] = 9'b111111111;
assign micromatrizz[25][578] = 9'b111111111;
assign micromatrizz[25][579] = 9'b111111111;
assign micromatrizz[25][580] = 9'b111111111;
assign micromatrizz[25][581] = 9'b111111111;
assign micromatrizz[25][582] = 9'b111111111;
assign micromatrizz[25][583] = 9'b111111111;
assign micromatrizz[25][584] = 9'b111111111;
assign micromatrizz[25][585] = 9'b111111111;
assign micromatrizz[25][586] = 9'b111111111;
assign micromatrizz[25][587] = 9'b111111111;
assign micromatrizz[25][588] = 9'b111111111;
assign micromatrizz[25][589] = 9'b111111111;
assign micromatrizz[25][590] = 9'b111111111;
assign micromatrizz[25][591] = 9'b111111111;
assign micromatrizz[25][592] = 9'b111111111;
assign micromatrizz[25][593] = 9'b111111111;
assign micromatrizz[25][594] = 9'b111111111;
assign micromatrizz[25][595] = 9'b111111111;
assign micromatrizz[25][596] = 9'b111111111;
assign micromatrizz[25][597] = 9'b111111111;
assign micromatrizz[25][598] = 9'b111111111;
assign micromatrizz[25][599] = 9'b111111111;
assign micromatrizz[25][600] = 9'b111111111;
assign micromatrizz[25][601] = 9'b111111111;
assign micromatrizz[25][602] = 9'b111111111;
assign micromatrizz[25][603] = 9'b111111111;
assign micromatrizz[25][604] = 9'b111111111;
assign micromatrizz[25][605] = 9'b111111111;
assign micromatrizz[25][606] = 9'b111111111;
assign micromatrizz[25][607] = 9'b111111111;
assign micromatrizz[25][608] = 9'b111111111;
assign micromatrizz[25][609] = 9'b111111111;
assign micromatrizz[25][610] = 9'b111111111;
assign micromatrizz[25][611] = 9'b111111111;
assign micromatrizz[25][612] = 9'b111111111;
assign micromatrizz[25][613] = 9'b111111111;
assign micromatrizz[25][614] = 9'b111111111;
assign micromatrizz[25][615] = 9'b111111111;
assign micromatrizz[25][616] = 9'b111111111;
assign micromatrizz[25][617] = 9'b111111111;
assign micromatrizz[25][618] = 9'b111111111;
assign micromatrizz[25][619] = 9'b111111111;
assign micromatrizz[25][620] = 9'b111111111;
assign micromatrizz[25][621] = 9'b111111111;
assign micromatrizz[25][622] = 9'b111111111;
assign micromatrizz[25][623] = 9'b111111111;
assign micromatrizz[25][624] = 9'b111111111;
assign micromatrizz[25][625] = 9'b111111111;
assign micromatrizz[25][626] = 9'b111111111;
assign micromatrizz[25][627] = 9'b111111111;
assign micromatrizz[25][628] = 9'b111111111;
assign micromatrizz[25][629] = 9'b111111111;
assign micromatrizz[25][630] = 9'b111111111;
assign micromatrizz[25][631] = 9'b111111111;
assign micromatrizz[25][632] = 9'b111111111;
assign micromatrizz[25][633] = 9'b111111111;
assign micromatrizz[25][634] = 9'b111111111;
assign micromatrizz[25][635] = 9'b111111111;
assign micromatrizz[25][636] = 9'b111111111;
assign micromatrizz[25][637] = 9'b111111111;
assign micromatrizz[25][638] = 9'b111111111;
assign micromatrizz[25][639] = 9'b111111111;
assign micromatrizz[26][0] = 9'b111111111;
assign micromatrizz[26][1] = 9'b111111111;
assign micromatrizz[26][2] = 9'b111111111;
assign micromatrizz[26][3] = 9'b111111111;
assign micromatrizz[26][4] = 9'b111111111;
assign micromatrizz[26][5] = 9'b111111111;
assign micromatrizz[26][6] = 9'b111111111;
assign micromatrizz[26][7] = 9'b111111111;
assign micromatrizz[26][8] = 9'b111111111;
assign micromatrizz[26][9] = 9'b111111111;
assign micromatrizz[26][10] = 9'b111111111;
assign micromatrizz[26][11] = 9'b111111111;
assign micromatrizz[26][12] = 9'b111111111;
assign micromatrizz[26][13] = 9'b111111111;
assign micromatrizz[26][14] = 9'b111111111;
assign micromatrizz[26][15] = 9'b111111111;
assign micromatrizz[26][16] = 9'b111111111;
assign micromatrizz[26][17] = 9'b111111111;
assign micromatrizz[26][18] = 9'b111111111;
assign micromatrizz[26][19] = 9'b111111111;
assign micromatrizz[26][20] = 9'b111111111;
assign micromatrizz[26][21] = 9'b111111111;
assign micromatrizz[26][22] = 9'b111111111;
assign micromatrizz[26][23] = 9'b111111111;
assign micromatrizz[26][24] = 9'b111111111;
assign micromatrizz[26][25] = 9'b111111111;
assign micromatrizz[26][26] = 9'b111111111;
assign micromatrizz[26][27] = 9'b111111111;
assign micromatrizz[26][28] = 9'b111111111;
assign micromatrizz[26][29] = 9'b111111111;
assign micromatrizz[26][30] = 9'b111111111;
assign micromatrizz[26][31] = 9'b111111111;
assign micromatrizz[26][32] = 9'b111111111;
assign micromatrizz[26][33] = 9'b111111111;
assign micromatrizz[26][34] = 9'b111111111;
assign micromatrizz[26][35] = 9'b111111111;
assign micromatrizz[26][36] = 9'b111111111;
assign micromatrizz[26][37] = 9'b111111111;
assign micromatrizz[26][38] = 9'b111111111;
assign micromatrizz[26][39] = 9'b111111111;
assign micromatrizz[26][40] = 9'b111111111;
assign micromatrizz[26][41] = 9'b111111111;
assign micromatrizz[26][42] = 9'b111111111;
assign micromatrizz[26][43] = 9'b111111111;
assign micromatrizz[26][44] = 9'b111111111;
assign micromatrizz[26][45] = 9'b111111111;
assign micromatrizz[26][46] = 9'b111111111;
assign micromatrizz[26][47] = 9'b111111111;
assign micromatrizz[26][48] = 9'b111111111;
assign micromatrizz[26][49] = 9'b111111111;
assign micromatrizz[26][50] = 9'b111111111;
assign micromatrizz[26][51] = 9'b111111111;
assign micromatrizz[26][52] = 9'b111111111;
assign micromatrizz[26][53] = 9'b111111111;
assign micromatrizz[26][54] = 9'b111111111;
assign micromatrizz[26][55] = 9'b111111111;
assign micromatrizz[26][56] = 9'b111111111;
assign micromatrizz[26][57] = 9'b111111111;
assign micromatrizz[26][58] = 9'b111111111;
assign micromatrizz[26][59] = 9'b111111111;
assign micromatrizz[26][60] = 9'b111111111;
assign micromatrizz[26][61] = 9'b111111111;
assign micromatrizz[26][62] = 9'b111111111;
assign micromatrizz[26][63] = 9'b111111111;
assign micromatrizz[26][64] = 9'b111111111;
assign micromatrizz[26][65] = 9'b111111111;
assign micromatrizz[26][66] = 9'b111111111;
assign micromatrizz[26][67] = 9'b111111111;
assign micromatrizz[26][68] = 9'b111111111;
assign micromatrizz[26][69] = 9'b111111111;
assign micromatrizz[26][70] = 9'b111111111;
assign micromatrizz[26][71] = 9'b111111111;
assign micromatrizz[26][72] = 9'b111111111;
assign micromatrizz[26][73] = 9'b111111111;
assign micromatrizz[26][74] = 9'b111111111;
assign micromatrizz[26][75] = 9'b111111111;
assign micromatrizz[26][76] = 9'b111111111;
assign micromatrizz[26][77] = 9'b111111111;
assign micromatrizz[26][78] = 9'b111111111;
assign micromatrizz[26][79] = 9'b111111111;
assign micromatrizz[26][80] = 9'b111111111;
assign micromatrizz[26][81] = 9'b111111111;
assign micromatrizz[26][82] = 9'b111111111;
assign micromatrizz[26][83] = 9'b111111111;
assign micromatrizz[26][84] = 9'b111111111;
assign micromatrizz[26][85] = 9'b111111111;
assign micromatrizz[26][86] = 9'b111111111;
assign micromatrizz[26][87] = 9'b111111111;
assign micromatrizz[26][88] = 9'b111111111;
assign micromatrizz[26][89] = 9'b111111111;
assign micromatrizz[26][90] = 9'b111111111;
assign micromatrizz[26][91] = 9'b111111111;
assign micromatrizz[26][92] = 9'b111111111;
assign micromatrizz[26][93] = 9'b111111111;
assign micromatrizz[26][94] = 9'b111111111;
assign micromatrizz[26][95] = 9'b111111111;
assign micromatrizz[26][96] = 9'b111111111;
assign micromatrizz[26][97] = 9'b111111111;
assign micromatrizz[26][98] = 9'b111111111;
assign micromatrizz[26][99] = 9'b111111111;
assign micromatrizz[26][100] = 9'b111111111;
assign micromatrizz[26][101] = 9'b111111111;
assign micromatrizz[26][102] = 9'b111111111;
assign micromatrizz[26][103] = 9'b111111111;
assign micromatrizz[26][104] = 9'b111111111;
assign micromatrizz[26][105] = 9'b111111111;
assign micromatrizz[26][106] = 9'b111111111;
assign micromatrizz[26][107] = 9'b111111111;
assign micromatrizz[26][108] = 9'b111111111;
assign micromatrizz[26][109] = 9'b111111111;
assign micromatrizz[26][110] = 9'b111111111;
assign micromatrizz[26][111] = 9'b111111111;
assign micromatrizz[26][112] = 9'b111111111;
assign micromatrizz[26][113] = 9'b111111111;
assign micromatrizz[26][114] = 9'b111111111;
assign micromatrizz[26][115] = 9'b111111111;
assign micromatrizz[26][116] = 9'b111111111;
assign micromatrizz[26][117] = 9'b111111111;
assign micromatrizz[26][118] = 9'b111111111;
assign micromatrizz[26][119] = 9'b111111111;
assign micromatrizz[26][120] = 9'b111111111;
assign micromatrizz[26][121] = 9'b111111111;
assign micromatrizz[26][122] = 9'b111111111;
assign micromatrizz[26][123] = 9'b111111111;
assign micromatrizz[26][124] = 9'b111111111;
assign micromatrizz[26][125] = 9'b111111111;
assign micromatrizz[26][126] = 9'b111111111;
assign micromatrizz[26][127] = 9'b111111111;
assign micromatrizz[26][128] = 9'b111111111;
assign micromatrizz[26][129] = 9'b111111111;
assign micromatrizz[26][130] = 9'b111111111;
assign micromatrizz[26][131] = 9'b111111111;
assign micromatrizz[26][132] = 9'b111111111;
assign micromatrizz[26][133] = 9'b111111111;
assign micromatrizz[26][134] = 9'b111111111;
assign micromatrizz[26][135] = 9'b111111111;
assign micromatrizz[26][136] = 9'b111111111;
assign micromatrizz[26][137] = 9'b111111111;
assign micromatrizz[26][138] = 9'b111111111;
assign micromatrizz[26][139] = 9'b111111111;
assign micromatrizz[26][140] = 9'b111111111;
assign micromatrizz[26][141] = 9'b111111111;
assign micromatrizz[26][142] = 9'b111111111;
assign micromatrizz[26][143] = 9'b111111111;
assign micromatrizz[26][144] = 9'b111111111;
assign micromatrizz[26][145] = 9'b111111111;
assign micromatrizz[26][146] = 9'b111111111;
assign micromatrizz[26][147] = 9'b111111111;
assign micromatrizz[26][148] = 9'b111111111;
assign micromatrizz[26][149] = 9'b111111111;
assign micromatrizz[26][150] = 9'b111111111;
assign micromatrizz[26][151] = 9'b111111111;
assign micromatrizz[26][152] = 9'b111111111;
assign micromatrizz[26][153] = 9'b111111111;
assign micromatrizz[26][154] = 9'b111111111;
assign micromatrizz[26][155] = 9'b111111111;
assign micromatrizz[26][156] = 9'b111111111;
assign micromatrizz[26][157] = 9'b111111111;
assign micromatrizz[26][158] = 9'b111111111;
assign micromatrizz[26][159] = 9'b111111111;
assign micromatrizz[26][160] = 9'b111111111;
assign micromatrizz[26][161] = 9'b111111111;
assign micromatrizz[26][162] = 9'b111111111;
assign micromatrizz[26][163] = 9'b111111111;
assign micromatrizz[26][164] = 9'b111111111;
assign micromatrizz[26][165] = 9'b111111111;
assign micromatrizz[26][166] = 9'b111111111;
assign micromatrizz[26][167] = 9'b111111111;
assign micromatrizz[26][168] = 9'b111111111;
assign micromatrizz[26][169] = 9'b111111111;
assign micromatrizz[26][170] = 9'b111111111;
assign micromatrizz[26][171] = 9'b111111111;
assign micromatrizz[26][172] = 9'b111111111;
assign micromatrizz[26][173] = 9'b111111111;
assign micromatrizz[26][174] = 9'b111111111;
assign micromatrizz[26][175] = 9'b111111111;
assign micromatrizz[26][176] = 9'b111111111;
assign micromatrizz[26][177] = 9'b111111111;
assign micromatrizz[26][178] = 9'b111111111;
assign micromatrizz[26][179] = 9'b111111111;
assign micromatrizz[26][180] = 9'b111111111;
assign micromatrizz[26][181] = 9'b111111111;
assign micromatrizz[26][182] = 9'b111111111;
assign micromatrizz[26][183] = 9'b111111111;
assign micromatrizz[26][184] = 9'b111111111;
assign micromatrizz[26][185] = 9'b111111111;
assign micromatrizz[26][186] = 9'b111111111;
assign micromatrizz[26][187] = 9'b111111111;
assign micromatrizz[26][188] = 9'b111111111;
assign micromatrizz[26][189] = 9'b111111111;
assign micromatrizz[26][190] = 9'b111111111;
assign micromatrizz[26][191] = 9'b111111111;
assign micromatrizz[26][192] = 9'b111111111;
assign micromatrizz[26][193] = 9'b111111111;
assign micromatrizz[26][194] = 9'b111111111;
assign micromatrizz[26][195] = 9'b111111111;
assign micromatrizz[26][196] = 9'b111111111;
assign micromatrizz[26][197] = 9'b111111111;
assign micromatrizz[26][198] = 9'b111111111;
assign micromatrizz[26][199] = 9'b111111111;
assign micromatrizz[26][200] = 9'b111111111;
assign micromatrizz[26][201] = 9'b111111111;
assign micromatrizz[26][202] = 9'b111111111;
assign micromatrizz[26][203] = 9'b111111111;
assign micromatrizz[26][204] = 9'b111111111;
assign micromatrizz[26][205] = 9'b111111111;
assign micromatrizz[26][206] = 9'b111111111;
assign micromatrizz[26][207] = 9'b111111111;
assign micromatrizz[26][208] = 9'b111111111;
assign micromatrizz[26][209] = 9'b111111111;
assign micromatrizz[26][210] = 9'b111111111;
assign micromatrizz[26][211] = 9'b111111111;
assign micromatrizz[26][212] = 9'b111111111;
assign micromatrizz[26][213] = 9'b111111111;
assign micromatrizz[26][214] = 9'b111111111;
assign micromatrizz[26][215] = 9'b111111111;
assign micromatrizz[26][216] = 9'b111111111;
assign micromatrizz[26][217] = 9'b111111111;
assign micromatrizz[26][218] = 9'b111111111;
assign micromatrizz[26][219] = 9'b111111111;
assign micromatrizz[26][220] = 9'b111111111;
assign micromatrizz[26][221] = 9'b111111111;
assign micromatrizz[26][222] = 9'b111111111;
assign micromatrizz[26][223] = 9'b111111111;
assign micromatrizz[26][224] = 9'b111111111;
assign micromatrizz[26][225] = 9'b111111111;
assign micromatrizz[26][226] = 9'b111111111;
assign micromatrizz[26][227] = 9'b111111111;
assign micromatrizz[26][228] = 9'b111111111;
assign micromatrizz[26][229] = 9'b111111111;
assign micromatrizz[26][230] = 9'b111111111;
assign micromatrizz[26][231] = 9'b111111111;
assign micromatrizz[26][232] = 9'b111111111;
assign micromatrizz[26][233] = 9'b111111111;
assign micromatrizz[26][234] = 9'b111111111;
assign micromatrizz[26][235] = 9'b111111111;
assign micromatrizz[26][236] = 9'b111111111;
assign micromatrizz[26][237] = 9'b111111111;
assign micromatrizz[26][238] = 9'b111111111;
assign micromatrizz[26][239] = 9'b111111111;
assign micromatrizz[26][240] = 9'b111111111;
assign micromatrizz[26][241] = 9'b111111111;
assign micromatrizz[26][242] = 9'b111111111;
assign micromatrizz[26][243] = 9'b111111111;
assign micromatrizz[26][244] = 9'b111111111;
assign micromatrizz[26][245] = 9'b111111111;
assign micromatrizz[26][246] = 9'b111111111;
assign micromatrizz[26][247] = 9'b111111111;
assign micromatrizz[26][248] = 9'b111111111;
assign micromatrizz[26][249] = 9'b111111111;
assign micromatrizz[26][250] = 9'b111111111;
assign micromatrizz[26][251] = 9'b111111111;
assign micromatrizz[26][252] = 9'b111111111;
assign micromatrizz[26][253] = 9'b111111111;
assign micromatrizz[26][254] = 9'b111111111;
assign micromatrizz[26][255] = 9'b111111111;
assign micromatrizz[26][256] = 9'b111111111;
assign micromatrizz[26][257] = 9'b111111111;
assign micromatrizz[26][258] = 9'b111111111;
assign micromatrizz[26][259] = 9'b111111111;
assign micromatrizz[26][260] = 9'b111111111;
assign micromatrizz[26][261] = 9'b111111111;
assign micromatrizz[26][262] = 9'b111111111;
assign micromatrizz[26][263] = 9'b111111111;
assign micromatrizz[26][264] = 9'b111111111;
assign micromatrizz[26][265] = 9'b111111111;
assign micromatrizz[26][266] = 9'b111111111;
assign micromatrizz[26][267] = 9'b111111111;
assign micromatrizz[26][268] = 9'b111111111;
assign micromatrizz[26][269] = 9'b111111111;
assign micromatrizz[26][270] = 9'b111110010;
assign micromatrizz[26][271] = 9'b111110010;
assign micromatrizz[26][272] = 9'b111110010;
assign micromatrizz[26][273] = 9'b111110010;
assign micromatrizz[26][274] = 9'b111110011;
assign micromatrizz[26][275] = 9'b111110011;
assign micromatrizz[26][276] = 9'b111110011;
assign micromatrizz[26][277] = 9'b111110011;
assign micromatrizz[26][278] = 9'b111110011;
assign micromatrizz[26][279] = 9'b111111111;
assign micromatrizz[26][280] = 9'b111111111;
assign micromatrizz[26][281] = 9'b111111111;
assign micromatrizz[26][282] = 9'b111111111;
assign micromatrizz[26][283] = 9'b111111111;
assign micromatrizz[26][284] = 9'b111111111;
assign micromatrizz[26][285] = 9'b111111111;
assign micromatrizz[26][286] = 9'b111111111;
assign micromatrizz[26][287] = 9'b111111111;
assign micromatrizz[26][288] = 9'b111111111;
assign micromatrizz[26][289] = 9'b111111111;
assign micromatrizz[26][290] = 9'b111110111;
assign micromatrizz[26][291] = 9'b111110010;
assign micromatrizz[26][292] = 9'b111110011;
assign micromatrizz[26][293] = 9'b111110010;
assign micromatrizz[26][294] = 9'b111110011;
assign micromatrizz[26][295] = 9'b111110011;
assign micromatrizz[26][296] = 9'b111110011;
assign micromatrizz[26][297] = 9'b111110111;
assign micromatrizz[26][298] = 9'b111111111;
assign micromatrizz[26][299] = 9'b111111111;
assign micromatrizz[26][300] = 9'b111111111;
assign micromatrizz[26][301] = 9'b111111111;
assign micromatrizz[26][302] = 9'b111111111;
assign micromatrizz[26][303] = 9'b111111111;
assign micromatrizz[26][304] = 9'b111110111;
assign micromatrizz[26][305] = 9'b111110111;
assign micromatrizz[26][306] = 9'b111111111;
assign micromatrizz[26][307] = 9'b111111111;
assign micromatrizz[26][308] = 9'b111110010;
assign micromatrizz[26][309] = 9'b111110010;
assign micromatrizz[26][310] = 9'b111110010;
assign micromatrizz[26][311] = 9'b111110010;
assign micromatrizz[26][312] = 9'b111110011;
assign micromatrizz[26][313] = 9'b111110010;
assign micromatrizz[26][314] = 9'b111110011;
assign micromatrizz[26][315] = 9'b111110011;
assign micromatrizz[26][316] = 9'b111111111;
assign micromatrizz[26][317] = 9'b111111111;
assign micromatrizz[26][318] = 9'b111111111;
assign micromatrizz[26][319] = 9'b111111111;
assign micromatrizz[26][320] = 9'b111111111;
assign micromatrizz[26][321] = 9'b111111111;
assign micromatrizz[26][322] = 9'b111111111;
assign micromatrizz[26][323] = 9'b111111111;
assign micromatrizz[26][324] = 9'b111111111;
assign micromatrizz[26][325] = 9'b111111111;
assign micromatrizz[26][326] = 9'b111111111;
assign micromatrizz[26][327] = 9'b111111111;
assign micromatrizz[26][328] = 9'b111111111;
assign micromatrizz[26][329] = 9'b111111111;
assign micromatrizz[26][330] = 9'b111111111;
assign micromatrizz[26][331] = 9'b111111111;
assign micromatrizz[26][332] = 9'b111111111;
assign micromatrizz[26][333] = 9'b111111111;
assign micromatrizz[26][334] = 9'b111111111;
assign micromatrizz[26][335] = 9'b111111111;
assign micromatrizz[26][336] = 9'b111111111;
assign micromatrizz[26][337] = 9'b111111111;
assign micromatrizz[26][338] = 9'b111111111;
assign micromatrizz[26][339] = 9'b111111111;
assign micromatrizz[26][340] = 9'b111111111;
assign micromatrizz[26][341] = 9'b111111111;
assign micromatrizz[26][342] = 9'b111111111;
assign micromatrizz[26][343] = 9'b111111111;
assign micromatrizz[26][344] = 9'b111111111;
assign micromatrizz[26][345] = 9'b111111111;
assign micromatrizz[26][346] = 9'b111111111;
assign micromatrizz[26][347] = 9'b111111111;
assign micromatrizz[26][348] = 9'b111111111;
assign micromatrizz[26][349] = 9'b111111111;
assign micromatrizz[26][350] = 9'b111111111;
assign micromatrizz[26][351] = 9'b111111111;
assign micromatrizz[26][352] = 9'b111111111;
assign micromatrizz[26][353] = 9'b111111111;
assign micromatrizz[26][354] = 9'b111111111;
assign micromatrizz[26][355] = 9'b111111111;
assign micromatrizz[26][356] = 9'b111111111;
assign micromatrizz[26][357] = 9'b111111111;
assign micromatrizz[26][358] = 9'b111111111;
assign micromatrizz[26][359] = 9'b111111111;
assign micromatrizz[26][360] = 9'b111111111;
assign micromatrizz[26][361] = 9'b111111111;
assign micromatrizz[26][362] = 9'b111111111;
assign micromatrizz[26][363] = 9'b111111111;
assign micromatrizz[26][364] = 9'b111111111;
assign micromatrizz[26][365] = 9'b111111111;
assign micromatrizz[26][366] = 9'b111111111;
assign micromatrizz[26][367] = 9'b111111111;
assign micromatrizz[26][368] = 9'b111111111;
assign micromatrizz[26][369] = 9'b111111111;
assign micromatrizz[26][370] = 9'b111111111;
assign micromatrizz[26][371] = 9'b111111111;
assign micromatrizz[26][372] = 9'b111111111;
assign micromatrizz[26][373] = 9'b111111111;
assign micromatrizz[26][374] = 9'b111111111;
assign micromatrizz[26][375] = 9'b111111111;
assign micromatrizz[26][376] = 9'b111111111;
assign micromatrizz[26][377] = 9'b111111111;
assign micromatrizz[26][378] = 9'b111111111;
assign micromatrizz[26][379] = 9'b111111111;
assign micromatrizz[26][380] = 9'b111111111;
assign micromatrizz[26][381] = 9'b111111111;
assign micromatrizz[26][382] = 9'b111111111;
assign micromatrizz[26][383] = 9'b111111111;
assign micromatrizz[26][384] = 9'b111111111;
assign micromatrizz[26][385] = 9'b111111111;
assign micromatrizz[26][386] = 9'b111111111;
assign micromatrizz[26][387] = 9'b111111111;
assign micromatrizz[26][388] = 9'b111111111;
assign micromatrizz[26][389] = 9'b111111111;
assign micromatrizz[26][390] = 9'b111111111;
assign micromatrizz[26][391] = 9'b111111111;
assign micromatrizz[26][392] = 9'b111111111;
assign micromatrizz[26][393] = 9'b111111111;
assign micromatrizz[26][394] = 9'b111111111;
assign micromatrizz[26][395] = 9'b111111111;
assign micromatrizz[26][396] = 9'b111111111;
assign micromatrizz[26][397] = 9'b111111111;
assign micromatrizz[26][398] = 9'b111111111;
assign micromatrizz[26][399] = 9'b111111111;
assign micromatrizz[26][400] = 9'b111111111;
assign micromatrizz[26][401] = 9'b111111111;
assign micromatrizz[26][402] = 9'b111111111;
assign micromatrizz[26][403] = 9'b111111111;
assign micromatrizz[26][404] = 9'b111111111;
assign micromatrizz[26][405] = 9'b111111111;
assign micromatrizz[26][406] = 9'b111111111;
assign micromatrizz[26][407] = 9'b111111111;
assign micromatrizz[26][408] = 9'b111111111;
assign micromatrizz[26][409] = 9'b111111111;
assign micromatrizz[26][410] = 9'b111111111;
assign micromatrizz[26][411] = 9'b111111111;
assign micromatrizz[26][412] = 9'b111111111;
assign micromatrizz[26][413] = 9'b111111111;
assign micromatrizz[26][414] = 9'b111111111;
assign micromatrizz[26][415] = 9'b111111111;
assign micromatrizz[26][416] = 9'b111111111;
assign micromatrizz[26][417] = 9'b111111111;
assign micromatrizz[26][418] = 9'b111111111;
assign micromatrizz[26][419] = 9'b111111111;
assign micromatrizz[26][420] = 9'b111111111;
assign micromatrizz[26][421] = 9'b111111111;
assign micromatrizz[26][422] = 9'b111111111;
assign micromatrizz[26][423] = 9'b111111111;
assign micromatrizz[26][424] = 9'b111111111;
assign micromatrizz[26][425] = 9'b111111111;
assign micromatrizz[26][426] = 9'b111111111;
assign micromatrizz[26][427] = 9'b111111111;
assign micromatrizz[26][428] = 9'b111111111;
assign micromatrizz[26][429] = 9'b111111111;
assign micromatrizz[26][430] = 9'b111111111;
assign micromatrizz[26][431] = 9'b111111111;
assign micromatrizz[26][432] = 9'b111111111;
assign micromatrizz[26][433] = 9'b111111111;
assign micromatrizz[26][434] = 9'b111111111;
assign micromatrizz[26][435] = 9'b111111111;
assign micromatrizz[26][436] = 9'b111111111;
assign micromatrizz[26][437] = 9'b111111111;
assign micromatrizz[26][438] = 9'b111111111;
assign micromatrizz[26][439] = 9'b111111111;
assign micromatrizz[26][440] = 9'b111111111;
assign micromatrizz[26][441] = 9'b111111111;
assign micromatrizz[26][442] = 9'b111111111;
assign micromatrizz[26][443] = 9'b111111111;
assign micromatrizz[26][444] = 9'b111111111;
assign micromatrizz[26][445] = 9'b111111111;
assign micromatrizz[26][446] = 9'b111111111;
assign micromatrizz[26][447] = 9'b111111111;
assign micromatrizz[26][448] = 9'b111111111;
assign micromatrizz[26][449] = 9'b111111111;
assign micromatrizz[26][450] = 9'b111111111;
assign micromatrizz[26][451] = 9'b111111111;
assign micromatrizz[26][452] = 9'b111111111;
assign micromatrizz[26][453] = 9'b111111111;
assign micromatrizz[26][454] = 9'b111111111;
assign micromatrizz[26][455] = 9'b111111111;
assign micromatrizz[26][456] = 9'b111111111;
assign micromatrizz[26][457] = 9'b111111111;
assign micromatrizz[26][458] = 9'b111111111;
assign micromatrizz[26][459] = 9'b111111111;
assign micromatrizz[26][460] = 9'b111111111;
assign micromatrizz[26][461] = 9'b111111111;
assign micromatrizz[26][462] = 9'b111111111;
assign micromatrizz[26][463] = 9'b111111111;
assign micromatrizz[26][464] = 9'b111111111;
assign micromatrizz[26][465] = 9'b111111111;
assign micromatrizz[26][466] = 9'b111111111;
assign micromatrizz[26][467] = 9'b111111111;
assign micromatrizz[26][468] = 9'b111111111;
assign micromatrizz[26][469] = 9'b111111111;
assign micromatrizz[26][470] = 9'b111111111;
assign micromatrizz[26][471] = 9'b111111111;
assign micromatrizz[26][472] = 9'b111111111;
assign micromatrizz[26][473] = 9'b111111111;
assign micromatrizz[26][474] = 9'b111111111;
assign micromatrizz[26][475] = 9'b111111111;
assign micromatrizz[26][476] = 9'b111111111;
assign micromatrizz[26][477] = 9'b111111111;
assign micromatrizz[26][478] = 9'b111111111;
assign micromatrizz[26][479] = 9'b111111111;
assign micromatrizz[26][480] = 9'b111111111;
assign micromatrizz[26][481] = 9'b111111111;
assign micromatrizz[26][482] = 9'b111111111;
assign micromatrizz[26][483] = 9'b111111111;
assign micromatrizz[26][484] = 9'b111111111;
assign micromatrizz[26][485] = 9'b111111111;
assign micromatrizz[26][486] = 9'b111111111;
assign micromatrizz[26][487] = 9'b111111111;
assign micromatrizz[26][488] = 9'b111111111;
assign micromatrizz[26][489] = 9'b111111111;
assign micromatrizz[26][490] = 9'b111111111;
assign micromatrizz[26][491] = 9'b111111111;
assign micromatrizz[26][492] = 9'b111111111;
assign micromatrizz[26][493] = 9'b111111111;
assign micromatrizz[26][494] = 9'b111111111;
assign micromatrizz[26][495] = 9'b111111111;
assign micromatrizz[26][496] = 9'b111111111;
assign micromatrizz[26][497] = 9'b111111111;
assign micromatrizz[26][498] = 9'b111111111;
assign micromatrizz[26][499] = 9'b111111111;
assign micromatrizz[26][500] = 9'b111111111;
assign micromatrizz[26][501] = 9'b111111111;
assign micromatrizz[26][502] = 9'b111111111;
assign micromatrizz[26][503] = 9'b111111111;
assign micromatrizz[26][504] = 9'b111111111;
assign micromatrizz[26][505] = 9'b111111111;
assign micromatrizz[26][506] = 9'b111111111;
assign micromatrizz[26][507] = 9'b111111111;
assign micromatrizz[26][508] = 9'b111111111;
assign micromatrizz[26][509] = 9'b111111111;
assign micromatrizz[26][510] = 9'b111111111;
assign micromatrizz[26][511] = 9'b111111111;
assign micromatrizz[26][512] = 9'b111111111;
assign micromatrizz[26][513] = 9'b111111111;
assign micromatrizz[26][514] = 9'b111111111;
assign micromatrizz[26][515] = 9'b111111111;
assign micromatrizz[26][516] = 9'b111111111;
assign micromatrizz[26][517] = 9'b111111111;
assign micromatrizz[26][518] = 9'b111111111;
assign micromatrizz[26][519] = 9'b111111111;
assign micromatrizz[26][520] = 9'b111111111;
assign micromatrizz[26][521] = 9'b111111111;
assign micromatrizz[26][522] = 9'b111111111;
assign micromatrizz[26][523] = 9'b111111111;
assign micromatrizz[26][524] = 9'b111111111;
assign micromatrizz[26][525] = 9'b111111111;
assign micromatrizz[26][526] = 9'b111111111;
assign micromatrizz[26][527] = 9'b111111111;
assign micromatrizz[26][528] = 9'b111111111;
assign micromatrizz[26][529] = 9'b111111111;
assign micromatrizz[26][530] = 9'b111111111;
assign micromatrizz[26][531] = 9'b111111111;
assign micromatrizz[26][532] = 9'b111111111;
assign micromatrizz[26][533] = 9'b111111111;
assign micromatrizz[26][534] = 9'b111111111;
assign micromatrizz[26][535] = 9'b111111111;
assign micromatrizz[26][536] = 9'b111111111;
assign micromatrizz[26][537] = 9'b111111111;
assign micromatrizz[26][538] = 9'b111111111;
assign micromatrizz[26][539] = 9'b111111111;
assign micromatrizz[26][540] = 9'b111111111;
assign micromatrizz[26][541] = 9'b111111111;
assign micromatrizz[26][542] = 9'b111111111;
assign micromatrizz[26][543] = 9'b111111111;
assign micromatrizz[26][544] = 9'b111111111;
assign micromatrizz[26][545] = 9'b111111111;
assign micromatrizz[26][546] = 9'b111111111;
assign micromatrizz[26][547] = 9'b111111111;
assign micromatrizz[26][548] = 9'b111111111;
assign micromatrizz[26][549] = 9'b111111111;
assign micromatrizz[26][550] = 9'b111111111;
assign micromatrizz[26][551] = 9'b111111111;
assign micromatrizz[26][552] = 9'b111111111;
assign micromatrizz[26][553] = 9'b111111111;
assign micromatrizz[26][554] = 9'b111111111;
assign micromatrizz[26][555] = 9'b111111111;
assign micromatrizz[26][556] = 9'b111111111;
assign micromatrizz[26][557] = 9'b111111111;
assign micromatrizz[26][558] = 9'b111111111;
assign micromatrizz[26][559] = 9'b111111111;
assign micromatrizz[26][560] = 9'b111111111;
assign micromatrizz[26][561] = 9'b111111111;
assign micromatrizz[26][562] = 9'b111111111;
assign micromatrizz[26][563] = 9'b111111111;
assign micromatrizz[26][564] = 9'b111111111;
assign micromatrizz[26][565] = 9'b111111111;
assign micromatrizz[26][566] = 9'b111111111;
assign micromatrizz[26][567] = 9'b111111111;
assign micromatrizz[26][568] = 9'b111111111;
assign micromatrizz[26][569] = 9'b111111111;
assign micromatrizz[26][570] = 9'b111111111;
assign micromatrizz[26][571] = 9'b111111111;
assign micromatrizz[26][572] = 9'b111111111;
assign micromatrizz[26][573] = 9'b111111111;
assign micromatrizz[26][574] = 9'b111111111;
assign micromatrizz[26][575] = 9'b111111111;
assign micromatrizz[26][576] = 9'b111111111;
assign micromatrizz[26][577] = 9'b111111111;
assign micromatrizz[26][578] = 9'b111111111;
assign micromatrizz[26][579] = 9'b111111111;
assign micromatrizz[26][580] = 9'b111111111;
assign micromatrizz[26][581] = 9'b111111111;
assign micromatrizz[26][582] = 9'b111111111;
assign micromatrizz[26][583] = 9'b111111111;
assign micromatrizz[26][584] = 9'b111111111;
assign micromatrizz[26][585] = 9'b111111111;
assign micromatrizz[26][586] = 9'b111111111;
assign micromatrizz[26][587] = 9'b111111111;
assign micromatrizz[26][588] = 9'b111111111;
assign micromatrizz[26][589] = 9'b111111111;
assign micromatrizz[26][590] = 9'b111111111;
assign micromatrizz[26][591] = 9'b111111111;
assign micromatrizz[26][592] = 9'b111111111;
assign micromatrizz[26][593] = 9'b111111111;
assign micromatrizz[26][594] = 9'b111111111;
assign micromatrizz[26][595] = 9'b111111111;
assign micromatrizz[26][596] = 9'b111111111;
assign micromatrizz[26][597] = 9'b111111111;
assign micromatrizz[26][598] = 9'b111111111;
assign micromatrizz[26][599] = 9'b111111111;
assign micromatrizz[26][600] = 9'b111111111;
assign micromatrizz[26][601] = 9'b111111111;
assign micromatrizz[26][602] = 9'b111111111;
assign micromatrizz[26][603] = 9'b111111111;
assign micromatrizz[26][604] = 9'b111111111;
assign micromatrizz[26][605] = 9'b111111111;
assign micromatrizz[26][606] = 9'b111111111;
assign micromatrizz[26][607] = 9'b111111111;
assign micromatrizz[26][608] = 9'b111111111;
assign micromatrizz[26][609] = 9'b111111111;
assign micromatrizz[26][610] = 9'b111111111;
assign micromatrizz[26][611] = 9'b111111111;
assign micromatrizz[26][612] = 9'b111111111;
assign micromatrizz[26][613] = 9'b111111111;
assign micromatrizz[26][614] = 9'b111111111;
assign micromatrizz[26][615] = 9'b111111111;
assign micromatrizz[26][616] = 9'b111111111;
assign micromatrizz[26][617] = 9'b111111111;
assign micromatrizz[26][618] = 9'b111111111;
assign micromatrizz[26][619] = 9'b111111111;
assign micromatrizz[26][620] = 9'b111111111;
assign micromatrizz[26][621] = 9'b111111111;
assign micromatrizz[26][622] = 9'b111111111;
assign micromatrizz[26][623] = 9'b111111111;
assign micromatrizz[26][624] = 9'b111111111;
assign micromatrizz[26][625] = 9'b111111111;
assign micromatrizz[26][626] = 9'b111111111;
assign micromatrizz[26][627] = 9'b111111111;
assign micromatrizz[26][628] = 9'b111111111;
assign micromatrizz[26][629] = 9'b111111111;
assign micromatrizz[26][630] = 9'b111111111;
assign micromatrizz[26][631] = 9'b111111111;
assign micromatrizz[26][632] = 9'b111111111;
assign micromatrizz[26][633] = 9'b111111111;
assign micromatrizz[26][634] = 9'b111111111;
assign micromatrizz[26][635] = 9'b111111111;
assign micromatrizz[26][636] = 9'b111111111;
assign micromatrizz[26][637] = 9'b111111111;
assign micromatrizz[26][638] = 9'b111111111;
assign micromatrizz[26][639] = 9'b111111111;
assign micromatrizz[27][0] = 9'b111111111;
assign micromatrizz[27][1] = 9'b111111111;
assign micromatrizz[27][2] = 9'b111111111;
assign micromatrizz[27][3] = 9'b111111111;
assign micromatrizz[27][4] = 9'b111111111;
assign micromatrizz[27][5] = 9'b111111111;
assign micromatrizz[27][6] = 9'b111111111;
assign micromatrizz[27][7] = 9'b111111111;
assign micromatrizz[27][8] = 9'b111111111;
assign micromatrizz[27][9] = 9'b111111111;
assign micromatrizz[27][10] = 9'b111111111;
assign micromatrizz[27][11] = 9'b111111111;
assign micromatrizz[27][12] = 9'b111111111;
assign micromatrizz[27][13] = 9'b111111111;
assign micromatrizz[27][14] = 9'b111111111;
assign micromatrizz[27][15] = 9'b111111111;
assign micromatrizz[27][16] = 9'b111111111;
assign micromatrizz[27][17] = 9'b111111111;
assign micromatrizz[27][18] = 9'b111111111;
assign micromatrizz[27][19] = 9'b111111111;
assign micromatrizz[27][20] = 9'b111111111;
assign micromatrizz[27][21] = 9'b111111111;
assign micromatrizz[27][22] = 9'b111111111;
assign micromatrizz[27][23] = 9'b111111111;
assign micromatrizz[27][24] = 9'b111111111;
assign micromatrizz[27][25] = 9'b111111111;
assign micromatrizz[27][26] = 9'b111111111;
assign micromatrizz[27][27] = 9'b111111111;
assign micromatrizz[27][28] = 9'b111111111;
assign micromatrizz[27][29] = 9'b111111111;
assign micromatrizz[27][30] = 9'b111111111;
assign micromatrizz[27][31] = 9'b111111111;
assign micromatrizz[27][32] = 9'b111111111;
assign micromatrizz[27][33] = 9'b111111111;
assign micromatrizz[27][34] = 9'b111111111;
assign micromatrizz[27][35] = 9'b111111111;
assign micromatrizz[27][36] = 9'b111111111;
assign micromatrizz[27][37] = 9'b111111111;
assign micromatrizz[27][38] = 9'b111111111;
assign micromatrizz[27][39] = 9'b111111111;
assign micromatrizz[27][40] = 9'b111111111;
assign micromatrizz[27][41] = 9'b111111111;
assign micromatrizz[27][42] = 9'b111111111;
assign micromatrizz[27][43] = 9'b111111111;
assign micromatrizz[27][44] = 9'b111111111;
assign micromatrizz[27][45] = 9'b111111111;
assign micromatrizz[27][46] = 9'b111111111;
assign micromatrizz[27][47] = 9'b111111111;
assign micromatrizz[27][48] = 9'b111111111;
assign micromatrizz[27][49] = 9'b111111111;
assign micromatrizz[27][50] = 9'b111111111;
assign micromatrizz[27][51] = 9'b111111111;
assign micromatrizz[27][52] = 9'b111111111;
assign micromatrizz[27][53] = 9'b111111111;
assign micromatrizz[27][54] = 9'b111111111;
assign micromatrizz[27][55] = 9'b111111111;
assign micromatrizz[27][56] = 9'b111111111;
assign micromatrizz[27][57] = 9'b111111111;
assign micromatrizz[27][58] = 9'b111111111;
assign micromatrizz[27][59] = 9'b111111111;
assign micromatrizz[27][60] = 9'b111111111;
assign micromatrizz[27][61] = 9'b111111111;
assign micromatrizz[27][62] = 9'b111111111;
assign micromatrizz[27][63] = 9'b111111111;
assign micromatrizz[27][64] = 9'b111111111;
assign micromatrizz[27][65] = 9'b111111111;
assign micromatrizz[27][66] = 9'b111111111;
assign micromatrizz[27][67] = 9'b111111111;
assign micromatrizz[27][68] = 9'b111111111;
assign micromatrizz[27][69] = 9'b111111111;
assign micromatrizz[27][70] = 9'b111111111;
assign micromatrizz[27][71] = 9'b111111111;
assign micromatrizz[27][72] = 9'b111111111;
assign micromatrizz[27][73] = 9'b111111111;
assign micromatrizz[27][74] = 9'b111111111;
assign micromatrizz[27][75] = 9'b111111111;
assign micromatrizz[27][76] = 9'b111111111;
assign micromatrizz[27][77] = 9'b111111111;
assign micromatrizz[27][78] = 9'b111111111;
assign micromatrizz[27][79] = 9'b111111111;
assign micromatrizz[27][80] = 9'b111111111;
assign micromatrizz[27][81] = 9'b111111111;
assign micromatrizz[27][82] = 9'b111111111;
assign micromatrizz[27][83] = 9'b111111111;
assign micromatrizz[27][84] = 9'b111111111;
assign micromatrizz[27][85] = 9'b111111111;
assign micromatrizz[27][86] = 9'b111111111;
assign micromatrizz[27][87] = 9'b111111111;
assign micromatrizz[27][88] = 9'b111111111;
assign micromatrizz[27][89] = 9'b111111111;
assign micromatrizz[27][90] = 9'b111111111;
assign micromatrizz[27][91] = 9'b111111111;
assign micromatrizz[27][92] = 9'b111111111;
assign micromatrizz[27][93] = 9'b111111111;
assign micromatrizz[27][94] = 9'b111111111;
assign micromatrizz[27][95] = 9'b111111111;
assign micromatrizz[27][96] = 9'b111111111;
assign micromatrizz[27][97] = 9'b111111111;
assign micromatrizz[27][98] = 9'b111111111;
assign micromatrizz[27][99] = 9'b111111111;
assign micromatrizz[27][100] = 9'b111111111;
assign micromatrizz[27][101] = 9'b111111111;
assign micromatrizz[27][102] = 9'b111111111;
assign micromatrizz[27][103] = 9'b111111111;
assign micromatrizz[27][104] = 9'b111111111;
assign micromatrizz[27][105] = 9'b111111111;
assign micromatrizz[27][106] = 9'b111111111;
assign micromatrizz[27][107] = 9'b111111111;
assign micromatrizz[27][108] = 9'b111111111;
assign micromatrizz[27][109] = 9'b111111111;
assign micromatrizz[27][110] = 9'b111111111;
assign micromatrizz[27][111] = 9'b111111111;
assign micromatrizz[27][112] = 9'b111111111;
assign micromatrizz[27][113] = 9'b111111111;
assign micromatrizz[27][114] = 9'b111111111;
assign micromatrizz[27][115] = 9'b111111111;
assign micromatrizz[27][116] = 9'b111111111;
assign micromatrizz[27][117] = 9'b111111111;
assign micromatrizz[27][118] = 9'b111111111;
assign micromatrizz[27][119] = 9'b111111111;
assign micromatrizz[27][120] = 9'b111111111;
assign micromatrizz[27][121] = 9'b111111111;
assign micromatrizz[27][122] = 9'b111111111;
assign micromatrizz[27][123] = 9'b111111111;
assign micromatrizz[27][124] = 9'b111111111;
assign micromatrizz[27][125] = 9'b111111111;
assign micromatrizz[27][126] = 9'b111111111;
assign micromatrizz[27][127] = 9'b111111111;
assign micromatrizz[27][128] = 9'b111111111;
assign micromatrizz[27][129] = 9'b111111111;
assign micromatrizz[27][130] = 9'b111111111;
assign micromatrizz[27][131] = 9'b111111111;
assign micromatrizz[27][132] = 9'b111111111;
assign micromatrizz[27][133] = 9'b111111111;
assign micromatrizz[27][134] = 9'b111111111;
assign micromatrizz[27][135] = 9'b111111111;
assign micromatrizz[27][136] = 9'b111111111;
assign micromatrizz[27][137] = 9'b111111111;
assign micromatrizz[27][138] = 9'b111111111;
assign micromatrizz[27][139] = 9'b111111111;
assign micromatrizz[27][140] = 9'b111111111;
assign micromatrizz[27][141] = 9'b111111111;
assign micromatrizz[27][142] = 9'b111111111;
assign micromatrizz[27][143] = 9'b111111111;
assign micromatrizz[27][144] = 9'b111111111;
assign micromatrizz[27][145] = 9'b111111111;
assign micromatrizz[27][146] = 9'b111111111;
assign micromatrizz[27][147] = 9'b111111111;
assign micromatrizz[27][148] = 9'b111111111;
assign micromatrizz[27][149] = 9'b111111111;
assign micromatrizz[27][150] = 9'b111111111;
assign micromatrizz[27][151] = 9'b111111111;
assign micromatrizz[27][152] = 9'b111111111;
assign micromatrizz[27][153] = 9'b111111111;
assign micromatrizz[27][154] = 9'b111111111;
assign micromatrizz[27][155] = 9'b111111111;
assign micromatrizz[27][156] = 9'b111111111;
assign micromatrizz[27][157] = 9'b111111111;
assign micromatrizz[27][158] = 9'b111111111;
assign micromatrizz[27][159] = 9'b111111111;
assign micromatrizz[27][160] = 9'b111111111;
assign micromatrizz[27][161] = 9'b111111111;
assign micromatrizz[27][162] = 9'b111111111;
assign micromatrizz[27][163] = 9'b111111111;
assign micromatrizz[27][164] = 9'b111111111;
assign micromatrizz[27][165] = 9'b111111111;
assign micromatrizz[27][166] = 9'b111111111;
assign micromatrizz[27][167] = 9'b111111111;
assign micromatrizz[27][168] = 9'b111111111;
assign micromatrizz[27][169] = 9'b111111111;
assign micromatrizz[27][170] = 9'b111111111;
assign micromatrizz[27][171] = 9'b111111111;
assign micromatrizz[27][172] = 9'b111111111;
assign micromatrizz[27][173] = 9'b111111111;
assign micromatrizz[27][174] = 9'b111111111;
assign micromatrizz[27][175] = 9'b111111111;
assign micromatrizz[27][176] = 9'b111111111;
assign micromatrizz[27][177] = 9'b111111111;
assign micromatrizz[27][178] = 9'b111111111;
assign micromatrizz[27][179] = 9'b111111111;
assign micromatrizz[27][180] = 9'b111111111;
assign micromatrizz[27][181] = 9'b111111111;
assign micromatrizz[27][182] = 9'b111111111;
assign micromatrizz[27][183] = 9'b111111111;
assign micromatrizz[27][184] = 9'b111111111;
assign micromatrizz[27][185] = 9'b111111111;
assign micromatrizz[27][186] = 9'b111111111;
assign micromatrizz[27][187] = 9'b111111111;
assign micromatrizz[27][188] = 9'b111111111;
assign micromatrizz[27][189] = 9'b111111111;
assign micromatrizz[27][190] = 9'b111111111;
assign micromatrizz[27][191] = 9'b111111111;
assign micromatrizz[27][192] = 9'b111111111;
assign micromatrizz[27][193] = 9'b111111111;
assign micromatrizz[27][194] = 9'b111111111;
assign micromatrizz[27][195] = 9'b111111111;
assign micromatrizz[27][196] = 9'b111111111;
assign micromatrizz[27][197] = 9'b111111111;
assign micromatrizz[27][198] = 9'b111111111;
assign micromatrizz[27][199] = 9'b111111111;
assign micromatrizz[27][200] = 9'b111111111;
assign micromatrizz[27][201] = 9'b111111111;
assign micromatrizz[27][202] = 9'b111111111;
assign micromatrizz[27][203] = 9'b111111111;
assign micromatrizz[27][204] = 9'b111111111;
assign micromatrizz[27][205] = 9'b111111111;
assign micromatrizz[27][206] = 9'b111111111;
assign micromatrizz[27][207] = 9'b111111111;
assign micromatrizz[27][208] = 9'b111111111;
assign micromatrizz[27][209] = 9'b111111111;
assign micromatrizz[27][210] = 9'b111111111;
assign micromatrizz[27][211] = 9'b111111111;
assign micromatrizz[27][212] = 9'b111111111;
assign micromatrizz[27][213] = 9'b111111111;
assign micromatrizz[27][214] = 9'b111111111;
assign micromatrizz[27][215] = 9'b111111111;
assign micromatrizz[27][216] = 9'b111111111;
assign micromatrizz[27][217] = 9'b111111111;
assign micromatrizz[27][218] = 9'b111111111;
assign micromatrizz[27][219] = 9'b111111111;
assign micromatrizz[27][220] = 9'b111111111;
assign micromatrizz[27][221] = 9'b111111111;
assign micromatrizz[27][222] = 9'b111111111;
assign micromatrizz[27][223] = 9'b111111111;
assign micromatrizz[27][224] = 9'b111111111;
assign micromatrizz[27][225] = 9'b111111111;
assign micromatrizz[27][226] = 9'b111111111;
assign micromatrizz[27][227] = 9'b111111111;
assign micromatrizz[27][228] = 9'b111111111;
assign micromatrizz[27][229] = 9'b111111111;
assign micromatrizz[27][230] = 9'b111111111;
assign micromatrizz[27][231] = 9'b111111111;
assign micromatrizz[27][232] = 9'b111111111;
assign micromatrizz[27][233] = 9'b111111111;
assign micromatrizz[27][234] = 9'b111111111;
assign micromatrizz[27][235] = 9'b111111111;
assign micromatrizz[27][236] = 9'b111111111;
assign micromatrizz[27][237] = 9'b111111111;
assign micromatrizz[27][238] = 9'b111111111;
assign micromatrizz[27][239] = 9'b111111111;
assign micromatrizz[27][240] = 9'b111111111;
assign micromatrizz[27][241] = 9'b111111111;
assign micromatrizz[27][242] = 9'b111111111;
assign micromatrizz[27][243] = 9'b111111111;
assign micromatrizz[27][244] = 9'b111111111;
assign micromatrizz[27][245] = 9'b111111111;
assign micromatrizz[27][246] = 9'b111111111;
assign micromatrizz[27][247] = 9'b111111111;
assign micromatrizz[27][248] = 9'b111111111;
assign micromatrizz[27][249] = 9'b111111111;
assign micromatrizz[27][250] = 9'b111111111;
assign micromatrizz[27][251] = 9'b111111111;
assign micromatrizz[27][252] = 9'b111111111;
assign micromatrizz[27][253] = 9'b111111111;
assign micromatrizz[27][254] = 9'b111111111;
assign micromatrizz[27][255] = 9'b111111111;
assign micromatrizz[27][256] = 9'b111111111;
assign micromatrizz[27][257] = 9'b111111111;
assign micromatrizz[27][258] = 9'b111111111;
assign micromatrizz[27][259] = 9'b111111111;
assign micromatrizz[27][260] = 9'b111111111;
assign micromatrizz[27][261] = 9'b111111111;
assign micromatrizz[27][262] = 9'b111111111;
assign micromatrizz[27][263] = 9'b111111111;
assign micromatrizz[27][264] = 9'b111111111;
assign micromatrizz[27][265] = 9'b111111111;
assign micromatrizz[27][266] = 9'b111111111;
assign micromatrizz[27][267] = 9'b111111111;
assign micromatrizz[27][268] = 9'b111111111;
assign micromatrizz[27][269] = 9'b111111111;
assign micromatrizz[27][270] = 9'b111110010;
assign micromatrizz[27][271] = 9'b111110010;
assign micromatrizz[27][272] = 9'b111110010;
assign micromatrizz[27][273] = 9'b111110011;
assign micromatrizz[27][274] = 9'b111110011;
assign micromatrizz[27][275] = 9'b111110011;
assign micromatrizz[27][276] = 9'b111110011;
assign micromatrizz[27][277] = 9'b111110011;
assign micromatrizz[27][278] = 9'b111110011;
assign micromatrizz[27][279] = 9'b111111111;
assign micromatrizz[27][280] = 9'b111111111;
assign micromatrizz[27][281] = 9'b111111111;
assign micromatrizz[27][282] = 9'b111111111;
assign micromatrizz[27][283] = 9'b111111111;
assign micromatrizz[27][284] = 9'b111111111;
assign micromatrizz[27][285] = 9'b111111111;
assign micromatrizz[27][286] = 9'b111111111;
assign micromatrizz[27][287] = 9'b111111111;
assign micromatrizz[27][288] = 9'b111111111;
assign micromatrizz[27][289] = 9'b111111111;
assign micromatrizz[27][290] = 9'b111110111;
assign micromatrizz[27][291] = 9'b111110010;
assign micromatrizz[27][292] = 9'b111110010;
assign micromatrizz[27][293] = 9'b111110011;
assign micromatrizz[27][294] = 9'b111110011;
assign micromatrizz[27][295] = 9'b111110011;
assign micromatrizz[27][296] = 9'b111110011;
assign micromatrizz[27][297] = 9'b111110111;
assign micromatrizz[27][298] = 9'b111111111;
assign micromatrizz[27][299] = 9'b111111111;
assign micromatrizz[27][300] = 9'b111111111;
assign micromatrizz[27][301] = 9'b111111111;
assign micromatrizz[27][302] = 9'b111111111;
assign micromatrizz[27][303] = 9'b111111111;
assign micromatrizz[27][304] = 9'b111111111;
assign micromatrizz[27][305] = 9'b111110010;
assign micromatrizz[27][306] = 9'b111111111;
assign micromatrizz[27][307] = 9'b111111111;
assign micromatrizz[27][308] = 9'b111110111;
assign micromatrizz[27][309] = 9'b111110010;
assign micromatrizz[27][310] = 9'b111110010;
assign micromatrizz[27][311] = 9'b111110011;
assign micromatrizz[27][312] = 9'b111110011;
assign micromatrizz[27][313] = 9'b111110010;
assign micromatrizz[27][314] = 9'b111110011;
assign micromatrizz[27][315] = 9'b111110011;
assign micromatrizz[27][316] = 9'b111110011;
assign micromatrizz[27][317] = 9'b111111111;
assign micromatrizz[27][318] = 9'b111111111;
assign micromatrizz[27][319] = 9'b111111111;
assign micromatrizz[27][320] = 9'b111111111;
assign micromatrizz[27][321] = 9'b111111111;
assign micromatrizz[27][322] = 9'b111111111;
assign micromatrizz[27][323] = 9'b111111111;
assign micromatrizz[27][324] = 9'b111111111;
assign micromatrizz[27][325] = 9'b111111111;
assign micromatrizz[27][326] = 9'b111111111;
assign micromatrizz[27][327] = 9'b111111111;
assign micromatrizz[27][328] = 9'b111111111;
assign micromatrizz[27][329] = 9'b111111111;
assign micromatrizz[27][330] = 9'b111111111;
assign micromatrizz[27][331] = 9'b111111111;
assign micromatrizz[27][332] = 9'b111111111;
assign micromatrizz[27][333] = 9'b111111111;
assign micromatrizz[27][334] = 9'b111111111;
assign micromatrizz[27][335] = 9'b111111111;
assign micromatrizz[27][336] = 9'b111111111;
assign micromatrizz[27][337] = 9'b111111111;
assign micromatrizz[27][338] = 9'b111111111;
assign micromatrizz[27][339] = 9'b111111111;
assign micromatrizz[27][340] = 9'b111111111;
assign micromatrizz[27][341] = 9'b111111111;
assign micromatrizz[27][342] = 9'b111111111;
assign micromatrizz[27][343] = 9'b111111111;
assign micromatrizz[27][344] = 9'b111111111;
assign micromatrizz[27][345] = 9'b111111111;
assign micromatrizz[27][346] = 9'b111111111;
assign micromatrizz[27][347] = 9'b111111111;
assign micromatrizz[27][348] = 9'b111111111;
assign micromatrizz[27][349] = 9'b111111111;
assign micromatrizz[27][350] = 9'b111111111;
assign micromatrizz[27][351] = 9'b111111111;
assign micromatrizz[27][352] = 9'b111111111;
assign micromatrizz[27][353] = 9'b111111111;
assign micromatrizz[27][354] = 9'b111111111;
assign micromatrizz[27][355] = 9'b111111111;
assign micromatrizz[27][356] = 9'b111111111;
assign micromatrizz[27][357] = 9'b111111111;
assign micromatrizz[27][358] = 9'b111111111;
assign micromatrizz[27][359] = 9'b111111111;
assign micromatrizz[27][360] = 9'b111111111;
assign micromatrizz[27][361] = 9'b111111111;
assign micromatrizz[27][362] = 9'b111111111;
assign micromatrizz[27][363] = 9'b111111111;
assign micromatrizz[27][364] = 9'b111111111;
assign micromatrizz[27][365] = 9'b111111111;
assign micromatrizz[27][366] = 9'b111111111;
assign micromatrizz[27][367] = 9'b111111111;
assign micromatrizz[27][368] = 9'b111111111;
assign micromatrizz[27][369] = 9'b111111111;
assign micromatrizz[27][370] = 9'b111111111;
assign micromatrizz[27][371] = 9'b111111111;
assign micromatrizz[27][372] = 9'b111111111;
assign micromatrizz[27][373] = 9'b111111111;
assign micromatrizz[27][374] = 9'b111111111;
assign micromatrizz[27][375] = 9'b111111111;
assign micromatrizz[27][376] = 9'b111111111;
assign micromatrizz[27][377] = 9'b111111111;
assign micromatrizz[27][378] = 9'b111111111;
assign micromatrizz[27][379] = 9'b111111111;
assign micromatrizz[27][380] = 9'b111111111;
assign micromatrizz[27][381] = 9'b111111111;
assign micromatrizz[27][382] = 9'b111111111;
assign micromatrizz[27][383] = 9'b111111111;
assign micromatrizz[27][384] = 9'b111111111;
assign micromatrizz[27][385] = 9'b111111111;
assign micromatrizz[27][386] = 9'b111111111;
assign micromatrizz[27][387] = 9'b111111111;
assign micromatrizz[27][388] = 9'b111111111;
assign micromatrizz[27][389] = 9'b111111111;
assign micromatrizz[27][390] = 9'b111111111;
assign micromatrizz[27][391] = 9'b111111111;
assign micromatrizz[27][392] = 9'b111111111;
assign micromatrizz[27][393] = 9'b111111111;
assign micromatrizz[27][394] = 9'b111111111;
assign micromatrizz[27][395] = 9'b111111111;
assign micromatrizz[27][396] = 9'b111111111;
assign micromatrizz[27][397] = 9'b111111111;
assign micromatrizz[27][398] = 9'b111111111;
assign micromatrizz[27][399] = 9'b111111111;
assign micromatrizz[27][400] = 9'b111111111;
assign micromatrizz[27][401] = 9'b111111111;
assign micromatrizz[27][402] = 9'b111111111;
assign micromatrizz[27][403] = 9'b111111111;
assign micromatrizz[27][404] = 9'b111111111;
assign micromatrizz[27][405] = 9'b111111111;
assign micromatrizz[27][406] = 9'b111111111;
assign micromatrizz[27][407] = 9'b111111111;
assign micromatrizz[27][408] = 9'b111111111;
assign micromatrizz[27][409] = 9'b111111111;
assign micromatrizz[27][410] = 9'b111111111;
assign micromatrizz[27][411] = 9'b111111111;
assign micromatrizz[27][412] = 9'b111111111;
assign micromatrizz[27][413] = 9'b111111111;
assign micromatrizz[27][414] = 9'b111111111;
assign micromatrizz[27][415] = 9'b111111111;
assign micromatrizz[27][416] = 9'b111111111;
assign micromatrizz[27][417] = 9'b111111111;
assign micromatrizz[27][418] = 9'b111111111;
assign micromatrizz[27][419] = 9'b111111111;
assign micromatrizz[27][420] = 9'b111111111;
assign micromatrizz[27][421] = 9'b111111111;
assign micromatrizz[27][422] = 9'b111111111;
assign micromatrizz[27][423] = 9'b111111111;
assign micromatrizz[27][424] = 9'b111111111;
assign micromatrizz[27][425] = 9'b111111111;
assign micromatrizz[27][426] = 9'b111111111;
assign micromatrizz[27][427] = 9'b111111111;
assign micromatrizz[27][428] = 9'b111111111;
assign micromatrizz[27][429] = 9'b111111111;
assign micromatrizz[27][430] = 9'b111111111;
assign micromatrizz[27][431] = 9'b111111111;
assign micromatrizz[27][432] = 9'b111111111;
assign micromatrizz[27][433] = 9'b111111111;
assign micromatrizz[27][434] = 9'b111111111;
assign micromatrizz[27][435] = 9'b111111111;
assign micromatrizz[27][436] = 9'b111111111;
assign micromatrizz[27][437] = 9'b111111111;
assign micromatrizz[27][438] = 9'b111111111;
assign micromatrizz[27][439] = 9'b111111111;
assign micromatrizz[27][440] = 9'b111111111;
assign micromatrizz[27][441] = 9'b111111111;
assign micromatrizz[27][442] = 9'b111111111;
assign micromatrizz[27][443] = 9'b111111111;
assign micromatrizz[27][444] = 9'b111111111;
assign micromatrizz[27][445] = 9'b111111111;
assign micromatrizz[27][446] = 9'b111111111;
assign micromatrizz[27][447] = 9'b111111111;
assign micromatrizz[27][448] = 9'b111111111;
assign micromatrizz[27][449] = 9'b111111111;
assign micromatrizz[27][450] = 9'b111111111;
assign micromatrizz[27][451] = 9'b111111111;
assign micromatrizz[27][452] = 9'b111111111;
assign micromatrizz[27][453] = 9'b111111111;
assign micromatrizz[27][454] = 9'b111111111;
assign micromatrizz[27][455] = 9'b111111111;
assign micromatrizz[27][456] = 9'b111111111;
assign micromatrizz[27][457] = 9'b111111111;
assign micromatrizz[27][458] = 9'b111111111;
assign micromatrizz[27][459] = 9'b111111111;
assign micromatrizz[27][460] = 9'b111111111;
assign micromatrizz[27][461] = 9'b111111111;
assign micromatrizz[27][462] = 9'b111111111;
assign micromatrizz[27][463] = 9'b111111111;
assign micromatrizz[27][464] = 9'b111111111;
assign micromatrizz[27][465] = 9'b111111111;
assign micromatrizz[27][466] = 9'b111111111;
assign micromatrizz[27][467] = 9'b111111111;
assign micromatrizz[27][468] = 9'b111111111;
assign micromatrizz[27][469] = 9'b111111111;
assign micromatrizz[27][470] = 9'b111111111;
assign micromatrizz[27][471] = 9'b111111111;
assign micromatrizz[27][472] = 9'b111111111;
assign micromatrizz[27][473] = 9'b111111111;
assign micromatrizz[27][474] = 9'b111111111;
assign micromatrizz[27][475] = 9'b111111111;
assign micromatrizz[27][476] = 9'b111111111;
assign micromatrizz[27][477] = 9'b111111111;
assign micromatrizz[27][478] = 9'b111111111;
assign micromatrizz[27][479] = 9'b111111111;
assign micromatrizz[27][480] = 9'b111111111;
assign micromatrizz[27][481] = 9'b111111111;
assign micromatrizz[27][482] = 9'b111111111;
assign micromatrizz[27][483] = 9'b111111111;
assign micromatrizz[27][484] = 9'b111111111;
assign micromatrizz[27][485] = 9'b111111111;
assign micromatrizz[27][486] = 9'b111111111;
assign micromatrizz[27][487] = 9'b111111111;
assign micromatrizz[27][488] = 9'b111111111;
assign micromatrizz[27][489] = 9'b111111111;
assign micromatrizz[27][490] = 9'b111111111;
assign micromatrizz[27][491] = 9'b111111111;
assign micromatrizz[27][492] = 9'b111111111;
assign micromatrizz[27][493] = 9'b111111111;
assign micromatrizz[27][494] = 9'b111111111;
assign micromatrizz[27][495] = 9'b111111111;
assign micromatrizz[27][496] = 9'b111111111;
assign micromatrizz[27][497] = 9'b111111111;
assign micromatrizz[27][498] = 9'b111111111;
assign micromatrizz[27][499] = 9'b111111111;
assign micromatrizz[27][500] = 9'b111111111;
assign micromatrizz[27][501] = 9'b111111111;
assign micromatrizz[27][502] = 9'b111111111;
assign micromatrizz[27][503] = 9'b111111111;
assign micromatrizz[27][504] = 9'b111111111;
assign micromatrizz[27][505] = 9'b111111111;
assign micromatrizz[27][506] = 9'b111111111;
assign micromatrizz[27][507] = 9'b111111111;
assign micromatrizz[27][508] = 9'b111111111;
assign micromatrizz[27][509] = 9'b111111111;
assign micromatrizz[27][510] = 9'b111111111;
assign micromatrizz[27][511] = 9'b111111111;
assign micromatrizz[27][512] = 9'b111111111;
assign micromatrizz[27][513] = 9'b111111111;
assign micromatrizz[27][514] = 9'b111111111;
assign micromatrizz[27][515] = 9'b111111111;
assign micromatrizz[27][516] = 9'b111111111;
assign micromatrizz[27][517] = 9'b111111111;
assign micromatrizz[27][518] = 9'b111111111;
assign micromatrizz[27][519] = 9'b111111111;
assign micromatrizz[27][520] = 9'b111111111;
assign micromatrizz[27][521] = 9'b111111111;
assign micromatrizz[27][522] = 9'b111111111;
assign micromatrizz[27][523] = 9'b111111111;
assign micromatrizz[27][524] = 9'b111111111;
assign micromatrizz[27][525] = 9'b111111111;
assign micromatrizz[27][526] = 9'b111111111;
assign micromatrizz[27][527] = 9'b111111111;
assign micromatrizz[27][528] = 9'b111111111;
assign micromatrizz[27][529] = 9'b111111111;
assign micromatrizz[27][530] = 9'b111111111;
assign micromatrizz[27][531] = 9'b111111111;
assign micromatrizz[27][532] = 9'b111111111;
assign micromatrizz[27][533] = 9'b111111111;
assign micromatrizz[27][534] = 9'b111111111;
assign micromatrizz[27][535] = 9'b111111111;
assign micromatrizz[27][536] = 9'b111111111;
assign micromatrizz[27][537] = 9'b111111111;
assign micromatrizz[27][538] = 9'b111111111;
assign micromatrizz[27][539] = 9'b111111111;
assign micromatrizz[27][540] = 9'b111111111;
assign micromatrizz[27][541] = 9'b111111111;
assign micromatrizz[27][542] = 9'b111111111;
assign micromatrizz[27][543] = 9'b111111111;
assign micromatrizz[27][544] = 9'b111111111;
assign micromatrizz[27][545] = 9'b111111111;
assign micromatrizz[27][546] = 9'b111111111;
assign micromatrizz[27][547] = 9'b111111111;
assign micromatrizz[27][548] = 9'b111111111;
assign micromatrizz[27][549] = 9'b111111111;
assign micromatrizz[27][550] = 9'b111111111;
assign micromatrizz[27][551] = 9'b111111111;
assign micromatrizz[27][552] = 9'b111111111;
assign micromatrizz[27][553] = 9'b111111111;
assign micromatrizz[27][554] = 9'b111111111;
assign micromatrizz[27][555] = 9'b111111111;
assign micromatrizz[27][556] = 9'b111111111;
assign micromatrizz[27][557] = 9'b111111111;
assign micromatrizz[27][558] = 9'b111111111;
assign micromatrizz[27][559] = 9'b111111111;
assign micromatrizz[27][560] = 9'b111111111;
assign micromatrizz[27][561] = 9'b111111111;
assign micromatrizz[27][562] = 9'b111111111;
assign micromatrizz[27][563] = 9'b111111111;
assign micromatrizz[27][564] = 9'b111111111;
assign micromatrizz[27][565] = 9'b111111111;
assign micromatrizz[27][566] = 9'b111111111;
assign micromatrizz[27][567] = 9'b111111111;
assign micromatrizz[27][568] = 9'b111111111;
assign micromatrizz[27][569] = 9'b111111111;
assign micromatrizz[27][570] = 9'b111111111;
assign micromatrizz[27][571] = 9'b111111111;
assign micromatrizz[27][572] = 9'b111111111;
assign micromatrizz[27][573] = 9'b111111111;
assign micromatrizz[27][574] = 9'b111111111;
assign micromatrizz[27][575] = 9'b111111111;
assign micromatrizz[27][576] = 9'b111111111;
assign micromatrizz[27][577] = 9'b111111111;
assign micromatrizz[27][578] = 9'b111111111;
assign micromatrizz[27][579] = 9'b111111111;
assign micromatrizz[27][580] = 9'b111111111;
assign micromatrizz[27][581] = 9'b111111111;
assign micromatrizz[27][582] = 9'b111111111;
assign micromatrizz[27][583] = 9'b111111111;
assign micromatrizz[27][584] = 9'b111111111;
assign micromatrizz[27][585] = 9'b111111111;
assign micromatrizz[27][586] = 9'b111111111;
assign micromatrizz[27][587] = 9'b111111111;
assign micromatrizz[27][588] = 9'b111111111;
assign micromatrizz[27][589] = 9'b111111111;
assign micromatrizz[27][590] = 9'b111111111;
assign micromatrizz[27][591] = 9'b111111111;
assign micromatrizz[27][592] = 9'b111111111;
assign micromatrizz[27][593] = 9'b111111111;
assign micromatrizz[27][594] = 9'b111111111;
assign micromatrizz[27][595] = 9'b111111111;
assign micromatrizz[27][596] = 9'b111111111;
assign micromatrizz[27][597] = 9'b111111111;
assign micromatrizz[27][598] = 9'b111111111;
assign micromatrizz[27][599] = 9'b111111111;
assign micromatrizz[27][600] = 9'b111111111;
assign micromatrizz[27][601] = 9'b111111111;
assign micromatrizz[27][602] = 9'b111111111;
assign micromatrizz[27][603] = 9'b111111111;
assign micromatrizz[27][604] = 9'b111111111;
assign micromatrizz[27][605] = 9'b111111111;
assign micromatrizz[27][606] = 9'b111111111;
assign micromatrizz[27][607] = 9'b111111111;
assign micromatrizz[27][608] = 9'b111111111;
assign micromatrizz[27][609] = 9'b111111111;
assign micromatrizz[27][610] = 9'b111111111;
assign micromatrizz[27][611] = 9'b111111111;
assign micromatrizz[27][612] = 9'b111111111;
assign micromatrizz[27][613] = 9'b111111111;
assign micromatrizz[27][614] = 9'b111111111;
assign micromatrizz[27][615] = 9'b111111111;
assign micromatrizz[27][616] = 9'b111111111;
assign micromatrizz[27][617] = 9'b111111111;
assign micromatrizz[27][618] = 9'b111111111;
assign micromatrizz[27][619] = 9'b111111111;
assign micromatrizz[27][620] = 9'b111111111;
assign micromatrizz[27][621] = 9'b111111111;
assign micromatrizz[27][622] = 9'b111111111;
assign micromatrizz[27][623] = 9'b111111111;
assign micromatrizz[27][624] = 9'b111111111;
assign micromatrizz[27][625] = 9'b111111111;
assign micromatrizz[27][626] = 9'b111111111;
assign micromatrizz[27][627] = 9'b111111111;
assign micromatrizz[27][628] = 9'b111111111;
assign micromatrizz[27][629] = 9'b111111111;
assign micromatrizz[27][630] = 9'b111111111;
assign micromatrizz[27][631] = 9'b111111111;
assign micromatrizz[27][632] = 9'b111111111;
assign micromatrizz[27][633] = 9'b111111111;
assign micromatrizz[27][634] = 9'b111111111;
assign micromatrizz[27][635] = 9'b111111111;
assign micromatrizz[27][636] = 9'b111111111;
assign micromatrizz[27][637] = 9'b111111111;
assign micromatrizz[27][638] = 9'b111111111;
assign micromatrizz[27][639] = 9'b111111111;
assign micromatrizz[28][0] = 9'b111111111;
assign micromatrizz[28][1] = 9'b111111111;
assign micromatrizz[28][2] = 9'b111111111;
assign micromatrizz[28][3] = 9'b111111111;
assign micromatrizz[28][4] = 9'b111111111;
assign micromatrizz[28][5] = 9'b111111111;
assign micromatrizz[28][6] = 9'b111111111;
assign micromatrizz[28][7] = 9'b111111111;
assign micromatrizz[28][8] = 9'b111111111;
assign micromatrizz[28][9] = 9'b111111111;
assign micromatrizz[28][10] = 9'b111111111;
assign micromatrizz[28][11] = 9'b111111111;
assign micromatrizz[28][12] = 9'b111111111;
assign micromatrizz[28][13] = 9'b111111111;
assign micromatrizz[28][14] = 9'b111111111;
assign micromatrizz[28][15] = 9'b111111111;
assign micromatrizz[28][16] = 9'b111111111;
assign micromatrizz[28][17] = 9'b111111111;
assign micromatrizz[28][18] = 9'b111111111;
assign micromatrizz[28][19] = 9'b111111111;
assign micromatrizz[28][20] = 9'b111111111;
assign micromatrizz[28][21] = 9'b111111111;
assign micromatrizz[28][22] = 9'b111111111;
assign micromatrizz[28][23] = 9'b111111111;
assign micromatrizz[28][24] = 9'b111111111;
assign micromatrizz[28][25] = 9'b111111111;
assign micromatrizz[28][26] = 9'b111111111;
assign micromatrizz[28][27] = 9'b111111111;
assign micromatrizz[28][28] = 9'b111111111;
assign micromatrizz[28][29] = 9'b111111111;
assign micromatrizz[28][30] = 9'b111111111;
assign micromatrizz[28][31] = 9'b111111111;
assign micromatrizz[28][32] = 9'b111111111;
assign micromatrizz[28][33] = 9'b111111111;
assign micromatrizz[28][34] = 9'b111111111;
assign micromatrizz[28][35] = 9'b111111111;
assign micromatrizz[28][36] = 9'b111111111;
assign micromatrizz[28][37] = 9'b111111111;
assign micromatrizz[28][38] = 9'b111111111;
assign micromatrizz[28][39] = 9'b111111111;
assign micromatrizz[28][40] = 9'b111111111;
assign micromatrizz[28][41] = 9'b111111111;
assign micromatrizz[28][42] = 9'b111111111;
assign micromatrizz[28][43] = 9'b111111111;
assign micromatrizz[28][44] = 9'b111111111;
assign micromatrizz[28][45] = 9'b111111111;
assign micromatrizz[28][46] = 9'b111111111;
assign micromatrizz[28][47] = 9'b111111111;
assign micromatrizz[28][48] = 9'b111111111;
assign micromatrizz[28][49] = 9'b111111111;
assign micromatrizz[28][50] = 9'b111111111;
assign micromatrizz[28][51] = 9'b111111111;
assign micromatrizz[28][52] = 9'b111111111;
assign micromatrizz[28][53] = 9'b111111111;
assign micromatrizz[28][54] = 9'b111111111;
assign micromatrizz[28][55] = 9'b111111111;
assign micromatrizz[28][56] = 9'b111111111;
assign micromatrizz[28][57] = 9'b111111111;
assign micromatrizz[28][58] = 9'b111111111;
assign micromatrizz[28][59] = 9'b111111111;
assign micromatrizz[28][60] = 9'b111111111;
assign micromatrizz[28][61] = 9'b111111111;
assign micromatrizz[28][62] = 9'b111111111;
assign micromatrizz[28][63] = 9'b111111111;
assign micromatrizz[28][64] = 9'b111111111;
assign micromatrizz[28][65] = 9'b111111111;
assign micromatrizz[28][66] = 9'b111111111;
assign micromatrizz[28][67] = 9'b111111111;
assign micromatrizz[28][68] = 9'b111111111;
assign micromatrizz[28][69] = 9'b111111111;
assign micromatrizz[28][70] = 9'b111111111;
assign micromatrizz[28][71] = 9'b111111111;
assign micromatrizz[28][72] = 9'b111111111;
assign micromatrizz[28][73] = 9'b111111111;
assign micromatrizz[28][74] = 9'b111111111;
assign micromatrizz[28][75] = 9'b111111111;
assign micromatrizz[28][76] = 9'b111111111;
assign micromatrizz[28][77] = 9'b111111111;
assign micromatrizz[28][78] = 9'b111111111;
assign micromatrizz[28][79] = 9'b111111111;
assign micromatrizz[28][80] = 9'b111111111;
assign micromatrizz[28][81] = 9'b111111111;
assign micromatrizz[28][82] = 9'b111111111;
assign micromatrizz[28][83] = 9'b111111111;
assign micromatrizz[28][84] = 9'b111111111;
assign micromatrizz[28][85] = 9'b111111111;
assign micromatrizz[28][86] = 9'b111111111;
assign micromatrizz[28][87] = 9'b111111111;
assign micromatrizz[28][88] = 9'b111111111;
assign micromatrizz[28][89] = 9'b111111111;
assign micromatrizz[28][90] = 9'b111111111;
assign micromatrizz[28][91] = 9'b111111111;
assign micromatrizz[28][92] = 9'b111111111;
assign micromatrizz[28][93] = 9'b111111111;
assign micromatrizz[28][94] = 9'b111111111;
assign micromatrizz[28][95] = 9'b111111111;
assign micromatrizz[28][96] = 9'b111111111;
assign micromatrizz[28][97] = 9'b111111111;
assign micromatrizz[28][98] = 9'b111111111;
assign micromatrizz[28][99] = 9'b111111111;
assign micromatrizz[28][100] = 9'b111111111;
assign micromatrizz[28][101] = 9'b111111111;
assign micromatrizz[28][102] = 9'b111111111;
assign micromatrizz[28][103] = 9'b111111111;
assign micromatrizz[28][104] = 9'b111111111;
assign micromatrizz[28][105] = 9'b111111111;
assign micromatrizz[28][106] = 9'b111111111;
assign micromatrizz[28][107] = 9'b111111111;
assign micromatrizz[28][108] = 9'b111111111;
assign micromatrizz[28][109] = 9'b111111111;
assign micromatrizz[28][110] = 9'b111111111;
assign micromatrizz[28][111] = 9'b111111111;
assign micromatrizz[28][112] = 9'b111111111;
assign micromatrizz[28][113] = 9'b111111111;
assign micromatrizz[28][114] = 9'b111111111;
assign micromatrizz[28][115] = 9'b111111111;
assign micromatrizz[28][116] = 9'b111111111;
assign micromatrizz[28][117] = 9'b111111111;
assign micromatrizz[28][118] = 9'b111111111;
assign micromatrizz[28][119] = 9'b111111111;
assign micromatrizz[28][120] = 9'b111111111;
assign micromatrizz[28][121] = 9'b111111111;
assign micromatrizz[28][122] = 9'b111111111;
assign micromatrizz[28][123] = 9'b111111111;
assign micromatrizz[28][124] = 9'b111111111;
assign micromatrizz[28][125] = 9'b111111111;
assign micromatrizz[28][126] = 9'b111111111;
assign micromatrizz[28][127] = 9'b111111111;
assign micromatrizz[28][128] = 9'b111111111;
assign micromatrizz[28][129] = 9'b111111111;
assign micromatrizz[28][130] = 9'b111111111;
assign micromatrizz[28][131] = 9'b111111111;
assign micromatrizz[28][132] = 9'b111111111;
assign micromatrizz[28][133] = 9'b111111111;
assign micromatrizz[28][134] = 9'b111111111;
assign micromatrizz[28][135] = 9'b111111111;
assign micromatrizz[28][136] = 9'b111111111;
assign micromatrizz[28][137] = 9'b111111111;
assign micromatrizz[28][138] = 9'b111111111;
assign micromatrizz[28][139] = 9'b111111111;
assign micromatrizz[28][140] = 9'b111111111;
assign micromatrizz[28][141] = 9'b111111111;
assign micromatrizz[28][142] = 9'b111111111;
assign micromatrizz[28][143] = 9'b111111111;
assign micromatrizz[28][144] = 9'b111111111;
assign micromatrizz[28][145] = 9'b111111111;
assign micromatrizz[28][146] = 9'b111111111;
assign micromatrizz[28][147] = 9'b111111111;
assign micromatrizz[28][148] = 9'b111111111;
assign micromatrizz[28][149] = 9'b111111111;
assign micromatrizz[28][150] = 9'b111111111;
assign micromatrizz[28][151] = 9'b111111111;
assign micromatrizz[28][152] = 9'b111111111;
assign micromatrizz[28][153] = 9'b111111111;
assign micromatrizz[28][154] = 9'b111111111;
assign micromatrizz[28][155] = 9'b111111111;
assign micromatrizz[28][156] = 9'b111111111;
assign micromatrizz[28][157] = 9'b111111111;
assign micromatrizz[28][158] = 9'b111111111;
assign micromatrizz[28][159] = 9'b111111111;
assign micromatrizz[28][160] = 9'b111111111;
assign micromatrizz[28][161] = 9'b111111111;
assign micromatrizz[28][162] = 9'b111111111;
assign micromatrizz[28][163] = 9'b111111111;
assign micromatrizz[28][164] = 9'b111111111;
assign micromatrizz[28][165] = 9'b111111111;
assign micromatrizz[28][166] = 9'b111111111;
assign micromatrizz[28][167] = 9'b111111111;
assign micromatrizz[28][168] = 9'b111111111;
assign micromatrizz[28][169] = 9'b111111111;
assign micromatrizz[28][170] = 9'b111111111;
assign micromatrizz[28][171] = 9'b111111111;
assign micromatrizz[28][172] = 9'b111111111;
assign micromatrizz[28][173] = 9'b111111111;
assign micromatrizz[28][174] = 9'b111111111;
assign micromatrizz[28][175] = 9'b111111111;
assign micromatrizz[28][176] = 9'b111111111;
assign micromatrizz[28][177] = 9'b111111111;
assign micromatrizz[28][178] = 9'b111111111;
assign micromatrizz[28][179] = 9'b111111111;
assign micromatrizz[28][180] = 9'b111111111;
assign micromatrizz[28][181] = 9'b111111111;
assign micromatrizz[28][182] = 9'b111111111;
assign micromatrizz[28][183] = 9'b111111111;
assign micromatrizz[28][184] = 9'b111111111;
assign micromatrizz[28][185] = 9'b111111111;
assign micromatrizz[28][186] = 9'b111111111;
assign micromatrizz[28][187] = 9'b111111111;
assign micromatrizz[28][188] = 9'b111111111;
assign micromatrizz[28][189] = 9'b111111111;
assign micromatrizz[28][190] = 9'b111111111;
assign micromatrizz[28][191] = 9'b111111111;
assign micromatrizz[28][192] = 9'b111111111;
assign micromatrizz[28][193] = 9'b111111111;
assign micromatrizz[28][194] = 9'b111111111;
assign micromatrizz[28][195] = 9'b111111111;
assign micromatrizz[28][196] = 9'b111111111;
assign micromatrizz[28][197] = 9'b111111111;
assign micromatrizz[28][198] = 9'b111111111;
assign micromatrizz[28][199] = 9'b111111111;
assign micromatrizz[28][200] = 9'b111111111;
assign micromatrizz[28][201] = 9'b111111111;
assign micromatrizz[28][202] = 9'b111111111;
assign micromatrizz[28][203] = 9'b111111111;
assign micromatrizz[28][204] = 9'b111111111;
assign micromatrizz[28][205] = 9'b111111111;
assign micromatrizz[28][206] = 9'b111111111;
assign micromatrizz[28][207] = 9'b111111111;
assign micromatrizz[28][208] = 9'b111111111;
assign micromatrizz[28][209] = 9'b111111111;
assign micromatrizz[28][210] = 9'b111111111;
assign micromatrizz[28][211] = 9'b111111111;
assign micromatrizz[28][212] = 9'b111111111;
assign micromatrizz[28][213] = 9'b111111111;
assign micromatrizz[28][214] = 9'b111111111;
assign micromatrizz[28][215] = 9'b111111111;
assign micromatrizz[28][216] = 9'b111111111;
assign micromatrizz[28][217] = 9'b111111111;
assign micromatrizz[28][218] = 9'b111111111;
assign micromatrizz[28][219] = 9'b111111111;
assign micromatrizz[28][220] = 9'b111111111;
assign micromatrizz[28][221] = 9'b111111111;
assign micromatrizz[28][222] = 9'b111111111;
assign micromatrizz[28][223] = 9'b111111111;
assign micromatrizz[28][224] = 9'b111111111;
assign micromatrizz[28][225] = 9'b111111111;
assign micromatrizz[28][226] = 9'b111111111;
assign micromatrizz[28][227] = 9'b111111111;
assign micromatrizz[28][228] = 9'b111111111;
assign micromatrizz[28][229] = 9'b111111111;
assign micromatrizz[28][230] = 9'b111111111;
assign micromatrizz[28][231] = 9'b111111111;
assign micromatrizz[28][232] = 9'b111111111;
assign micromatrizz[28][233] = 9'b111111111;
assign micromatrizz[28][234] = 9'b111111111;
assign micromatrizz[28][235] = 9'b111111111;
assign micromatrizz[28][236] = 9'b111111111;
assign micromatrizz[28][237] = 9'b111111111;
assign micromatrizz[28][238] = 9'b111111111;
assign micromatrizz[28][239] = 9'b111111111;
assign micromatrizz[28][240] = 9'b111111111;
assign micromatrizz[28][241] = 9'b111111111;
assign micromatrizz[28][242] = 9'b111111111;
assign micromatrizz[28][243] = 9'b111111111;
assign micromatrizz[28][244] = 9'b111111111;
assign micromatrizz[28][245] = 9'b111111111;
assign micromatrizz[28][246] = 9'b111111111;
assign micromatrizz[28][247] = 9'b111111111;
assign micromatrizz[28][248] = 9'b111111111;
assign micromatrizz[28][249] = 9'b111111111;
assign micromatrizz[28][250] = 9'b111111111;
assign micromatrizz[28][251] = 9'b111111111;
assign micromatrizz[28][252] = 9'b111111111;
assign micromatrizz[28][253] = 9'b111111111;
assign micromatrizz[28][254] = 9'b111111111;
assign micromatrizz[28][255] = 9'b111111111;
assign micromatrizz[28][256] = 9'b111111111;
assign micromatrizz[28][257] = 9'b111111111;
assign micromatrizz[28][258] = 9'b111111111;
assign micromatrizz[28][259] = 9'b111111111;
assign micromatrizz[28][260] = 9'b111111111;
assign micromatrizz[28][261] = 9'b111111111;
assign micromatrizz[28][262] = 9'b111111111;
assign micromatrizz[28][263] = 9'b111111111;
assign micromatrizz[28][264] = 9'b111111111;
assign micromatrizz[28][265] = 9'b111111111;
assign micromatrizz[28][266] = 9'b111111111;
assign micromatrizz[28][267] = 9'b111111111;
assign micromatrizz[28][268] = 9'b111111111;
assign micromatrizz[28][269] = 9'b111111111;
assign micromatrizz[28][270] = 9'b111110010;
assign micromatrizz[28][271] = 9'b111110010;
assign micromatrizz[28][272] = 9'b111110010;
assign micromatrizz[28][273] = 9'b111110010;
assign micromatrizz[28][274] = 9'b111110011;
assign micromatrizz[28][275] = 9'b111110011;
assign micromatrizz[28][276] = 9'b111110011;
assign micromatrizz[28][277] = 9'b111110011;
assign micromatrizz[28][278] = 9'b111110011;
assign micromatrizz[28][279] = 9'b111111111;
assign micromatrizz[28][280] = 9'b111111111;
assign micromatrizz[28][281] = 9'b111111111;
assign micromatrizz[28][282] = 9'b111111111;
assign micromatrizz[28][283] = 9'b111111111;
assign micromatrizz[28][284] = 9'b111111111;
assign micromatrizz[28][285] = 9'b111111111;
assign micromatrizz[28][286] = 9'b111111111;
assign micromatrizz[28][287] = 9'b111111111;
assign micromatrizz[28][288] = 9'b111111111;
assign micromatrizz[28][289] = 9'b111111111;
assign micromatrizz[28][290] = 9'b111110010;
assign micromatrizz[28][291] = 9'b111110010;
assign micromatrizz[28][292] = 9'b111110010;
assign micromatrizz[28][293] = 9'b111110011;
assign micromatrizz[28][294] = 9'b111110011;
assign micromatrizz[28][295] = 9'b111110011;
assign micromatrizz[28][296] = 9'b111110011;
assign micromatrizz[28][297] = 9'b111110111;
assign micromatrizz[28][298] = 9'b111111111;
assign micromatrizz[28][299] = 9'b111111111;
assign micromatrizz[28][300] = 9'b111111111;
assign micromatrizz[28][301] = 9'b111111111;
assign micromatrizz[28][302] = 9'b111111111;
assign micromatrizz[28][303] = 9'b111111111;
assign micromatrizz[28][304] = 9'b111111111;
assign micromatrizz[28][305] = 9'b111110010;
assign micromatrizz[28][306] = 9'b111111111;
assign micromatrizz[28][307] = 9'b111111111;
assign micromatrizz[28][308] = 9'b111111111;
assign micromatrizz[28][309] = 9'b111110010;
assign micromatrizz[28][310] = 9'b111110010;
assign micromatrizz[28][311] = 9'b111110011;
assign micromatrizz[28][312] = 9'b111110010;
assign micromatrizz[28][313] = 9'b111110010;
assign micromatrizz[28][314] = 9'b111110011;
assign micromatrizz[28][315] = 9'b111110011;
assign micromatrizz[28][316] = 9'b111110011;
assign micromatrizz[28][317] = 9'b111110010;
assign micromatrizz[28][318] = 9'b111111111;
assign micromatrizz[28][319] = 9'b111111111;
assign micromatrizz[28][320] = 9'b111111111;
assign micromatrizz[28][321] = 9'b111111111;
assign micromatrizz[28][322] = 9'b111111111;
assign micromatrizz[28][323] = 9'b111111111;
assign micromatrizz[28][324] = 9'b111111111;
assign micromatrizz[28][325] = 9'b111111111;
assign micromatrizz[28][326] = 9'b111111111;
assign micromatrizz[28][327] = 9'b111111111;
assign micromatrizz[28][328] = 9'b111111111;
assign micromatrizz[28][329] = 9'b111111111;
assign micromatrizz[28][330] = 9'b111111111;
assign micromatrizz[28][331] = 9'b111111111;
assign micromatrizz[28][332] = 9'b111111111;
assign micromatrizz[28][333] = 9'b111111111;
assign micromatrizz[28][334] = 9'b111111111;
assign micromatrizz[28][335] = 9'b111111111;
assign micromatrizz[28][336] = 9'b111111111;
assign micromatrizz[28][337] = 9'b111111111;
assign micromatrizz[28][338] = 9'b111111111;
assign micromatrizz[28][339] = 9'b111111111;
assign micromatrizz[28][340] = 9'b111111111;
assign micromatrizz[28][341] = 9'b111111111;
assign micromatrizz[28][342] = 9'b111111111;
assign micromatrizz[28][343] = 9'b111111111;
assign micromatrizz[28][344] = 9'b111111111;
assign micromatrizz[28][345] = 9'b111111111;
assign micromatrizz[28][346] = 9'b111111111;
assign micromatrizz[28][347] = 9'b111111111;
assign micromatrizz[28][348] = 9'b111111111;
assign micromatrizz[28][349] = 9'b111111111;
assign micromatrizz[28][350] = 9'b111111111;
assign micromatrizz[28][351] = 9'b111111111;
assign micromatrizz[28][352] = 9'b111111111;
assign micromatrizz[28][353] = 9'b111111111;
assign micromatrizz[28][354] = 9'b111111111;
assign micromatrizz[28][355] = 9'b111111111;
assign micromatrizz[28][356] = 9'b111111111;
assign micromatrizz[28][357] = 9'b111111111;
assign micromatrizz[28][358] = 9'b111111111;
assign micromatrizz[28][359] = 9'b111111111;
assign micromatrizz[28][360] = 9'b111111111;
assign micromatrizz[28][361] = 9'b111111111;
assign micromatrizz[28][362] = 9'b111111111;
assign micromatrizz[28][363] = 9'b111111111;
assign micromatrizz[28][364] = 9'b111111111;
assign micromatrizz[28][365] = 9'b111111111;
assign micromatrizz[28][366] = 9'b111111111;
assign micromatrizz[28][367] = 9'b111111111;
assign micromatrizz[28][368] = 9'b111111111;
assign micromatrizz[28][369] = 9'b111111111;
assign micromatrizz[28][370] = 9'b111111111;
assign micromatrizz[28][371] = 9'b111111111;
assign micromatrizz[28][372] = 9'b111111111;
assign micromatrizz[28][373] = 9'b111111111;
assign micromatrizz[28][374] = 9'b111111111;
assign micromatrizz[28][375] = 9'b111111111;
assign micromatrizz[28][376] = 9'b111111111;
assign micromatrizz[28][377] = 9'b111111111;
assign micromatrizz[28][378] = 9'b111111111;
assign micromatrizz[28][379] = 9'b111111111;
assign micromatrizz[28][380] = 9'b111111111;
assign micromatrizz[28][381] = 9'b111111111;
assign micromatrizz[28][382] = 9'b111111111;
assign micromatrizz[28][383] = 9'b111111111;
assign micromatrizz[28][384] = 9'b111111111;
assign micromatrizz[28][385] = 9'b111111111;
assign micromatrizz[28][386] = 9'b111111111;
assign micromatrizz[28][387] = 9'b111111111;
assign micromatrizz[28][388] = 9'b111111111;
assign micromatrizz[28][389] = 9'b111111111;
assign micromatrizz[28][390] = 9'b111111111;
assign micromatrizz[28][391] = 9'b111111111;
assign micromatrizz[28][392] = 9'b111111111;
assign micromatrizz[28][393] = 9'b111111111;
assign micromatrizz[28][394] = 9'b111111111;
assign micromatrizz[28][395] = 9'b111111111;
assign micromatrizz[28][396] = 9'b111111111;
assign micromatrizz[28][397] = 9'b111111111;
assign micromatrizz[28][398] = 9'b111111111;
assign micromatrizz[28][399] = 9'b111111111;
assign micromatrizz[28][400] = 9'b111111111;
assign micromatrizz[28][401] = 9'b111111111;
assign micromatrizz[28][402] = 9'b111111111;
assign micromatrizz[28][403] = 9'b111111111;
assign micromatrizz[28][404] = 9'b111111111;
assign micromatrizz[28][405] = 9'b111111111;
assign micromatrizz[28][406] = 9'b111111111;
assign micromatrizz[28][407] = 9'b111111111;
assign micromatrizz[28][408] = 9'b111111111;
assign micromatrizz[28][409] = 9'b111111111;
assign micromatrizz[28][410] = 9'b111111111;
assign micromatrizz[28][411] = 9'b111111111;
assign micromatrizz[28][412] = 9'b111111111;
assign micromatrizz[28][413] = 9'b111111111;
assign micromatrizz[28][414] = 9'b111111111;
assign micromatrizz[28][415] = 9'b111111111;
assign micromatrizz[28][416] = 9'b111111111;
assign micromatrizz[28][417] = 9'b111111111;
assign micromatrizz[28][418] = 9'b111111111;
assign micromatrizz[28][419] = 9'b111111111;
assign micromatrizz[28][420] = 9'b111111111;
assign micromatrizz[28][421] = 9'b111111111;
assign micromatrizz[28][422] = 9'b111111111;
assign micromatrizz[28][423] = 9'b111111111;
assign micromatrizz[28][424] = 9'b111111111;
assign micromatrizz[28][425] = 9'b111111111;
assign micromatrizz[28][426] = 9'b111111111;
assign micromatrizz[28][427] = 9'b111111111;
assign micromatrizz[28][428] = 9'b111111111;
assign micromatrizz[28][429] = 9'b111111111;
assign micromatrizz[28][430] = 9'b111111111;
assign micromatrizz[28][431] = 9'b111111111;
assign micromatrizz[28][432] = 9'b111111111;
assign micromatrizz[28][433] = 9'b111111111;
assign micromatrizz[28][434] = 9'b111111111;
assign micromatrizz[28][435] = 9'b111111111;
assign micromatrizz[28][436] = 9'b111111111;
assign micromatrizz[28][437] = 9'b111111111;
assign micromatrizz[28][438] = 9'b111111111;
assign micromatrizz[28][439] = 9'b111111111;
assign micromatrizz[28][440] = 9'b111111111;
assign micromatrizz[28][441] = 9'b111111111;
assign micromatrizz[28][442] = 9'b111111111;
assign micromatrizz[28][443] = 9'b111111111;
assign micromatrizz[28][444] = 9'b111111111;
assign micromatrizz[28][445] = 9'b111111111;
assign micromatrizz[28][446] = 9'b111111111;
assign micromatrizz[28][447] = 9'b111111111;
assign micromatrizz[28][448] = 9'b111111111;
assign micromatrizz[28][449] = 9'b111111111;
assign micromatrizz[28][450] = 9'b111111111;
assign micromatrizz[28][451] = 9'b111111111;
assign micromatrizz[28][452] = 9'b111111111;
assign micromatrizz[28][453] = 9'b111111111;
assign micromatrizz[28][454] = 9'b111111111;
assign micromatrizz[28][455] = 9'b111111111;
assign micromatrizz[28][456] = 9'b111111111;
assign micromatrizz[28][457] = 9'b111111111;
assign micromatrizz[28][458] = 9'b111111111;
assign micromatrizz[28][459] = 9'b111111111;
assign micromatrizz[28][460] = 9'b111111111;
assign micromatrizz[28][461] = 9'b111111111;
assign micromatrizz[28][462] = 9'b111111111;
assign micromatrizz[28][463] = 9'b111111111;
assign micromatrizz[28][464] = 9'b111111111;
assign micromatrizz[28][465] = 9'b111111111;
assign micromatrizz[28][466] = 9'b111111111;
assign micromatrizz[28][467] = 9'b111111111;
assign micromatrizz[28][468] = 9'b111111111;
assign micromatrizz[28][469] = 9'b111111111;
assign micromatrizz[28][470] = 9'b111111111;
assign micromatrizz[28][471] = 9'b111111111;
assign micromatrizz[28][472] = 9'b111111111;
assign micromatrizz[28][473] = 9'b111111111;
assign micromatrizz[28][474] = 9'b111111111;
assign micromatrizz[28][475] = 9'b111111111;
assign micromatrizz[28][476] = 9'b111111111;
assign micromatrizz[28][477] = 9'b111111111;
assign micromatrizz[28][478] = 9'b111111111;
assign micromatrizz[28][479] = 9'b111111111;
assign micromatrizz[28][480] = 9'b111111111;
assign micromatrizz[28][481] = 9'b111111111;
assign micromatrizz[28][482] = 9'b111111111;
assign micromatrizz[28][483] = 9'b111111111;
assign micromatrizz[28][484] = 9'b111111111;
assign micromatrizz[28][485] = 9'b111111111;
assign micromatrizz[28][486] = 9'b111111111;
assign micromatrizz[28][487] = 9'b111111111;
assign micromatrizz[28][488] = 9'b111111111;
assign micromatrizz[28][489] = 9'b111111111;
assign micromatrizz[28][490] = 9'b111111111;
assign micromatrizz[28][491] = 9'b111111111;
assign micromatrizz[28][492] = 9'b111111111;
assign micromatrizz[28][493] = 9'b111111111;
assign micromatrizz[28][494] = 9'b111111111;
assign micromatrizz[28][495] = 9'b111111111;
assign micromatrizz[28][496] = 9'b111111111;
assign micromatrizz[28][497] = 9'b111111111;
assign micromatrizz[28][498] = 9'b111111111;
assign micromatrizz[28][499] = 9'b111111111;
assign micromatrizz[28][500] = 9'b111111111;
assign micromatrizz[28][501] = 9'b111111111;
assign micromatrizz[28][502] = 9'b111111111;
assign micromatrizz[28][503] = 9'b111111111;
assign micromatrizz[28][504] = 9'b111111111;
assign micromatrizz[28][505] = 9'b111111111;
assign micromatrizz[28][506] = 9'b111111111;
assign micromatrizz[28][507] = 9'b111111111;
assign micromatrizz[28][508] = 9'b111111111;
assign micromatrizz[28][509] = 9'b111111111;
assign micromatrizz[28][510] = 9'b111111111;
assign micromatrizz[28][511] = 9'b111111111;
assign micromatrizz[28][512] = 9'b111111111;
assign micromatrizz[28][513] = 9'b111111111;
assign micromatrizz[28][514] = 9'b111111111;
assign micromatrizz[28][515] = 9'b111111111;
assign micromatrizz[28][516] = 9'b111111111;
assign micromatrizz[28][517] = 9'b111111111;
assign micromatrizz[28][518] = 9'b111111111;
assign micromatrizz[28][519] = 9'b111111111;
assign micromatrizz[28][520] = 9'b111111111;
assign micromatrizz[28][521] = 9'b111111111;
assign micromatrizz[28][522] = 9'b111111111;
assign micromatrizz[28][523] = 9'b111111111;
assign micromatrizz[28][524] = 9'b111111111;
assign micromatrizz[28][525] = 9'b111111111;
assign micromatrizz[28][526] = 9'b111111111;
assign micromatrizz[28][527] = 9'b111111111;
assign micromatrizz[28][528] = 9'b111111111;
assign micromatrizz[28][529] = 9'b111111111;
assign micromatrizz[28][530] = 9'b111111111;
assign micromatrizz[28][531] = 9'b111111111;
assign micromatrizz[28][532] = 9'b111111111;
assign micromatrizz[28][533] = 9'b111111111;
assign micromatrizz[28][534] = 9'b111111111;
assign micromatrizz[28][535] = 9'b111111111;
assign micromatrizz[28][536] = 9'b111111111;
assign micromatrizz[28][537] = 9'b111111111;
assign micromatrizz[28][538] = 9'b111111111;
assign micromatrizz[28][539] = 9'b111111111;
assign micromatrizz[28][540] = 9'b111111111;
assign micromatrizz[28][541] = 9'b111111111;
assign micromatrizz[28][542] = 9'b111111111;
assign micromatrizz[28][543] = 9'b111111111;
assign micromatrizz[28][544] = 9'b111111111;
assign micromatrizz[28][545] = 9'b111111111;
assign micromatrizz[28][546] = 9'b111111111;
assign micromatrizz[28][547] = 9'b111111111;
assign micromatrizz[28][548] = 9'b111111111;
assign micromatrizz[28][549] = 9'b111111111;
assign micromatrizz[28][550] = 9'b111111111;
assign micromatrizz[28][551] = 9'b111111111;
assign micromatrizz[28][552] = 9'b111111111;
assign micromatrizz[28][553] = 9'b111111111;
assign micromatrizz[28][554] = 9'b111111111;
assign micromatrizz[28][555] = 9'b111111111;
assign micromatrizz[28][556] = 9'b111111111;
assign micromatrizz[28][557] = 9'b111111111;
assign micromatrizz[28][558] = 9'b111111111;
assign micromatrizz[28][559] = 9'b111111111;
assign micromatrizz[28][560] = 9'b111111111;
assign micromatrizz[28][561] = 9'b111111111;
assign micromatrizz[28][562] = 9'b111111111;
assign micromatrizz[28][563] = 9'b111111111;
assign micromatrizz[28][564] = 9'b111111111;
assign micromatrizz[28][565] = 9'b111111111;
assign micromatrizz[28][566] = 9'b111111111;
assign micromatrizz[28][567] = 9'b111111111;
assign micromatrizz[28][568] = 9'b111111111;
assign micromatrizz[28][569] = 9'b111111111;
assign micromatrizz[28][570] = 9'b111111111;
assign micromatrizz[28][571] = 9'b111111111;
assign micromatrizz[28][572] = 9'b111111111;
assign micromatrizz[28][573] = 9'b111111111;
assign micromatrizz[28][574] = 9'b111111111;
assign micromatrizz[28][575] = 9'b111111111;
assign micromatrizz[28][576] = 9'b111111111;
assign micromatrizz[28][577] = 9'b111111111;
assign micromatrizz[28][578] = 9'b111111111;
assign micromatrizz[28][579] = 9'b111111111;
assign micromatrizz[28][580] = 9'b111111111;
assign micromatrizz[28][581] = 9'b111111111;
assign micromatrizz[28][582] = 9'b111111111;
assign micromatrizz[28][583] = 9'b111111111;
assign micromatrizz[28][584] = 9'b111111111;
assign micromatrizz[28][585] = 9'b111111111;
assign micromatrizz[28][586] = 9'b111111111;
assign micromatrizz[28][587] = 9'b111111111;
assign micromatrizz[28][588] = 9'b111111111;
assign micromatrizz[28][589] = 9'b111111111;
assign micromatrizz[28][590] = 9'b111111111;
assign micromatrizz[28][591] = 9'b111111111;
assign micromatrizz[28][592] = 9'b111111111;
assign micromatrizz[28][593] = 9'b111111111;
assign micromatrizz[28][594] = 9'b111111111;
assign micromatrizz[28][595] = 9'b111111111;
assign micromatrizz[28][596] = 9'b111111111;
assign micromatrizz[28][597] = 9'b111111111;
assign micromatrizz[28][598] = 9'b111111111;
assign micromatrizz[28][599] = 9'b111111111;
assign micromatrizz[28][600] = 9'b111111111;
assign micromatrizz[28][601] = 9'b111111111;
assign micromatrizz[28][602] = 9'b111111111;
assign micromatrizz[28][603] = 9'b111111111;
assign micromatrizz[28][604] = 9'b111111111;
assign micromatrizz[28][605] = 9'b111111111;
assign micromatrizz[28][606] = 9'b111111111;
assign micromatrizz[28][607] = 9'b111111111;
assign micromatrizz[28][608] = 9'b111111111;
assign micromatrizz[28][609] = 9'b111111111;
assign micromatrizz[28][610] = 9'b111111111;
assign micromatrizz[28][611] = 9'b111111111;
assign micromatrizz[28][612] = 9'b111111111;
assign micromatrizz[28][613] = 9'b111111111;
assign micromatrizz[28][614] = 9'b111111111;
assign micromatrizz[28][615] = 9'b111111111;
assign micromatrizz[28][616] = 9'b111111111;
assign micromatrizz[28][617] = 9'b111111111;
assign micromatrizz[28][618] = 9'b111111111;
assign micromatrizz[28][619] = 9'b111111111;
assign micromatrizz[28][620] = 9'b111111111;
assign micromatrizz[28][621] = 9'b111111111;
assign micromatrizz[28][622] = 9'b111111111;
assign micromatrizz[28][623] = 9'b111111111;
assign micromatrizz[28][624] = 9'b111111111;
assign micromatrizz[28][625] = 9'b111111111;
assign micromatrizz[28][626] = 9'b111111111;
assign micromatrizz[28][627] = 9'b111111111;
assign micromatrizz[28][628] = 9'b111111111;
assign micromatrizz[28][629] = 9'b111111111;
assign micromatrizz[28][630] = 9'b111111111;
assign micromatrizz[28][631] = 9'b111111111;
assign micromatrizz[28][632] = 9'b111111111;
assign micromatrizz[28][633] = 9'b111111111;
assign micromatrizz[28][634] = 9'b111111111;
assign micromatrizz[28][635] = 9'b111111111;
assign micromatrizz[28][636] = 9'b111111111;
assign micromatrizz[28][637] = 9'b111111111;
assign micromatrizz[28][638] = 9'b111111111;
assign micromatrizz[28][639] = 9'b111111111;
assign micromatrizz[29][0] = 9'b111111111;
assign micromatrizz[29][1] = 9'b111111111;
assign micromatrizz[29][2] = 9'b111111111;
assign micromatrizz[29][3] = 9'b111111111;
assign micromatrizz[29][4] = 9'b111111111;
assign micromatrizz[29][5] = 9'b111111111;
assign micromatrizz[29][6] = 9'b111111111;
assign micromatrizz[29][7] = 9'b111111111;
assign micromatrizz[29][8] = 9'b111111111;
assign micromatrizz[29][9] = 9'b111111111;
assign micromatrizz[29][10] = 9'b111111111;
assign micromatrizz[29][11] = 9'b111111111;
assign micromatrizz[29][12] = 9'b111111111;
assign micromatrizz[29][13] = 9'b111111111;
assign micromatrizz[29][14] = 9'b111111111;
assign micromatrizz[29][15] = 9'b111111111;
assign micromatrizz[29][16] = 9'b111111111;
assign micromatrizz[29][17] = 9'b111111111;
assign micromatrizz[29][18] = 9'b111111111;
assign micromatrizz[29][19] = 9'b111111111;
assign micromatrizz[29][20] = 9'b111111111;
assign micromatrizz[29][21] = 9'b111111111;
assign micromatrizz[29][22] = 9'b111111111;
assign micromatrizz[29][23] = 9'b111111111;
assign micromatrizz[29][24] = 9'b111111111;
assign micromatrizz[29][25] = 9'b111111111;
assign micromatrizz[29][26] = 9'b111111111;
assign micromatrizz[29][27] = 9'b111111111;
assign micromatrizz[29][28] = 9'b111111111;
assign micromatrizz[29][29] = 9'b111111111;
assign micromatrizz[29][30] = 9'b111111111;
assign micromatrizz[29][31] = 9'b111111111;
assign micromatrizz[29][32] = 9'b111111111;
assign micromatrizz[29][33] = 9'b111111111;
assign micromatrizz[29][34] = 9'b111111111;
assign micromatrizz[29][35] = 9'b111111111;
assign micromatrizz[29][36] = 9'b111111111;
assign micromatrizz[29][37] = 9'b111111111;
assign micromatrizz[29][38] = 9'b111111111;
assign micromatrizz[29][39] = 9'b111111111;
assign micromatrizz[29][40] = 9'b111111111;
assign micromatrizz[29][41] = 9'b111111111;
assign micromatrizz[29][42] = 9'b111111111;
assign micromatrizz[29][43] = 9'b111111111;
assign micromatrizz[29][44] = 9'b111111111;
assign micromatrizz[29][45] = 9'b111111111;
assign micromatrizz[29][46] = 9'b111111111;
assign micromatrizz[29][47] = 9'b111111111;
assign micromatrizz[29][48] = 9'b111111111;
assign micromatrizz[29][49] = 9'b111111111;
assign micromatrizz[29][50] = 9'b111111111;
assign micromatrizz[29][51] = 9'b111111111;
assign micromatrizz[29][52] = 9'b111111111;
assign micromatrizz[29][53] = 9'b111111111;
assign micromatrizz[29][54] = 9'b111111111;
assign micromatrizz[29][55] = 9'b111111111;
assign micromatrizz[29][56] = 9'b111111111;
assign micromatrizz[29][57] = 9'b111111111;
assign micromatrizz[29][58] = 9'b111111111;
assign micromatrizz[29][59] = 9'b111111111;
assign micromatrizz[29][60] = 9'b111111111;
assign micromatrizz[29][61] = 9'b111111111;
assign micromatrizz[29][62] = 9'b111111111;
assign micromatrizz[29][63] = 9'b111111111;
assign micromatrizz[29][64] = 9'b111111111;
assign micromatrizz[29][65] = 9'b111111111;
assign micromatrizz[29][66] = 9'b111111111;
assign micromatrizz[29][67] = 9'b111111111;
assign micromatrizz[29][68] = 9'b111111111;
assign micromatrizz[29][69] = 9'b111111111;
assign micromatrizz[29][70] = 9'b111111111;
assign micromatrizz[29][71] = 9'b111111111;
assign micromatrizz[29][72] = 9'b111111111;
assign micromatrizz[29][73] = 9'b111111111;
assign micromatrizz[29][74] = 9'b111111111;
assign micromatrizz[29][75] = 9'b111111111;
assign micromatrizz[29][76] = 9'b111111111;
assign micromatrizz[29][77] = 9'b111111111;
assign micromatrizz[29][78] = 9'b111111111;
assign micromatrizz[29][79] = 9'b111111111;
assign micromatrizz[29][80] = 9'b111111111;
assign micromatrizz[29][81] = 9'b111111111;
assign micromatrizz[29][82] = 9'b111111111;
assign micromatrizz[29][83] = 9'b111111111;
assign micromatrizz[29][84] = 9'b111111111;
assign micromatrizz[29][85] = 9'b111111111;
assign micromatrizz[29][86] = 9'b111111111;
assign micromatrizz[29][87] = 9'b111111111;
assign micromatrizz[29][88] = 9'b111111111;
assign micromatrizz[29][89] = 9'b111111111;
assign micromatrizz[29][90] = 9'b111111111;
assign micromatrizz[29][91] = 9'b111111111;
assign micromatrizz[29][92] = 9'b111111111;
assign micromatrizz[29][93] = 9'b111111111;
assign micromatrizz[29][94] = 9'b111111111;
assign micromatrizz[29][95] = 9'b111111111;
assign micromatrizz[29][96] = 9'b111111111;
assign micromatrizz[29][97] = 9'b111111111;
assign micromatrizz[29][98] = 9'b111111111;
assign micromatrizz[29][99] = 9'b111111111;
assign micromatrizz[29][100] = 9'b111111111;
assign micromatrizz[29][101] = 9'b111111111;
assign micromatrizz[29][102] = 9'b111111111;
assign micromatrizz[29][103] = 9'b111111111;
assign micromatrizz[29][104] = 9'b111111111;
assign micromatrizz[29][105] = 9'b111111111;
assign micromatrizz[29][106] = 9'b111111111;
assign micromatrizz[29][107] = 9'b111111111;
assign micromatrizz[29][108] = 9'b111111111;
assign micromatrizz[29][109] = 9'b111111111;
assign micromatrizz[29][110] = 9'b111111111;
assign micromatrizz[29][111] = 9'b111111111;
assign micromatrizz[29][112] = 9'b111111111;
assign micromatrizz[29][113] = 9'b111111111;
assign micromatrizz[29][114] = 9'b111111111;
assign micromatrizz[29][115] = 9'b111111111;
assign micromatrizz[29][116] = 9'b111111111;
assign micromatrizz[29][117] = 9'b111111111;
assign micromatrizz[29][118] = 9'b111111111;
assign micromatrizz[29][119] = 9'b111111111;
assign micromatrizz[29][120] = 9'b111111111;
assign micromatrizz[29][121] = 9'b111111111;
assign micromatrizz[29][122] = 9'b111111111;
assign micromatrizz[29][123] = 9'b111111111;
assign micromatrizz[29][124] = 9'b111111111;
assign micromatrizz[29][125] = 9'b111111111;
assign micromatrizz[29][126] = 9'b111111111;
assign micromatrizz[29][127] = 9'b111111111;
assign micromatrizz[29][128] = 9'b111111111;
assign micromatrizz[29][129] = 9'b111111111;
assign micromatrizz[29][130] = 9'b111111111;
assign micromatrizz[29][131] = 9'b111111111;
assign micromatrizz[29][132] = 9'b111111111;
assign micromatrizz[29][133] = 9'b111111111;
assign micromatrizz[29][134] = 9'b111111111;
assign micromatrizz[29][135] = 9'b111111111;
assign micromatrizz[29][136] = 9'b111111111;
assign micromatrizz[29][137] = 9'b111111111;
assign micromatrizz[29][138] = 9'b111111111;
assign micromatrizz[29][139] = 9'b111111111;
assign micromatrizz[29][140] = 9'b111111111;
assign micromatrizz[29][141] = 9'b111111111;
assign micromatrizz[29][142] = 9'b111111111;
assign micromatrizz[29][143] = 9'b111111111;
assign micromatrizz[29][144] = 9'b111111111;
assign micromatrizz[29][145] = 9'b111111111;
assign micromatrizz[29][146] = 9'b111111111;
assign micromatrizz[29][147] = 9'b111111111;
assign micromatrizz[29][148] = 9'b111111111;
assign micromatrizz[29][149] = 9'b111111111;
assign micromatrizz[29][150] = 9'b111111111;
assign micromatrizz[29][151] = 9'b111111111;
assign micromatrizz[29][152] = 9'b111111111;
assign micromatrizz[29][153] = 9'b111111111;
assign micromatrizz[29][154] = 9'b111111111;
assign micromatrizz[29][155] = 9'b111111111;
assign micromatrizz[29][156] = 9'b111111111;
assign micromatrizz[29][157] = 9'b111111111;
assign micromatrizz[29][158] = 9'b111111111;
assign micromatrizz[29][159] = 9'b111111111;
assign micromatrizz[29][160] = 9'b111111111;
assign micromatrizz[29][161] = 9'b111111111;
assign micromatrizz[29][162] = 9'b111111111;
assign micromatrizz[29][163] = 9'b111111111;
assign micromatrizz[29][164] = 9'b111111111;
assign micromatrizz[29][165] = 9'b111111111;
assign micromatrizz[29][166] = 9'b111111111;
assign micromatrizz[29][167] = 9'b111111111;
assign micromatrizz[29][168] = 9'b111111111;
assign micromatrizz[29][169] = 9'b111111111;
assign micromatrizz[29][170] = 9'b111111111;
assign micromatrizz[29][171] = 9'b111111111;
assign micromatrizz[29][172] = 9'b111111111;
assign micromatrizz[29][173] = 9'b111111111;
assign micromatrizz[29][174] = 9'b111111111;
assign micromatrizz[29][175] = 9'b111111111;
assign micromatrizz[29][176] = 9'b111111111;
assign micromatrizz[29][177] = 9'b111111111;
assign micromatrizz[29][178] = 9'b111111111;
assign micromatrizz[29][179] = 9'b111111111;
assign micromatrizz[29][180] = 9'b111111111;
assign micromatrizz[29][181] = 9'b111111111;
assign micromatrizz[29][182] = 9'b111111111;
assign micromatrizz[29][183] = 9'b111111111;
assign micromatrizz[29][184] = 9'b111111111;
assign micromatrizz[29][185] = 9'b111111111;
assign micromatrizz[29][186] = 9'b111111111;
assign micromatrizz[29][187] = 9'b111111111;
assign micromatrizz[29][188] = 9'b111111111;
assign micromatrizz[29][189] = 9'b111111111;
assign micromatrizz[29][190] = 9'b111111111;
assign micromatrizz[29][191] = 9'b111111111;
assign micromatrizz[29][192] = 9'b111111111;
assign micromatrizz[29][193] = 9'b111111111;
assign micromatrizz[29][194] = 9'b111111111;
assign micromatrizz[29][195] = 9'b111111111;
assign micromatrizz[29][196] = 9'b111111111;
assign micromatrizz[29][197] = 9'b111111111;
assign micromatrizz[29][198] = 9'b111111111;
assign micromatrizz[29][199] = 9'b111111111;
assign micromatrizz[29][200] = 9'b111111111;
assign micromatrizz[29][201] = 9'b111111111;
assign micromatrizz[29][202] = 9'b111111111;
assign micromatrizz[29][203] = 9'b111111111;
assign micromatrizz[29][204] = 9'b111111111;
assign micromatrizz[29][205] = 9'b111111111;
assign micromatrizz[29][206] = 9'b111111111;
assign micromatrizz[29][207] = 9'b111111111;
assign micromatrizz[29][208] = 9'b111111111;
assign micromatrizz[29][209] = 9'b111111111;
assign micromatrizz[29][210] = 9'b111111111;
assign micromatrizz[29][211] = 9'b111111111;
assign micromatrizz[29][212] = 9'b111111111;
assign micromatrizz[29][213] = 9'b111111111;
assign micromatrizz[29][214] = 9'b111111111;
assign micromatrizz[29][215] = 9'b111111111;
assign micromatrizz[29][216] = 9'b111111111;
assign micromatrizz[29][217] = 9'b111111111;
assign micromatrizz[29][218] = 9'b111111111;
assign micromatrizz[29][219] = 9'b111111111;
assign micromatrizz[29][220] = 9'b111111111;
assign micromatrizz[29][221] = 9'b111111111;
assign micromatrizz[29][222] = 9'b111111111;
assign micromatrizz[29][223] = 9'b111111111;
assign micromatrizz[29][224] = 9'b111111111;
assign micromatrizz[29][225] = 9'b111111111;
assign micromatrizz[29][226] = 9'b111111111;
assign micromatrizz[29][227] = 9'b111111111;
assign micromatrizz[29][228] = 9'b111111111;
assign micromatrizz[29][229] = 9'b111111111;
assign micromatrizz[29][230] = 9'b111111111;
assign micromatrizz[29][231] = 9'b111111111;
assign micromatrizz[29][232] = 9'b111111111;
assign micromatrizz[29][233] = 9'b111111111;
assign micromatrizz[29][234] = 9'b111111111;
assign micromatrizz[29][235] = 9'b111111111;
assign micromatrizz[29][236] = 9'b111111111;
assign micromatrizz[29][237] = 9'b111111111;
assign micromatrizz[29][238] = 9'b111111111;
assign micromatrizz[29][239] = 9'b111111111;
assign micromatrizz[29][240] = 9'b111111111;
assign micromatrizz[29][241] = 9'b111111111;
assign micromatrizz[29][242] = 9'b111111111;
assign micromatrizz[29][243] = 9'b111111111;
assign micromatrizz[29][244] = 9'b111111111;
assign micromatrizz[29][245] = 9'b111111111;
assign micromatrizz[29][246] = 9'b111111111;
assign micromatrizz[29][247] = 9'b111111111;
assign micromatrizz[29][248] = 9'b111111111;
assign micromatrizz[29][249] = 9'b111111111;
assign micromatrizz[29][250] = 9'b111111111;
assign micromatrizz[29][251] = 9'b111111111;
assign micromatrizz[29][252] = 9'b111111111;
assign micromatrizz[29][253] = 9'b111111111;
assign micromatrizz[29][254] = 9'b111111111;
assign micromatrizz[29][255] = 9'b111111111;
assign micromatrizz[29][256] = 9'b111111111;
assign micromatrizz[29][257] = 9'b111111111;
assign micromatrizz[29][258] = 9'b111111111;
assign micromatrizz[29][259] = 9'b111111111;
assign micromatrizz[29][260] = 9'b111111111;
assign micromatrizz[29][261] = 9'b111111111;
assign micromatrizz[29][262] = 9'b111111111;
assign micromatrizz[29][263] = 9'b111111111;
assign micromatrizz[29][264] = 9'b111111111;
assign micromatrizz[29][265] = 9'b111111111;
assign micromatrizz[29][266] = 9'b111111111;
assign micromatrizz[29][267] = 9'b111111111;
assign micromatrizz[29][268] = 9'b111111111;
assign micromatrizz[29][269] = 9'b111111111;
assign micromatrizz[29][270] = 9'b111110010;
assign micromatrizz[29][271] = 9'b111110010;
assign micromatrizz[29][272] = 9'b111110010;
assign micromatrizz[29][273] = 9'b111110010;
assign micromatrizz[29][274] = 9'b111110011;
assign micromatrizz[29][275] = 9'b111110011;
assign micromatrizz[29][276] = 9'b111110011;
assign micromatrizz[29][277] = 9'b111110011;
assign micromatrizz[29][278] = 9'b111110011;
assign micromatrizz[29][279] = 9'b111111111;
assign micromatrizz[29][280] = 9'b111111111;
assign micromatrizz[29][281] = 9'b111111111;
assign micromatrizz[29][282] = 9'b111111111;
assign micromatrizz[29][283] = 9'b111111111;
assign micromatrizz[29][284] = 9'b111111111;
assign micromatrizz[29][285] = 9'b111111111;
assign micromatrizz[29][286] = 9'b111111111;
assign micromatrizz[29][287] = 9'b111111111;
assign micromatrizz[29][288] = 9'b111111111;
assign micromatrizz[29][289] = 9'b111111111;
assign micromatrizz[29][290] = 9'b111110010;
assign micromatrizz[29][291] = 9'b111110010;
assign micromatrizz[29][292] = 9'b111110011;
assign micromatrizz[29][293] = 9'b111110010;
assign micromatrizz[29][294] = 9'b111110011;
assign micromatrizz[29][295] = 9'b111110011;
assign micromatrizz[29][296] = 9'b111110011;
assign micromatrizz[29][297] = 9'b111110111;
assign micromatrizz[29][298] = 9'b111111111;
assign micromatrizz[29][299] = 9'b111111111;
assign micromatrizz[29][300] = 9'b111111111;
assign micromatrizz[29][301] = 9'b111111111;
assign micromatrizz[29][302] = 9'b111111111;
assign micromatrizz[29][303] = 9'b111111111;
assign micromatrizz[29][304] = 9'b111111111;
assign micromatrizz[29][305] = 9'b111110111;
assign micromatrizz[29][306] = 9'b111111111;
assign micromatrizz[29][307] = 9'b111111111;
assign micromatrizz[29][308] = 9'b111111111;
assign micromatrizz[29][309] = 9'b111111111;
assign micromatrizz[29][310] = 9'b111110010;
assign micromatrizz[29][311] = 9'b111110010;
assign micromatrizz[29][312] = 9'b111110010;
assign micromatrizz[29][313] = 9'b111110011;
assign micromatrizz[29][314] = 9'b111110010;
assign micromatrizz[29][315] = 9'b111110011;
assign micromatrizz[29][316] = 9'b111110011;
assign micromatrizz[29][317] = 9'b111110011;
assign micromatrizz[29][318] = 9'b111110010;
assign micromatrizz[29][319] = 9'b111110011;
assign micromatrizz[29][320] = 9'b111111111;
assign micromatrizz[29][321] = 9'b111111111;
assign micromatrizz[29][322] = 9'b111111111;
assign micromatrizz[29][323] = 9'b111111111;
assign micromatrizz[29][324] = 9'b111111111;
assign micromatrizz[29][325] = 9'b111111111;
assign micromatrizz[29][326] = 9'b111111111;
assign micromatrizz[29][327] = 9'b111111111;
assign micromatrizz[29][328] = 9'b111111111;
assign micromatrizz[29][329] = 9'b111111111;
assign micromatrizz[29][330] = 9'b111111111;
assign micromatrizz[29][331] = 9'b111111111;
assign micromatrizz[29][332] = 9'b111111111;
assign micromatrizz[29][333] = 9'b111111111;
assign micromatrizz[29][334] = 9'b111111111;
assign micromatrizz[29][335] = 9'b111111111;
assign micromatrizz[29][336] = 9'b111111111;
assign micromatrizz[29][337] = 9'b111111111;
assign micromatrizz[29][338] = 9'b111111111;
assign micromatrizz[29][339] = 9'b111111111;
assign micromatrizz[29][340] = 9'b111111111;
assign micromatrizz[29][341] = 9'b111111111;
assign micromatrizz[29][342] = 9'b111111111;
assign micromatrizz[29][343] = 9'b111111111;
assign micromatrizz[29][344] = 9'b111111111;
assign micromatrizz[29][345] = 9'b111111111;
assign micromatrizz[29][346] = 9'b111111111;
assign micromatrizz[29][347] = 9'b111111111;
assign micromatrizz[29][348] = 9'b111111111;
assign micromatrizz[29][349] = 9'b111111111;
assign micromatrizz[29][350] = 9'b111111111;
assign micromatrizz[29][351] = 9'b111111111;
assign micromatrizz[29][352] = 9'b111111111;
assign micromatrizz[29][353] = 9'b111111111;
assign micromatrizz[29][354] = 9'b111111111;
assign micromatrizz[29][355] = 9'b111111111;
assign micromatrizz[29][356] = 9'b111111111;
assign micromatrizz[29][357] = 9'b111111111;
assign micromatrizz[29][358] = 9'b111111111;
assign micromatrizz[29][359] = 9'b111111111;
assign micromatrizz[29][360] = 9'b111111111;
assign micromatrizz[29][361] = 9'b111111111;
assign micromatrizz[29][362] = 9'b111111111;
assign micromatrizz[29][363] = 9'b111111111;
assign micromatrizz[29][364] = 9'b111111111;
assign micromatrizz[29][365] = 9'b111111111;
assign micromatrizz[29][366] = 9'b111111111;
assign micromatrizz[29][367] = 9'b111111111;
assign micromatrizz[29][368] = 9'b111111111;
assign micromatrizz[29][369] = 9'b111111111;
assign micromatrizz[29][370] = 9'b111111111;
assign micromatrizz[29][371] = 9'b111111111;
assign micromatrizz[29][372] = 9'b111111111;
assign micromatrizz[29][373] = 9'b111111111;
assign micromatrizz[29][374] = 9'b111111111;
assign micromatrizz[29][375] = 9'b111111111;
assign micromatrizz[29][376] = 9'b111111111;
assign micromatrizz[29][377] = 9'b111111111;
assign micromatrizz[29][378] = 9'b111111111;
assign micromatrizz[29][379] = 9'b111111111;
assign micromatrizz[29][380] = 9'b111111111;
assign micromatrizz[29][381] = 9'b111111111;
assign micromatrizz[29][382] = 9'b111111111;
assign micromatrizz[29][383] = 9'b111111111;
assign micromatrizz[29][384] = 9'b111111111;
assign micromatrizz[29][385] = 9'b111111111;
assign micromatrizz[29][386] = 9'b111111111;
assign micromatrizz[29][387] = 9'b111111111;
assign micromatrizz[29][388] = 9'b111111111;
assign micromatrizz[29][389] = 9'b111111111;
assign micromatrizz[29][390] = 9'b111111111;
assign micromatrizz[29][391] = 9'b111111111;
assign micromatrizz[29][392] = 9'b111111111;
assign micromatrizz[29][393] = 9'b111111111;
assign micromatrizz[29][394] = 9'b111111111;
assign micromatrizz[29][395] = 9'b111111111;
assign micromatrizz[29][396] = 9'b111111111;
assign micromatrizz[29][397] = 9'b111111111;
assign micromatrizz[29][398] = 9'b111111111;
assign micromatrizz[29][399] = 9'b111111111;
assign micromatrizz[29][400] = 9'b111111111;
assign micromatrizz[29][401] = 9'b111111111;
assign micromatrizz[29][402] = 9'b111111111;
assign micromatrizz[29][403] = 9'b111111111;
assign micromatrizz[29][404] = 9'b111111111;
assign micromatrizz[29][405] = 9'b111111111;
assign micromatrizz[29][406] = 9'b111111111;
assign micromatrizz[29][407] = 9'b111111111;
assign micromatrizz[29][408] = 9'b111111111;
assign micromatrizz[29][409] = 9'b111111111;
assign micromatrizz[29][410] = 9'b111111111;
assign micromatrizz[29][411] = 9'b111111111;
assign micromatrizz[29][412] = 9'b111111111;
assign micromatrizz[29][413] = 9'b111111111;
assign micromatrizz[29][414] = 9'b111111111;
assign micromatrizz[29][415] = 9'b111111111;
assign micromatrizz[29][416] = 9'b111111111;
assign micromatrizz[29][417] = 9'b111111111;
assign micromatrizz[29][418] = 9'b111111111;
assign micromatrizz[29][419] = 9'b111111111;
assign micromatrizz[29][420] = 9'b111111111;
assign micromatrizz[29][421] = 9'b111111111;
assign micromatrizz[29][422] = 9'b111111111;
assign micromatrizz[29][423] = 9'b111111111;
assign micromatrizz[29][424] = 9'b111111111;
assign micromatrizz[29][425] = 9'b111111111;
assign micromatrizz[29][426] = 9'b111111111;
assign micromatrizz[29][427] = 9'b111111111;
assign micromatrizz[29][428] = 9'b111111111;
assign micromatrizz[29][429] = 9'b111111111;
assign micromatrizz[29][430] = 9'b111111111;
assign micromatrizz[29][431] = 9'b111111111;
assign micromatrizz[29][432] = 9'b111111111;
assign micromatrizz[29][433] = 9'b111111111;
assign micromatrizz[29][434] = 9'b111111111;
assign micromatrizz[29][435] = 9'b111111111;
assign micromatrizz[29][436] = 9'b111111111;
assign micromatrizz[29][437] = 9'b111111111;
assign micromatrizz[29][438] = 9'b111111111;
assign micromatrizz[29][439] = 9'b111111111;
assign micromatrizz[29][440] = 9'b111111111;
assign micromatrizz[29][441] = 9'b111111111;
assign micromatrizz[29][442] = 9'b111111111;
assign micromatrizz[29][443] = 9'b111111111;
assign micromatrizz[29][444] = 9'b111111111;
assign micromatrizz[29][445] = 9'b111111111;
assign micromatrizz[29][446] = 9'b111111111;
assign micromatrizz[29][447] = 9'b111111111;
assign micromatrizz[29][448] = 9'b111111111;
assign micromatrizz[29][449] = 9'b111111111;
assign micromatrizz[29][450] = 9'b111111111;
assign micromatrizz[29][451] = 9'b111111111;
assign micromatrizz[29][452] = 9'b111111111;
assign micromatrizz[29][453] = 9'b111111111;
assign micromatrizz[29][454] = 9'b111111111;
assign micromatrizz[29][455] = 9'b111111111;
assign micromatrizz[29][456] = 9'b111111111;
assign micromatrizz[29][457] = 9'b111111111;
assign micromatrizz[29][458] = 9'b111111111;
assign micromatrizz[29][459] = 9'b111111111;
assign micromatrizz[29][460] = 9'b111111111;
assign micromatrizz[29][461] = 9'b111111111;
assign micromatrizz[29][462] = 9'b111111111;
assign micromatrizz[29][463] = 9'b111111111;
assign micromatrizz[29][464] = 9'b111111111;
assign micromatrizz[29][465] = 9'b111111111;
assign micromatrizz[29][466] = 9'b111111111;
assign micromatrizz[29][467] = 9'b111111111;
assign micromatrizz[29][468] = 9'b111111111;
assign micromatrizz[29][469] = 9'b111111111;
assign micromatrizz[29][470] = 9'b111111111;
assign micromatrizz[29][471] = 9'b111111111;
assign micromatrizz[29][472] = 9'b111111111;
assign micromatrizz[29][473] = 9'b111111111;
assign micromatrizz[29][474] = 9'b111111111;
assign micromatrizz[29][475] = 9'b111111111;
assign micromatrizz[29][476] = 9'b111111111;
assign micromatrizz[29][477] = 9'b111111111;
assign micromatrizz[29][478] = 9'b111111111;
assign micromatrizz[29][479] = 9'b111111111;
assign micromatrizz[29][480] = 9'b111111111;
assign micromatrizz[29][481] = 9'b111111111;
assign micromatrizz[29][482] = 9'b111111111;
assign micromatrizz[29][483] = 9'b111111111;
assign micromatrizz[29][484] = 9'b111111111;
assign micromatrizz[29][485] = 9'b111111111;
assign micromatrizz[29][486] = 9'b111111111;
assign micromatrizz[29][487] = 9'b111111111;
assign micromatrizz[29][488] = 9'b111111111;
assign micromatrizz[29][489] = 9'b111111111;
assign micromatrizz[29][490] = 9'b111111111;
assign micromatrizz[29][491] = 9'b111111111;
assign micromatrizz[29][492] = 9'b111111111;
assign micromatrizz[29][493] = 9'b111111111;
assign micromatrizz[29][494] = 9'b111111111;
assign micromatrizz[29][495] = 9'b111111111;
assign micromatrizz[29][496] = 9'b111111111;
assign micromatrizz[29][497] = 9'b111111111;
assign micromatrizz[29][498] = 9'b111111111;
assign micromatrizz[29][499] = 9'b111111111;
assign micromatrizz[29][500] = 9'b111111111;
assign micromatrizz[29][501] = 9'b111111111;
assign micromatrizz[29][502] = 9'b111111111;
assign micromatrizz[29][503] = 9'b111111111;
assign micromatrizz[29][504] = 9'b111111111;
assign micromatrizz[29][505] = 9'b111111111;
assign micromatrizz[29][506] = 9'b111111111;
assign micromatrizz[29][507] = 9'b111111111;
assign micromatrizz[29][508] = 9'b111111111;
assign micromatrizz[29][509] = 9'b111111111;
assign micromatrizz[29][510] = 9'b111111111;
assign micromatrizz[29][511] = 9'b111111111;
assign micromatrizz[29][512] = 9'b111111111;
assign micromatrizz[29][513] = 9'b111111111;
assign micromatrizz[29][514] = 9'b111111111;
assign micromatrizz[29][515] = 9'b111111111;
assign micromatrizz[29][516] = 9'b111111111;
assign micromatrizz[29][517] = 9'b111111111;
assign micromatrizz[29][518] = 9'b111111111;
assign micromatrizz[29][519] = 9'b111111111;
assign micromatrizz[29][520] = 9'b111111111;
assign micromatrizz[29][521] = 9'b111111111;
assign micromatrizz[29][522] = 9'b111111111;
assign micromatrizz[29][523] = 9'b111111111;
assign micromatrizz[29][524] = 9'b111111111;
assign micromatrizz[29][525] = 9'b111111111;
assign micromatrizz[29][526] = 9'b111111111;
assign micromatrizz[29][527] = 9'b111111111;
assign micromatrizz[29][528] = 9'b111111111;
assign micromatrizz[29][529] = 9'b111111111;
assign micromatrizz[29][530] = 9'b111111111;
assign micromatrizz[29][531] = 9'b111111111;
assign micromatrizz[29][532] = 9'b111111111;
assign micromatrizz[29][533] = 9'b111111111;
assign micromatrizz[29][534] = 9'b111111111;
assign micromatrizz[29][535] = 9'b111111111;
assign micromatrizz[29][536] = 9'b111111111;
assign micromatrizz[29][537] = 9'b111111111;
assign micromatrizz[29][538] = 9'b111111111;
assign micromatrizz[29][539] = 9'b111111111;
assign micromatrizz[29][540] = 9'b111111111;
assign micromatrizz[29][541] = 9'b111111111;
assign micromatrizz[29][542] = 9'b111111111;
assign micromatrizz[29][543] = 9'b111111111;
assign micromatrizz[29][544] = 9'b111111111;
assign micromatrizz[29][545] = 9'b111111111;
assign micromatrizz[29][546] = 9'b111111111;
assign micromatrizz[29][547] = 9'b111111111;
assign micromatrizz[29][548] = 9'b111111111;
assign micromatrizz[29][549] = 9'b111111111;
assign micromatrizz[29][550] = 9'b111111111;
assign micromatrizz[29][551] = 9'b111111111;
assign micromatrizz[29][552] = 9'b111111111;
assign micromatrizz[29][553] = 9'b111111111;
assign micromatrizz[29][554] = 9'b111111111;
assign micromatrizz[29][555] = 9'b111111111;
assign micromatrizz[29][556] = 9'b111111111;
assign micromatrizz[29][557] = 9'b111111111;
assign micromatrizz[29][558] = 9'b111111111;
assign micromatrizz[29][559] = 9'b111111111;
assign micromatrizz[29][560] = 9'b111111111;
assign micromatrizz[29][561] = 9'b111111111;
assign micromatrizz[29][562] = 9'b111111111;
assign micromatrizz[29][563] = 9'b111111111;
assign micromatrizz[29][564] = 9'b111111111;
assign micromatrizz[29][565] = 9'b111111111;
assign micromatrizz[29][566] = 9'b111111111;
assign micromatrizz[29][567] = 9'b111111111;
assign micromatrizz[29][568] = 9'b111111111;
assign micromatrizz[29][569] = 9'b111111111;
assign micromatrizz[29][570] = 9'b111111111;
assign micromatrizz[29][571] = 9'b111111111;
assign micromatrizz[29][572] = 9'b111111111;
assign micromatrizz[29][573] = 9'b111111111;
assign micromatrizz[29][574] = 9'b111111111;
assign micromatrizz[29][575] = 9'b111111111;
assign micromatrizz[29][576] = 9'b111111111;
assign micromatrizz[29][577] = 9'b111111111;
assign micromatrizz[29][578] = 9'b111111111;
assign micromatrizz[29][579] = 9'b111111111;
assign micromatrizz[29][580] = 9'b111111111;
assign micromatrizz[29][581] = 9'b111111111;
assign micromatrizz[29][582] = 9'b111111111;
assign micromatrizz[29][583] = 9'b111111111;
assign micromatrizz[29][584] = 9'b111111111;
assign micromatrizz[29][585] = 9'b111111111;
assign micromatrizz[29][586] = 9'b111111111;
assign micromatrizz[29][587] = 9'b111111111;
assign micromatrizz[29][588] = 9'b111111111;
assign micromatrizz[29][589] = 9'b111111111;
assign micromatrizz[29][590] = 9'b111111111;
assign micromatrizz[29][591] = 9'b111111111;
assign micromatrizz[29][592] = 9'b111111111;
assign micromatrizz[29][593] = 9'b111111111;
assign micromatrizz[29][594] = 9'b111111111;
assign micromatrizz[29][595] = 9'b111111111;
assign micromatrizz[29][596] = 9'b111111111;
assign micromatrizz[29][597] = 9'b111111111;
assign micromatrizz[29][598] = 9'b111111111;
assign micromatrizz[29][599] = 9'b111111111;
assign micromatrizz[29][600] = 9'b111111111;
assign micromatrizz[29][601] = 9'b111111111;
assign micromatrizz[29][602] = 9'b111111111;
assign micromatrizz[29][603] = 9'b111111111;
assign micromatrizz[29][604] = 9'b111111111;
assign micromatrizz[29][605] = 9'b111111111;
assign micromatrizz[29][606] = 9'b111111111;
assign micromatrizz[29][607] = 9'b111111111;
assign micromatrizz[29][608] = 9'b111111111;
assign micromatrizz[29][609] = 9'b111111111;
assign micromatrizz[29][610] = 9'b111111111;
assign micromatrizz[29][611] = 9'b111111111;
assign micromatrizz[29][612] = 9'b111111111;
assign micromatrizz[29][613] = 9'b111111111;
assign micromatrizz[29][614] = 9'b111111111;
assign micromatrizz[29][615] = 9'b111111111;
assign micromatrizz[29][616] = 9'b111111111;
assign micromatrizz[29][617] = 9'b111111111;
assign micromatrizz[29][618] = 9'b111111111;
assign micromatrizz[29][619] = 9'b111111111;
assign micromatrizz[29][620] = 9'b111111111;
assign micromatrizz[29][621] = 9'b111111111;
assign micromatrizz[29][622] = 9'b111111111;
assign micromatrizz[29][623] = 9'b111111111;
assign micromatrizz[29][624] = 9'b111111111;
assign micromatrizz[29][625] = 9'b111111111;
assign micromatrizz[29][626] = 9'b111111111;
assign micromatrizz[29][627] = 9'b111111111;
assign micromatrizz[29][628] = 9'b111111111;
assign micromatrizz[29][629] = 9'b111111111;
assign micromatrizz[29][630] = 9'b111111111;
assign micromatrizz[29][631] = 9'b111111111;
assign micromatrizz[29][632] = 9'b111111111;
assign micromatrizz[29][633] = 9'b111111111;
assign micromatrizz[29][634] = 9'b111111111;
assign micromatrizz[29][635] = 9'b111111111;
assign micromatrizz[29][636] = 9'b111111111;
assign micromatrizz[29][637] = 9'b111111111;
assign micromatrizz[29][638] = 9'b111111111;
assign micromatrizz[29][639] = 9'b111111111;
assign micromatrizz[30][0] = 9'b111111111;
assign micromatrizz[30][1] = 9'b111111111;
assign micromatrizz[30][2] = 9'b111111111;
assign micromatrizz[30][3] = 9'b111111111;
assign micromatrizz[30][4] = 9'b111111111;
assign micromatrizz[30][5] = 9'b111111111;
assign micromatrizz[30][6] = 9'b111111111;
assign micromatrizz[30][7] = 9'b111111111;
assign micromatrizz[30][8] = 9'b111111111;
assign micromatrizz[30][9] = 9'b111111111;
assign micromatrizz[30][10] = 9'b111111111;
assign micromatrizz[30][11] = 9'b111111111;
assign micromatrizz[30][12] = 9'b111111111;
assign micromatrizz[30][13] = 9'b111111111;
assign micromatrizz[30][14] = 9'b111111111;
assign micromatrizz[30][15] = 9'b111111111;
assign micromatrizz[30][16] = 9'b111111111;
assign micromatrizz[30][17] = 9'b111111111;
assign micromatrizz[30][18] = 9'b111111111;
assign micromatrizz[30][19] = 9'b111111111;
assign micromatrizz[30][20] = 9'b111111111;
assign micromatrizz[30][21] = 9'b111111111;
assign micromatrizz[30][22] = 9'b111111111;
assign micromatrizz[30][23] = 9'b111111111;
assign micromatrizz[30][24] = 9'b111111111;
assign micromatrizz[30][25] = 9'b111111111;
assign micromatrizz[30][26] = 9'b111111111;
assign micromatrizz[30][27] = 9'b111111111;
assign micromatrizz[30][28] = 9'b111111111;
assign micromatrizz[30][29] = 9'b111111111;
assign micromatrizz[30][30] = 9'b111111111;
assign micromatrizz[30][31] = 9'b111111111;
assign micromatrizz[30][32] = 9'b111111111;
assign micromatrizz[30][33] = 9'b111111111;
assign micromatrizz[30][34] = 9'b111111111;
assign micromatrizz[30][35] = 9'b111111111;
assign micromatrizz[30][36] = 9'b111111111;
assign micromatrizz[30][37] = 9'b111111111;
assign micromatrizz[30][38] = 9'b111111111;
assign micromatrizz[30][39] = 9'b111111111;
assign micromatrizz[30][40] = 9'b111111111;
assign micromatrizz[30][41] = 9'b111111111;
assign micromatrizz[30][42] = 9'b111111111;
assign micromatrizz[30][43] = 9'b111111111;
assign micromatrizz[30][44] = 9'b111111111;
assign micromatrizz[30][45] = 9'b111111111;
assign micromatrizz[30][46] = 9'b111111111;
assign micromatrizz[30][47] = 9'b111111111;
assign micromatrizz[30][48] = 9'b111111111;
assign micromatrizz[30][49] = 9'b111111111;
assign micromatrizz[30][50] = 9'b111111111;
assign micromatrizz[30][51] = 9'b111111111;
assign micromatrizz[30][52] = 9'b111111111;
assign micromatrizz[30][53] = 9'b111111111;
assign micromatrizz[30][54] = 9'b111111111;
assign micromatrizz[30][55] = 9'b111111111;
assign micromatrizz[30][56] = 9'b111111111;
assign micromatrizz[30][57] = 9'b111111111;
assign micromatrizz[30][58] = 9'b111111111;
assign micromatrizz[30][59] = 9'b111111111;
assign micromatrizz[30][60] = 9'b111111111;
assign micromatrizz[30][61] = 9'b111111111;
assign micromatrizz[30][62] = 9'b111111111;
assign micromatrizz[30][63] = 9'b111111111;
assign micromatrizz[30][64] = 9'b111111111;
assign micromatrizz[30][65] = 9'b111111111;
assign micromatrizz[30][66] = 9'b111111111;
assign micromatrizz[30][67] = 9'b111111111;
assign micromatrizz[30][68] = 9'b111111111;
assign micromatrizz[30][69] = 9'b111111111;
assign micromatrizz[30][70] = 9'b111111111;
assign micromatrizz[30][71] = 9'b111111111;
assign micromatrizz[30][72] = 9'b111111111;
assign micromatrizz[30][73] = 9'b111111111;
assign micromatrizz[30][74] = 9'b111111111;
assign micromatrizz[30][75] = 9'b111111111;
assign micromatrizz[30][76] = 9'b111111111;
assign micromatrizz[30][77] = 9'b111111111;
assign micromatrizz[30][78] = 9'b111111111;
assign micromatrizz[30][79] = 9'b111111111;
assign micromatrizz[30][80] = 9'b111111111;
assign micromatrizz[30][81] = 9'b111111111;
assign micromatrizz[30][82] = 9'b111111111;
assign micromatrizz[30][83] = 9'b111111111;
assign micromatrizz[30][84] = 9'b111111111;
assign micromatrizz[30][85] = 9'b111111111;
assign micromatrizz[30][86] = 9'b111111111;
assign micromatrizz[30][87] = 9'b111111111;
assign micromatrizz[30][88] = 9'b111111111;
assign micromatrizz[30][89] = 9'b111111111;
assign micromatrizz[30][90] = 9'b111111111;
assign micromatrizz[30][91] = 9'b111111111;
assign micromatrizz[30][92] = 9'b111111111;
assign micromatrizz[30][93] = 9'b111111111;
assign micromatrizz[30][94] = 9'b111111111;
assign micromatrizz[30][95] = 9'b111111111;
assign micromatrizz[30][96] = 9'b111111111;
assign micromatrizz[30][97] = 9'b111111111;
assign micromatrizz[30][98] = 9'b111111111;
assign micromatrizz[30][99] = 9'b111111111;
assign micromatrizz[30][100] = 9'b111111111;
assign micromatrizz[30][101] = 9'b111111111;
assign micromatrizz[30][102] = 9'b111111111;
assign micromatrizz[30][103] = 9'b111111111;
assign micromatrizz[30][104] = 9'b111111111;
assign micromatrizz[30][105] = 9'b111111111;
assign micromatrizz[30][106] = 9'b111111111;
assign micromatrizz[30][107] = 9'b111111111;
assign micromatrizz[30][108] = 9'b111111111;
assign micromatrizz[30][109] = 9'b111111111;
assign micromatrizz[30][110] = 9'b111111111;
assign micromatrizz[30][111] = 9'b111111111;
assign micromatrizz[30][112] = 9'b111111111;
assign micromatrizz[30][113] = 9'b111111111;
assign micromatrizz[30][114] = 9'b111111111;
assign micromatrizz[30][115] = 9'b111111111;
assign micromatrizz[30][116] = 9'b111111111;
assign micromatrizz[30][117] = 9'b111111111;
assign micromatrizz[30][118] = 9'b111111111;
assign micromatrizz[30][119] = 9'b111111111;
assign micromatrizz[30][120] = 9'b111111111;
assign micromatrizz[30][121] = 9'b111111111;
assign micromatrizz[30][122] = 9'b111111111;
assign micromatrizz[30][123] = 9'b111111111;
assign micromatrizz[30][124] = 9'b111111111;
assign micromatrizz[30][125] = 9'b111111111;
assign micromatrizz[30][126] = 9'b111111111;
assign micromatrizz[30][127] = 9'b111111111;
assign micromatrizz[30][128] = 9'b111111111;
assign micromatrizz[30][129] = 9'b111111111;
assign micromatrizz[30][130] = 9'b111111111;
assign micromatrizz[30][131] = 9'b111111111;
assign micromatrizz[30][132] = 9'b111111111;
assign micromatrizz[30][133] = 9'b111111111;
assign micromatrizz[30][134] = 9'b111111111;
assign micromatrizz[30][135] = 9'b111111111;
assign micromatrizz[30][136] = 9'b111111111;
assign micromatrizz[30][137] = 9'b111111111;
assign micromatrizz[30][138] = 9'b111111111;
assign micromatrizz[30][139] = 9'b111111111;
assign micromatrizz[30][140] = 9'b111111111;
assign micromatrizz[30][141] = 9'b111111111;
assign micromatrizz[30][142] = 9'b111111111;
assign micromatrizz[30][143] = 9'b111111111;
assign micromatrizz[30][144] = 9'b111111111;
assign micromatrizz[30][145] = 9'b111111111;
assign micromatrizz[30][146] = 9'b111111111;
assign micromatrizz[30][147] = 9'b111111111;
assign micromatrizz[30][148] = 9'b111111111;
assign micromatrizz[30][149] = 9'b111111111;
assign micromatrizz[30][150] = 9'b111111111;
assign micromatrizz[30][151] = 9'b111111111;
assign micromatrizz[30][152] = 9'b111111111;
assign micromatrizz[30][153] = 9'b111111111;
assign micromatrizz[30][154] = 9'b111111111;
assign micromatrizz[30][155] = 9'b111111111;
assign micromatrizz[30][156] = 9'b111111111;
assign micromatrizz[30][157] = 9'b111111111;
assign micromatrizz[30][158] = 9'b111111111;
assign micromatrizz[30][159] = 9'b111111111;
assign micromatrizz[30][160] = 9'b111111111;
assign micromatrizz[30][161] = 9'b111111111;
assign micromatrizz[30][162] = 9'b111111111;
assign micromatrizz[30][163] = 9'b111111111;
assign micromatrizz[30][164] = 9'b111111111;
assign micromatrizz[30][165] = 9'b111111111;
assign micromatrizz[30][166] = 9'b111111111;
assign micromatrizz[30][167] = 9'b111111111;
assign micromatrizz[30][168] = 9'b111111111;
assign micromatrizz[30][169] = 9'b111111111;
assign micromatrizz[30][170] = 9'b111111111;
assign micromatrizz[30][171] = 9'b111111111;
assign micromatrizz[30][172] = 9'b111111111;
assign micromatrizz[30][173] = 9'b111111111;
assign micromatrizz[30][174] = 9'b111111111;
assign micromatrizz[30][175] = 9'b111111111;
assign micromatrizz[30][176] = 9'b111111111;
assign micromatrizz[30][177] = 9'b111111111;
assign micromatrizz[30][178] = 9'b111111111;
assign micromatrizz[30][179] = 9'b111111111;
assign micromatrizz[30][180] = 9'b111111111;
assign micromatrizz[30][181] = 9'b111111111;
assign micromatrizz[30][182] = 9'b111111111;
assign micromatrizz[30][183] = 9'b111111111;
assign micromatrizz[30][184] = 9'b111111111;
assign micromatrizz[30][185] = 9'b111111111;
assign micromatrizz[30][186] = 9'b111111111;
assign micromatrizz[30][187] = 9'b111111111;
assign micromatrizz[30][188] = 9'b111111111;
assign micromatrizz[30][189] = 9'b111111111;
assign micromatrizz[30][190] = 9'b111111111;
assign micromatrizz[30][191] = 9'b111111111;
assign micromatrizz[30][192] = 9'b111111111;
assign micromatrizz[30][193] = 9'b111111111;
assign micromatrizz[30][194] = 9'b111111111;
assign micromatrizz[30][195] = 9'b111111111;
assign micromatrizz[30][196] = 9'b111111111;
assign micromatrizz[30][197] = 9'b111111111;
assign micromatrizz[30][198] = 9'b111111111;
assign micromatrizz[30][199] = 9'b111111111;
assign micromatrizz[30][200] = 9'b111111111;
assign micromatrizz[30][201] = 9'b111111111;
assign micromatrizz[30][202] = 9'b111111111;
assign micromatrizz[30][203] = 9'b111111111;
assign micromatrizz[30][204] = 9'b111111111;
assign micromatrizz[30][205] = 9'b111111111;
assign micromatrizz[30][206] = 9'b111111111;
assign micromatrizz[30][207] = 9'b111111111;
assign micromatrizz[30][208] = 9'b111111111;
assign micromatrizz[30][209] = 9'b111111111;
assign micromatrizz[30][210] = 9'b111111111;
assign micromatrizz[30][211] = 9'b111111111;
assign micromatrizz[30][212] = 9'b111111111;
assign micromatrizz[30][213] = 9'b111111111;
assign micromatrizz[30][214] = 9'b111111111;
assign micromatrizz[30][215] = 9'b111111111;
assign micromatrizz[30][216] = 9'b111111111;
assign micromatrizz[30][217] = 9'b111111111;
assign micromatrizz[30][218] = 9'b111111111;
assign micromatrizz[30][219] = 9'b111111111;
assign micromatrizz[30][220] = 9'b111111111;
assign micromatrizz[30][221] = 9'b111111111;
assign micromatrizz[30][222] = 9'b111111111;
assign micromatrizz[30][223] = 9'b111111111;
assign micromatrizz[30][224] = 9'b111111111;
assign micromatrizz[30][225] = 9'b111111111;
assign micromatrizz[30][226] = 9'b111111111;
assign micromatrizz[30][227] = 9'b111111111;
assign micromatrizz[30][228] = 9'b111111111;
assign micromatrizz[30][229] = 9'b111111111;
assign micromatrizz[30][230] = 9'b111111111;
assign micromatrizz[30][231] = 9'b111111111;
assign micromatrizz[30][232] = 9'b111111111;
assign micromatrizz[30][233] = 9'b111111111;
assign micromatrizz[30][234] = 9'b111111111;
assign micromatrizz[30][235] = 9'b111111111;
assign micromatrizz[30][236] = 9'b111111111;
assign micromatrizz[30][237] = 9'b111111111;
assign micromatrizz[30][238] = 9'b111111111;
assign micromatrizz[30][239] = 9'b111111111;
assign micromatrizz[30][240] = 9'b111111111;
assign micromatrizz[30][241] = 9'b111111111;
assign micromatrizz[30][242] = 9'b111111111;
assign micromatrizz[30][243] = 9'b111111111;
assign micromatrizz[30][244] = 9'b111111111;
assign micromatrizz[30][245] = 9'b111111111;
assign micromatrizz[30][246] = 9'b111111111;
assign micromatrizz[30][247] = 9'b111111111;
assign micromatrizz[30][248] = 9'b111111111;
assign micromatrizz[30][249] = 9'b111111111;
assign micromatrizz[30][250] = 9'b111111111;
assign micromatrizz[30][251] = 9'b111111111;
assign micromatrizz[30][252] = 9'b111111111;
assign micromatrizz[30][253] = 9'b111111111;
assign micromatrizz[30][254] = 9'b111111111;
assign micromatrizz[30][255] = 9'b111111111;
assign micromatrizz[30][256] = 9'b111111111;
assign micromatrizz[30][257] = 9'b111111111;
assign micromatrizz[30][258] = 9'b111111111;
assign micromatrizz[30][259] = 9'b111111111;
assign micromatrizz[30][260] = 9'b111111111;
assign micromatrizz[30][261] = 9'b111111111;
assign micromatrizz[30][262] = 9'b111111111;
assign micromatrizz[30][263] = 9'b111111111;
assign micromatrizz[30][264] = 9'b111111111;
assign micromatrizz[30][265] = 9'b111111111;
assign micromatrizz[30][266] = 9'b111111111;
assign micromatrizz[30][267] = 9'b111111111;
assign micromatrizz[30][268] = 9'b111111111;
assign micromatrizz[30][269] = 9'b111111111;
assign micromatrizz[30][270] = 9'b111110010;
assign micromatrizz[30][271] = 9'b111110010;
assign micromatrizz[30][272] = 9'b111110010;
assign micromatrizz[30][273] = 9'b111110010;
assign micromatrizz[30][274] = 9'b111110010;
assign micromatrizz[30][275] = 9'b111110011;
assign micromatrizz[30][276] = 9'b111110011;
assign micromatrizz[30][277] = 9'b111110011;
assign micromatrizz[30][278] = 9'b111110011;
assign micromatrizz[30][279] = 9'b111111111;
assign micromatrizz[30][280] = 9'b111111111;
assign micromatrizz[30][281] = 9'b111111111;
assign micromatrizz[30][282] = 9'b111111111;
assign micromatrizz[30][283] = 9'b111111111;
assign micromatrizz[30][284] = 9'b111111111;
assign micromatrizz[30][285] = 9'b111111111;
assign micromatrizz[30][286] = 9'b111111111;
assign micromatrizz[30][287] = 9'b111111111;
assign micromatrizz[30][288] = 9'b111111111;
assign micromatrizz[30][289] = 9'b111111111;
assign micromatrizz[30][290] = 9'b111110010;
assign micromatrizz[30][291] = 9'b111110010;
assign micromatrizz[30][292] = 9'b111110011;
assign micromatrizz[30][293] = 9'b111110011;
assign micromatrizz[30][294] = 9'b111110011;
assign micromatrizz[30][295] = 9'b111110011;
assign micromatrizz[30][296] = 9'b111110011;
assign micromatrizz[30][297] = 9'b111110111;
assign micromatrizz[30][298] = 9'b111111111;
assign micromatrizz[30][299] = 9'b111111111;
assign micromatrizz[30][300] = 9'b111111111;
assign micromatrizz[30][301] = 9'b111111111;
assign micromatrizz[30][302] = 9'b111111111;
assign micromatrizz[30][303] = 9'b111111111;
assign micromatrizz[30][304] = 9'b111111111;
assign micromatrizz[30][305] = 9'b111110111;
assign micromatrizz[30][306] = 9'b111111111;
assign micromatrizz[30][307] = 9'b111111111;
assign micromatrizz[30][308] = 9'b111111111;
assign micromatrizz[30][309] = 9'b111111111;
assign micromatrizz[30][310] = 9'b111110111;
assign micromatrizz[30][311] = 9'b111110010;
assign micromatrizz[30][312] = 9'b111110010;
assign micromatrizz[30][313] = 9'b111110010;
assign micromatrizz[30][314] = 9'b111110010;
assign micromatrizz[30][315] = 9'b111110010;
assign micromatrizz[30][316] = 9'b111110011;
assign micromatrizz[30][317] = 9'b111110011;
assign micromatrizz[30][318] = 9'b111110011;
assign micromatrizz[30][319] = 9'b111110011;
assign micromatrizz[30][320] = 9'b111110111;
assign micromatrizz[30][321] = 9'b111111111;
assign micromatrizz[30][322] = 9'b111111111;
assign micromatrizz[30][323] = 9'b111111111;
assign micromatrizz[30][324] = 9'b111111111;
assign micromatrizz[30][325] = 9'b111111111;
assign micromatrizz[30][326] = 9'b111111111;
assign micromatrizz[30][327] = 9'b111111111;
assign micromatrizz[30][328] = 9'b111111111;
assign micromatrizz[30][329] = 9'b111111111;
assign micromatrizz[30][330] = 9'b111111111;
assign micromatrizz[30][331] = 9'b111111111;
assign micromatrizz[30][332] = 9'b111111111;
assign micromatrizz[30][333] = 9'b111111111;
assign micromatrizz[30][334] = 9'b111111111;
assign micromatrizz[30][335] = 9'b111111111;
assign micromatrizz[30][336] = 9'b111111111;
assign micromatrizz[30][337] = 9'b111111111;
assign micromatrizz[30][338] = 9'b111111111;
assign micromatrizz[30][339] = 9'b111111111;
assign micromatrizz[30][340] = 9'b111111111;
assign micromatrizz[30][341] = 9'b111111111;
assign micromatrizz[30][342] = 9'b111111111;
assign micromatrizz[30][343] = 9'b111111111;
assign micromatrizz[30][344] = 9'b111111111;
assign micromatrizz[30][345] = 9'b111111111;
assign micromatrizz[30][346] = 9'b111111111;
assign micromatrizz[30][347] = 9'b111111111;
assign micromatrizz[30][348] = 9'b111111111;
assign micromatrizz[30][349] = 9'b111111111;
assign micromatrizz[30][350] = 9'b111111111;
assign micromatrizz[30][351] = 9'b111111111;
assign micromatrizz[30][352] = 9'b111111111;
assign micromatrizz[30][353] = 9'b111111111;
assign micromatrizz[30][354] = 9'b111111111;
assign micromatrizz[30][355] = 9'b111111111;
assign micromatrizz[30][356] = 9'b111111111;
assign micromatrizz[30][357] = 9'b111111111;
assign micromatrizz[30][358] = 9'b111111111;
assign micromatrizz[30][359] = 9'b111111111;
assign micromatrizz[30][360] = 9'b111111111;
assign micromatrizz[30][361] = 9'b111111111;
assign micromatrizz[30][362] = 9'b111111111;
assign micromatrizz[30][363] = 9'b111111111;
assign micromatrizz[30][364] = 9'b111111111;
assign micromatrizz[30][365] = 9'b111111111;
assign micromatrizz[30][366] = 9'b111111111;
assign micromatrizz[30][367] = 9'b111111111;
assign micromatrizz[30][368] = 9'b111111111;
assign micromatrizz[30][369] = 9'b111111111;
assign micromatrizz[30][370] = 9'b111111111;
assign micromatrizz[30][371] = 9'b111111111;
assign micromatrizz[30][372] = 9'b111111111;
assign micromatrizz[30][373] = 9'b111111111;
assign micromatrizz[30][374] = 9'b111111111;
assign micromatrizz[30][375] = 9'b111111111;
assign micromatrizz[30][376] = 9'b111111111;
assign micromatrizz[30][377] = 9'b111111111;
assign micromatrizz[30][378] = 9'b111111111;
assign micromatrizz[30][379] = 9'b111111111;
assign micromatrizz[30][380] = 9'b111111111;
assign micromatrizz[30][381] = 9'b111111111;
assign micromatrizz[30][382] = 9'b111111111;
assign micromatrizz[30][383] = 9'b111111111;
assign micromatrizz[30][384] = 9'b111111111;
assign micromatrizz[30][385] = 9'b111111111;
assign micromatrizz[30][386] = 9'b111111111;
assign micromatrizz[30][387] = 9'b111111111;
assign micromatrizz[30][388] = 9'b111111111;
assign micromatrizz[30][389] = 9'b111111111;
assign micromatrizz[30][390] = 9'b111111111;
assign micromatrizz[30][391] = 9'b111111111;
assign micromatrizz[30][392] = 9'b111111111;
assign micromatrizz[30][393] = 9'b111111111;
assign micromatrizz[30][394] = 9'b111111111;
assign micromatrizz[30][395] = 9'b111111111;
assign micromatrizz[30][396] = 9'b111111111;
assign micromatrizz[30][397] = 9'b111111111;
assign micromatrizz[30][398] = 9'b111111111;
assign micromatrizz[30][399] = 9'b111111111;
assign micromatrizz[30][400] = 9'b111111111;
assign micromatrizz[30][401] = 9'b111111111;
assign micromatrizz[30][402] = 9'b111111111;
assign micromatrizz[30][403] = 9'b111111111;
assign micromatrizz[30][404] = 9'b111111111;
assign micromatrizz[30][405] = 9'b111111111;
assign micromatrizz[30][406] = 9'b111111111;
assign micromatrizz[30][407] = 9'b111111111;
assign micromatrizz[30][408] = 9'b111111111;
assign micromatrizz[30][409] = 9'b111111111;
assign micromatrizz[30][410] = 9'b111111111;
assign micromatrizz[30][411] = 9'b111111111;
assign micromatrizz[30][412] = 9'b111111111;
assign micromatrizz[30][413] = 9'b111111111;
assign micromatrizz[30][414] = 9'b111111111;
assign micromatrizz[30][415] = 9'b111111111;
assign micromatrizz[30][416] = 9'b111111111;
assign micromatrizz[30][417] = 9'b111111111;
assign micromatrizz[30][418] = 9'b111111111;
assign micromatrizz[30][419] = 9'b111111111;
assign micromatrizz[30][420] = 9'b111111111;
assign micromatrizz[30][421] = 9'b111111111;
assign micromatrizz[30][422] = 9'b111111111;
assign micromatrizz[30][423] = 9'b111111111;
assign micromatrizz[30][424] = 9'b111111111;
assign micromatrizz[30][425] = 9'b111111111;
assign micromatrizz[30][426] = 9'b111111111;
assign micromatrizz[30][427] = 9'b111111111;
assign micromatrizz[30][428] = 9'b111111111;
assign micromatrizz[30][429] = 9'b111111111;
assign micromatrizz[30][430] = 9'b111111111;
assign micromatrizz[30][431] = 9'b111111111;
assign micromatrizz[30][432] = 9'b111111111;
assign micromatrizz[30][433] = 9'b111111111;
assign micromatrizz[30][434] = 9'b111111111;
assign micromatrizz[30][435] = 9'b111111111;
assign micromatrizz[30][436] = 9'b111111111;
assign micromatrizz[30][437] = 9'b111111111;
assign micromatrizz[30][438] = 9'b111111111;
assign micromatrizz[30][439] = 9'b111111111;
assign micromatrizz[30][440] = 9'b111111111;
assign micromatrizz[30][441] = 9'b111111111;
assign micromatrizz[30][442] = 9'b111111111;
assign micromatrizz[30][443] = 9'b111111111;
assign micromatrizz[30][444] = 9'b111111111;
assign micromatrizz[30][445] = 9'b111111111;
assign micromatrizz[30][446] = 9'b111111111;
assign micromatrizz[30][447] = 9'b111111111;
assign micromatrizz[30][448] = 9'b111111111;
assign micromatrizz[30][449] = 9'b111111111;
assign micromatrizz[30][450] = 9'b111111111;
assign micromatrizz[30][451] = 9'b111111111;
assign micromatrizz[30][452] = 9'b111111111;
assign micromatrizz[30][453] = 9'b111111111;
assign micromatrizz[30][454] = 9'b111111111;
assign micromatrizz[30][455] = 9'b111111111;
assign micromatrizz[30][456] = 9'b111111111;
assign micromatrizz[30][457] = 9'b111111111;
assign micromatrizz[30][458] = 9'b111111111;
assign micromatrizz[30][459] = 9'b111111111;
assign micromatrizz[30][460] = 9'b111111111;
assign micromatrizz[30][461] = 9'b111111111;
assign micromatrizz[30][462] = 9'b111111111;
assign micromatrizz[30][463] = 9'b111111111;
assign micromatrizz[30][464] = 9'b111111111;
assign micromatrizz[30][465] = 9'b111111111;
assign micromatrizz[30][466] = 9'b111111111;
assign micromatrizz[30][467] = 9'b111111111;
assign micromatrizz[30][468] = 9'b111111111;
assign micromatrizz[30][469] = 9'b111111111;
assign micromatrizz[30][470] = 9'b111111111;
assign micromatrizz[30][471] = 9'b111111111;
assign micromatrizz[30][472] = 9'b111111111;
assign micromatrizz[30][473] = 9'b111111111;
assign micromatrizz[30][474] = 9'b111111111;
assign micromatrizz[30][475] = 9'b111111111;
assign micromatrizz[30][476] = 9'b111111111;
assign micromatrizz[30][477] = 9'b111111111;
assign micromatrizz[30][478] = 9'b111111111;
assign micromatrizz[30][479] = 9'b111111111;
assign micromatrizz[30][480] = 9'b111111111;
assign micromatrizz[30][481] = 9'b111111111;
assign micromatrizz[30][482] = 9'b111111111;
assign micromatrizz[30][483] = 9'b111111111;
assign micromatrizz[30][484] = 9'b111111111;
assign micromatrizz[30][485] = 9'b111111111;
assign micromatrizz[30][486] = 9'b111111111;
assign micromatrizz[30][487] = 9'b111111111;
assign micromatrizz[30][488] = 9'b111111111;
assign micromatrizz[30][489] = 9'b111111111;
assign micromatrizz[30][490] = 9'b111111111;
assign micromatrizz[30][491] = 9'b111111111;
assign micromatrizz[30][492] = 9'b111111111;
assign micromatrizz[30][493] = 9'b111111111;
assign micromatrizz[30][494] = 9'b111111111;
assign micromatrizz[30][495] = 9'b111111111;
assign micromatrizz[30][496] = 9'b111111111;
assign micromatrizz[30][497] = 9'b111111111;
assign micromatrizz[30][498] = 9'b111111111;
assign micromatrizz[30][499] = 9'b111111111;
assign micromatrizz[30][500] = 9'b111111111;
assign micromatrizz[30][501] = 9'b111111111;
assign micromatrizz[30][502] = 9'b111111111;
assign micromatrizz[30][503] = 9'b111111111;
assign micromatrizz[30][504] = 9'b111111111;
assign micromatrizz[30][505] = 9'b111111111;
assign micromatrizz[30][506] = 9'b111111111;
assign micromatrizz[30][507] = 9'b111111111;
assign micromatrizz[30][508] = 9'b111111111;
assign micromatrizz[30][509] = 9'b111111111;
assign micromatrizz[30][510] = 9'b111111111;
assign micromatrizz[30][511] = 9'b111111111;
assign micromatrizz[30][512] = 9'b111111111;
assign micromatrizz[30][513] = 9'b111111111;
assign micromatrizz[30][514] = 9'b111111111;
assign micromatrizz[30][515] = 9'b111111111;
assign micromatrizz[30][516] = 9'b111111111;
assign micromatrizz[30][517] = 9'b111111111;
assign micromatrizz[30][518] = 9'b111111111;
assign micromatrizz[30][519] = 9'b111111111;
assign micromatrizz[30][520] = 9'b111111111;
assign micromatrizz[30][521] = 9'b111111111;
assign micromatrizz[30][522] = 9'b111111111;
assign micromatrizz[30][523] = 9'b111111111;
assign micromatrizz[30][524] = 9'b111111111;
assign micromatrizz[30][525] = 9'b111111111;
assign micromatrizz[30][526] = 9'b111111111;
assign micromatrizz[30][527] = 9'b111111111;
assign micromatrizz[30][528] = 9'b111111111;
assign micromatrizz[30][529] = 9'b111111111;
assign micromatrizz[30][530] = 9'b111111111;
assign micromatrizz[30][531] = 9'b111111111;
assign micromatrizz[30][532] = 9'b111111111;
assign micromatrizz[30][533] = 9'b111111111;
assign micromatrizz[30][534] = 9'b111111111;
assign micromatrizz[30][535] = 9'b111111111;
assign micromatrizz[30][536] = 9'b111111111;
assign micromatrizz[30][537] = 9'b111111111;
assign micromatrizz[30][538] = 9'b111111111;
assign micromatrizz[30][539] = 9'b111111111;
assign micromatrizz[30][540] = 9'b111111111;
assign micromatrizz[30][541] = 9'b111111111;
assign micromatrizz[30][542] = 9'b111111111;
assign micromatrizz[30][543] = 9'b111111111;
assign micromatrizz[30][544] = 9'b111111111;
assign micromatrizz[30][545] = 9'b111111111;
assign micromatrizz[30][546] = 9'b111111111;
assign micromatrizz[30][547] = 9'b111111111;
assign micromatrizz[30][548] = 9'b111111111;
assign micromatrizz[30][549] = 9'b111111111;
assign micromatrizz[30][550] = 9'b111111111;
assign micromatrizz[30][551] = 9'b111111111;
assign micromatrizz[30][552] = 9'b111111111;
assign micromatrizz[30][553] = 9'b111111111;
assign micromatrizz[30][554] = 9'b111111111;
assign micromatrizz[30][555] = 9'b111111111;
assign micromatrizz[30][556] = 9'b111111111;
assign micromatrizz[30][557] = 9'b111111111;
assign micromatrizz[30][558] = 9'b111111111;
assign micromatrizz[30][559] = 9'b111111111;
assign micromatrizz[30][560] = 9'b111111111;
assign micromatrizz[30][561] = 9'b111111111;
assign micromatrizz[30][562] = 9'b111111111;
assign micromatrizz[30][563] = 9'b111111111;
assign micromatrizz[30][564] = 9'b111111111;
assign micromatrizz[30][565] = 9'b111111111;
assign micromatrizz[30][566] = 9'b111111111;
assign micromatrizz[30][567] = 9'b111111111;
assign micromatrizz[30][568] = 9'b111111111;
assign micromatrizz[30][569] = 9'b111111111;
assign micromatrizz[30][570] = 9'b111111111;
assign micromatrizz[30][571] = 9'b111111111;
assign micromatrizz[30][572] = 9'b111111111;
assign micromatrizz[30][573] = 9'b111111111;
assign micromatrizz[30][574] = 9'b111111111;
assign micromatrizz[30][575] = 9'b111111111;
assign micromatrizz[30][576] = 9'b111111111;
assign micromatrizz[30][577] = 9'b111111111;
assign micromatrizz[30][578] = 9'b111111111;
assign micromatrizz[30][579] = 9'b111111111;
assign micromatrizz[30][580] = 9'b111111111;
assign micromatrizz[30][581] = 9'b111111111;
assign micromatrizz[30][582] = 9'b111111111;
assign micromatrizz[30][583] = 9'b111111111;
assign micromatrizz[30][584] = 9'b111111111;
assign micromatrizz[30][585] = 9'b111111111;
assign micromatrizz[30][586] = 9'b111111111;
assign micromatrizz[30][587] = 9'b111111111;
assign micromatrizz[30][588] = 9'b111111111;
assign micromatrizz[30][589] = 9'b111111111;
assign micromatrizz[30][590] = 9'b111111111;
assign micromatrizz[30][591] = 9'b111111111;
assign micromatrizz[30][592] = 9'b111111111;
assign micromatrizz[30][593] = 9'b111111111;
assign micromatrizz[30][594] = 9'b111111111;
assign micromatrizz[30][595] = 9'b111111111;
assign micromatrizz[30][596] = 9'b111111111;
assign micromatrizz[30][597] = 9'b111111111;
assign micromatrizz[30][598] = 9'b111111111;
assign micromatrizz[30][599] = 9'b111111111;
assign micromatrizz[30][600] = 9'b111111111;
assign micromatrizz[30][601] = 9'b111111111;
assign micromatrizz[30][602] = 9'b111111111;
assign micromatrizz[30][603] = 9'b111111111;
assign micromatrizz[30][604] = 9'b111111111;
assign micromatrizz[30][605] = 9'b111111111;
assign micromatrizz[30][606] = 9'b111111111;
assign micromatrizz[30][607] = 9'b111111111;
assign micromatrizz[30][608] = 9'b111111111;
assign micromatrizz[30][609] = 9'b111111111;
assign micromatrizz[30][610] = 9'b111111111;
assign micromatrizz[30][611] = 9'b111111111;
assign micromatrizz[30][612] = 9'b111111111;
assign micromatrizz[30][613] = 9'b111111111;
assign micromatrizz[30][614] = 9'b111111111;
assign micromatrizz[30][615] = 9'b111111111;
assign micromatrizz[30][616] = 9'b111111111;
assign micromatrizz[30][617] = 9'b111111111;
assign micromatrizz[30][618] = 9'b111111111;
assign micromatrizz[30][619] = 9'b111111111;
assign micromatrizz[30][620] = 9'b111111111;
assign micromatrizz[30][621] = 9'b111111111;
assign micromatrizz[30][622] = 9'b111111111;
assign micromatrizz[30][623] = 9'b111111111;
assign micromatrizz[30][624] = 9'b111111111;
assign micromatrizz[30][625] = 9'b111111111;
assign micromatrizz[30][626] = 9'b111111111;
assign micromatrizz[30][627] = 9'b111111111;
assign micromatrizz[30][628] = 9'b111111111;
assign micromatrizz[30][629] = 9'b111111111;
assign micromatrizz[30][630] = 9'b111111111;
assign micromatrizz[30][631] = 9'b111111111;
assign micromatrizz[30][632] = 9'b111111111;
assign micromatrizz[30][633] = 9'b111111111;
assign micromatrizz[30][634] = 9'b111111111;
assign micromatrizz[30][635] = 9'b111111111;
assign micromatrizz[30][636] = 9'b111111111;
assign micromatrizz[30][637] = 9'b111111111;
assign micromatrizz[30][638] = 9'b111111111;
assign micromatrizz[30][639] = 9'b111111111;
assign micromatrizz[31][0] = 9'b111111111;
assign micromatrizz[31][1] = 9'b111111111;
assign micromatrizz[31][2] = 9'b111111111;
assign micromatrizz[31][3] = 9'b111111111;
assign micromatrizz[31][4] = 9'b111111111;
assign micromatrizz[31][5] = 9'b111111111;
assign micromatrizz[31][6] = 9'b111111111;
assign micromatrizz[31][7] = 9'b111111111;
assign micromatrizz[31][8] = 9'b111111111;
assign micromatrizz[31][9] = 9'b111111111;
assign micromatrizz[31][10] = 9'b111111111;
assign micromatrizz[31][11] = 9'b111111111;
assign micromatrizz[31][12] = 9'b111111111;
assign micromatrizz[31][13] = 9'b111111111;
assign micromatrizz[31][14] = 9'b111111111;
assign micromatrizz[31][15] = 9'b111111111;
assign micromatrizz[31][16] = 9'b111111111;
assign micromatrizz[31][17] = 9'b111111111;
assign micromatrizz[31][18] = 9'b111111111;
assign micromatrizz[31][19] = 9'b111111111;
assign micromatrizz[31][20] = 9'b111111111;
assign micromatrizz[31][21] = 9'b111111111;
assign micromatrizz[31][22] = 9'b111111111;
assign micromatrizz[31][23] = 9'b111111111;
assign micromatrizz[31][24] = 9'b111111111;
assign micromatrizz[31][25] = 9'b111111111;
assign micromatrizz[31][26] = 9'b111111111;
assign micromatrizz[31][27] = 9'b111111111;
assign micromatrizz[31][28] = 9'b111111111;
assign micromatrizz[31][29] = 9'b111111111;
assign micromatrizz[31][30] = 9'b111111111;
assign micromatrizz[31][31] = 9'b111111111;
assign micromatrizz[31][32] = 9'b111111111;
assign micromatrizz[31][33] = 9'b111111111;
assign micromatrizz[31][34] = 9'b111111111;
assign micromatrizz[31][35] = 9'b111111111;
assign micromatrizz[31][36] = 9'b111111111;
assign micromatrizz[31][37] = 9'b111111111;
assign micromatrizz[31][38] = 9'b111111111;
assign micromatrizz[31][39] = 9'b111111111;
assign micromatrizz[31][40] = 9'b111111111;
assign micromatrizz[31][41] = 9'b111111111;
assign micromatrizz[31][42] = 9'b111111111;
assign micromatrizz[31][43] = 9'b111111111;
assign micromatrizz[31][44] = 9'b111111111;
assign micromatrizz[31][45] = 9'b111111111;
assign micromatrizz[31][46] = 9'b111111111;
assign micromatrizz[31][47] = 9'b111111111;
assign micromatrizz[31][48] = 9'b111111111;
assign micromatrizz[31][49] = 9'b111111111;
assign micromatrizz[31][50] = 9'b111111111;
assign micromatrizz[31][51] = 9'b111111111;
assign micromatrizz[31][52] = 9'b111111111;
assign micromatrizz[31][53] = 9'b111111111;
assign micromatrizz[31][54] = 9'b111111111;
assign micromatrizz[31][55] = 9'b111111111;
assign micromatrizz[31][56] = 9'b111111111;
assign micromatrizz[31][57] = 9'b111111111;
assign micromatrizz[31][58] = 9'b111111111;
assign micromatrizz[31][59] = 9'b111111111;
assign micromatrizz[31][60] = 9'b111111111;
assign micromatrizz[31][61] = 9'b111111111;
assign micromatrizz[31][62] = 9'b111111111;
assign micromatrizz[31][63] = 9'b111111111;
assign micromatrizz[31][64] = 9'b111111111;
assign micromatrizz[31][65] = 9'b111111111;
assign micromatrizz[31][66] = 9'b111111111;
assign micromatrizz[31][67] = 9'b111111111;
assign micromatrizz[31][68] = 9'b111111111;
assign micromatrizz[31][69] = 9'b111111111;
assign micromatrizz[31][70] = 9'b111111111;
assign micromatrizz[31][71] = 9'b111111111;
assign micromatrizz[31][72] = 9'b111111111;
assign micromatrizz[31][73] = 9'b111111111;
assign micromatrizz[31][74] = 9'b111111111;
assign micromatrizz[31][75] = 9'b111111111;
assign micromatrizz[31][76] = 9'b111111111;
assign micromatrizz[31][77] = 9'b111111111;
assign micromatrizz[31][78] = 9'b111111111;
assign micromatrizz[31][79] = 9'b111111111;
assign micromatrizz[31][80] = 9'b111111111;
assign micromatrizz[31][81] = 9'b111111111;
assign micromatrizz[31][82] = 9'b111111111;
assign micromatrizz[31][83] = 9'b111111111;
assign micromatrizz[31][84] = 9'b111111111;
assign micromatrizz[31][85] = 9'b111111111;
assign micromatrizz[31][86] = 9'b111111111;
assign micromatrizz[31][87] = 9'b111111111;
assign micromatrizz[31][88] = 9'b111111111;
assign micromatrizz[31][89] = 9'b111111111;
assign micromatrizz[31][90] = 9'b111111111;
assign micromatrizz[31][91] = 9'b111111111;
assign micromatrizz[31][92] = 9'b111111111;
assign micromatrizz[31][93] = 9'b111111111;
assign micromatrizz[31][94] = 9'b111111111;
assign micromatrizz[31][95] = 9'b111111111;
assign micromatrizz[31][96] = 9'b111111111;
assign micromatrizz[31][97] = 9'b111111111;
assign micromatrizz[31][98] = 9'b111111111;
assign micromatrizz[31][99] = 9'b111111111;
assign micromatrizz[31][100] = 9'b111111111;
assign micromatrizz[31][101] = 9'b111111111;
assign micromatrizz[31][102] = 9'b111111111;
assign micromatrizz[31][103] = 9'b111111111;
assign micromatrizz[31][104] = 9'b111111111;
assign micromatrizz[31][105] = 9'b111111111;
assign micromatrizz[31][106] = 9'b111111111;
assign micromatrizz[31][107] = 9'b111111111;
assign micromatrizz[31][108] = 9'b111111111;
assign micromatrizz[31][109] = 9'b111111111;
assign micromatrizz[31][110] = 9'b111111111;
assign micromatrizz[31][111] = 9'b111111111;
assign micromatrizz[31][112] = 9'b111111111;
assign micromatrizz[31][113] = 9'b111111111;
assign micromatrizz[31][114] = 9'b111111111;
assign micromatrizz[31][115] = 9'b111111111;
assign micromatrizz[31][116] = 9'b111111111;
assign micromatrizz[31][117] = 9'b111111111;
assign micromatrizz[31][118] = 9'b111111111;
assign micromatrizz[31][119] = 9'b111111111;
assign micromatrizz[31][120] = 9'b111111111;
assign micromatrizz[31][121] = 9'b111111111;
assign micromatrizz[31][122] = 9'b111111111;
assign micromatrizz[31][123] = 9'b111111111;
assign micromatrizz[31][124] = 9'b111111111;
assign micromatrizz[31][125] = 9'b111111111;
assign micromatrizz[31][126] = 9'b111111111;
assign micromatrizz[31][127] = 9'b111111111;
assign micromatrizz[31][128] = 9'b111111111;
assign micromatrizz[31][129] = 9'b111111111;
assign micromatrizz[31][130] = 9'b111111111;
assign micromatrizz[31][131] = 9'b111111111;
assign micromatrizz[31][132] = 9'b111111111;
assign micromatrizz[31][133] = 9'b111111111;
assign micromatrizz[31][134] = 9'b111111111;
assign micromatrizz[31][135] = 9'b111111111;
assign micromatrizz[31][136] = 9'b111111111;
assign micromatrizz[31][137] = 9'b111111111;
assign micromatrizz[31][138] = 9'b111111111;
assign micromatrizz[31][139] = 9'b111111111;
assign micromatrizz[31][140] = 9'b111111111;
assign micromatrizz[31][141] = 9'b111111111;
assign micromatrizz[31][142] = 9'b111111111;
assign micromatrizz[31][143] = 9'b111111111;
assign micromatrizz[31][144] = 9'b111111111;
assign micromatrizz[31][145] = 9'b111111111;
assign micromatrizz[31][146] = 9'b111111111;
assign micromatrizz[31][147] = 9'b111111111;
assign micromatrizz[31][148] = 9'b111111111;
assign micromatrizz[31][149] = 9'b111111111;
assign micromatrizz[31][150] = 9'b111111111;
assign micromatrizz[31][151] = 9'b111111111;
assign micromatrizz[31][152] = 9'b111111111;
assign micromatrizz[31][153] = 9'b111111111;
assign micromatrizz[31][154] = 9'b111111111;
assign micromatrizz[31][155] = 9'b111111111;
assign micromatrizz[31][156] = 9'b111111111;
assign micromatrizz[31][157] = 9'b111111111;
assign micromatrizz[31][158] = 9'b111111111;
assign micromatrizz[31][159] = 9'b111111111;
assign micromatrizz[31][160] = 9'b111111111;
assign micromatrizz[31][161] = 9'b111111111;
assign micromatrizz[31][162] = 9'b111111111;
assign micromatrizz[31][163] = 9'b111111111;
assign micromatrizz[31][164] = 9'b111111111;
assign micromatrizz[31][165] = 9'b111111111;
assign micromatrizz[31][166] = 9'b111111111;
assign micromatrizz[31][167] = 9'b111111111;
assign micromatrizz[31][168] = 9'b111111111;
assign micromatrizz[31][169] = 9'b111111111;
assign micromatrizz[31][170] = 9'b111111111;
assign micromatrizz[31][171] = 9'b111111111;
assign micromatrizz[31][172] = 9'b111111111;
assign micromatrizz[31][173] = 9'b111111111;
assign micromatrizz[31][174] = 9'b111111111;
assign micromatrizz[31][175] = 9'b111111111;
assign micromatrizz[31][176] = 9'b111111111;
assign micromatrizz[31][177] = 9'b111111111;
assign micromatrizz[31][178] = 9'b111111111;
assign micromatrizz[31][179] = 9'b111111111;
assign micromatrizz[31][180] = 9'b111111111;
assign micromatrizz[31][181] = 9'b111111111;
assign micromatrizz[31][182] = 9'b111111111;
assign micromatrizz[31][183] = 9'b111111111;
assign micromatrizz[31][184] = 9'b111111111;
assign micromatrizz[31][185] = 9'b111111111;
assign micromatrizz[31][186] = 9'b111111111;
assign micromatrizz[31][187] = 9'b111111111;
assign micromatrizz[31][188] = 9'b111111111;
assign micromatrizz[31][189] = 9'b111111111;
assign micromatrizz[31][190] = 9'b111111111;
assign micromatrizz[31][191] = 9'b111111111;
assign micromatrizz[31][192] = 9'b111111111;
assign micromatrizz[31][193] = 9'b111111111;
assign micromatrizz[31][194] = 9'b111111111;
assign micromatrizz[31][195] = 9'b111111111;
assign micromatrizz[31][196] = 9'b111111111;
assign micromatrizz[31][197] = 9'b111111111;
assign micromatrizz[31][198] = 9'b111111111;
assign micromatrizz[31][199] = 9'b111111111;
assign micromatrizz[31][200] = 9'b111111111;
assign micromatrizz[31][201] = 9'b111111111;
assign micromatrizz[31][202] = 9'b111111111;
assign micromatrizz[31][203] = 9'b111111111;
assign micromatrizz[31][204] = 9'b111111111;
assign micromatrizz[31][205] = 9'b111111111;
assign micromatrizz[31][206] = 9'b111111111;
assign micromatrizz[31][207] = 9'b111111111;
assign micromatrizz[31][208] = 9'b111111111;
assign micromatrizz[31][209] = 9'b111111111;
assign micromatrizz[31][210] = 9'b111111111;
assign micromatrizz[31][211] = 9'b111111111;
assign micromatrizz[31][212] = 9'b111111111;
assign micromatrizz[31][213] = 9'b111111111;
assign micromatrizz[31][214] = 9'b111111111;
assign micromatrizz[31][215] = 9'b111111111;
assign micromatrizz[31][216] = 9'b111111111;
assign micromatrizz[31][217] = 9'b111111111;
assign micromatrizz[31][218] = 9'b111111111;
assign micromatrizz[31][219] = 9'b111111111;
assign micromatrizz[31][220] = 9'b111111111;
assign micromatrizz[31][221] = 9'b111111111;
assign micromatrizz[31][222] = 9'b111111111;
assign micromatrizz[31][223] = 9'b111111111;
assign micromatrizz[31][224] = 9'b111111111;
assign micromatrizz[31][225] = 9'b111111111;
assign micromatrizz[31][226] = 9'b111111111;
assign micromatrizz[31][227] = 9'b111111111;
assign micromatrizz[31][228] = 9'b111111111;
assign micromatrizz[31][229] = 9'b111111111;
assign micromatrizz[31][230] = 9'b111111111;
assign micromatrizz[31][231] = 9'b111111111;
assign micromatrizz[31][232] = 9'b111111111;
assign micromatrizz[31][233] = 9'b111111111;
assign micromatrizz[31][234] = 9'b111111111;
assign micromatrizz[31][235] = 9'b111111111;
assign micromatrizz[31][236] = 9'b111111111;
assign micromatrizz[31][237] = 9'b111111111;
assign micromatrizz[31][238] = 9'b111111111;
assign micromatrizz[31][239] = 9'b111111111;
assign micromatrizz[31][240] = 9'b111111111;
assign micromatrizz[31][241] = 9'b111111111;
assign micromatrizz[31][242] = 9'b111111111;
assign micromatrizz[31][243] = 9'b111111111;
assign micromatrizz[31][244] = 9'b111111111;
assign micromatrizz[31][245] = 9'b111111111;
assign micromatrizz[31][246] = 9'b111111111;
assign micromatrizz[31][247] = 9'b111111111;
assign micromatrizz[31][248] = 9'b111111111;
assign micromatrizz[31][249] = 9'b111111111;
assign micromatrizz[31][250] = 9'b111111111;
assign micromatrizz[31][251] = 9'b111111111;
assign micromatrizz[31][252] = 9'b111111111;
assign micromatrizz[31][253] = 9'b111111111;
assign micromatrizz[31][254] = 9'b111111111;
assign micromatrizz[31][255] = 9'b111111111;
assign micromatrizz[31][256] = 9'b111111111;
assign micromatrizz[31][257] = 9'b111111111;
assign micromatrizz[31][258] = 9'b111111111;
assign micromatrizz[31][259] = 9'b111111111;
assign micromatrizz[31][260] = 9'b111111111;
assign micromatrizz[31][261] = 9'b111111111;
assign micromatrizz[31][262] = 9'b111111111;
assign micromatrizz[31][263] = 9'b111111111;
assign micromatrizz[31][264] = 9'b111111111;
assign micromatrizz[31][265] = 9'b111111111;
assign micromatrizz[31][266] = 9'b111111111;
assign micromatrizz[31][267] = 9'b111111111;
assign micromatrizz[31][268] = 9'b111111111;
assign micromatrizz[31][269] = 9'b111111111;
assign micromatrizz[31][270] = 9'b111110010;
assign micromatrizz[31][271] = 9'b111110010;
assign micromatrizz[31][272] = 9'b111110010;
assign micromatrizz[31][273] = 9'b111110010;
assign micromatrizz[31][274] = 9'b111110010;
assign micromatrizz[31][275] = 9'b111110011;
assign micromatrizz[31][276] = 9'b111110011;
assign micromatrizz[31][277] = 9'b111110011;
assign micromatrizz[31][278] = 9'b111110011;
assign micromatrizz[31][279] = 9'b111111111;
assign micromatrizz[31][280] = 9'b111111111;
assign micromatrizz[31][281] = 9'b111111111;
assign micromatrizz[31][282] = 9'b111111111;
assign micromatrizz[31][283] = 9'b111111111;
assign micromatrizz[31][284] = 9'b111111111;
assign micromatrizz[31][285] = 9'b111111111;
assign micromatrizz[31][286] = 9'b111111111;
assign micromatrizz[31][287] = 9'b111111111;
assign micromatrizz[31][288] = 9'b111111111;
assign micromatrizz[31][289] = 9'b111111111;
assign micromatrizz[31][290] = 9'b111110010;
assign micromatrizz[31][291] = 9'b111110010;
assign micromatrizz[31][292] = 9'b111110011;
assign micromatrizz[31][293] = 9'b111110010;
assign micromatrizz[31][294] = 9'b111110011;
assign micromatrizz[31][295] = 9'b111110011;
assign micromatrizz[31][296] = 9'b111110011;
assign micromatrizz[31][297] = 9'b111110111;
assign micromatrizz[31][298] = 9'b111111111;
assign micromatrizz[31][299] = 9'b111111111;
assign micromatrizz[31][300] = 9'b111111111;
assign micromatrizz[31][301] = 9'b111111111;
assign micromatrizz[31][302] = 9'b111111111;
assign micromatrizz[31][303] = 9'b111111111;
assign micromatrizz[31][304] = 9'b111111111;
assign micromatrizz[31][305] = 9'b111110111;
assign micromatrizz[31][306] = 9'b111111111;
assign micromatrizz[31][307] = 9'b111111111;
assign micromatrizz[31][308] = 9'b111111111;
assign micromatrizz[31][309] = 9'b111111111;
assign micromatrizz[31][310] = 9'b111111111;
assign micromatrizz[31][311] = 9'b111110111;
assign micromatrizz[31][312] = 9'b111110010;
assign micromatrizz[31][313] = 9'b111110010;
assign micromatrizz[31][314] = 9'b111110010;
assign micromatrizz[31][315] = 9'b111110010;
assign micromatrizz[31][316] = 9'b111110011;
assign micromatrizz[31][317] = 9'b111110010;
assign micromatrizz[31][318] = 9'b111110011;
assign micromatrizz[31][319] = 9'b111110011;
assign micromatrizz[31][320] = 9'b111110011;
assign micromatrizz[31][321] = 9'b111111111;
assign micromatrizz[31][322] = 9'b111111111;
assign micromatrizz[31][323] = 9'b111111111;
assign micromatrizz[31][324] = 9'b111111111;
assign micromatrizz[31][325] = 9'b111111111;
assign micromatrizz[31][326] = 9'b111111111;
assign micromatrizz[31][327] = 9'b111111111;
assign micromatrizz[31][328] = 9'b111111111;
assign micromatrizz[31][329] = 9'b111111111;
assign micromatrizz[31][330] = 9'b111111111;
assign micromatrizz[31][331] = 9'b111111111;
assign micromatrizz[31][332] = 9'b111111111;
assign micromatrizz[31][333] = 9'b111111111;
assign micromatrizz[31][334] = 9'b111111111;
assign micromatrizz[31][335] = 9'b111111111;
assign micromatrizz[31][336] = 9'b111111111;
assign micromatrizz[31][337] = 9'b111111111;
assign micromatrizz[31][338] = 9'b111111111;
assign micromatrizz[31][339] = 9'b111111111;
assign micromatrizz[31][340] = 9'b111111111;
assign micromatrizz[31][341] = 9'b111111111;
assign micromatrizz[31][342] = 9'b111111111;
assign micromatrizz[31][343] = 9'b111111111;
assign micromatrizz[31][344] = 9'b111111111;
assign micromatrizz[31][345] = 9'b111111111;
assign micromatrizz[31][346] = 9'b111111111;
assign micromatrizz[31][347] = 9'b111111111;
assign micromatrizz[31][348] = 9'b111111111;
assign micromatrizz[31][349] = 9'b111111111;
assign micromatrizz[31][350] = 9'b111111111;
assign micromatrizz[31][351] = 9'b111111111;
assign micromatrizz[31][352] = 9'b111111111;
assign micromatrizz[31][353] = 9'b111111111;
assign micromatrizz[31][354] = 9'b111111111;
assign micromatrizz[31][355] = 9'b111111111;
assign micromatrizz[31][356] = 9'b111111111;
assign micromatrizz[31][357] = 9'b111111111;
assign micromatrizz[31][358] = 9'b111111111;
assign micromatrizz[31][359] = 9'b111111111;
assign micromatrizz[31][360] = 9'b111111111;
assign micromatrizz[31][361] = 9'b111111111;
assign micromatrizz[31][362] = 9'b111111111;
assign micromatrizz[31][363] = 9'b111111111;
assign micromatrizz[31][364] = 9'b111111111;
assign micromatrizz[31][365] = 9'b111111111;
assign micromatrizz[31][366] = 9'b111111111;
assign micromatrizz[31][367] = 9'b111111111;
assign micromatrizz[31][368] = 9'b111111111;
assign micromatrizz[31][369] = 9'b111111111;
assign micromatrizz[31][370] = 9'b111111111;
assign micromatrizz[31][371] = 9'b111111111;
assign micromatrizz[31][372] = 9'b111111111;
assign micromatrizz[31][373] = 9'b111111111;
assign micromatrizz[31][374] = 9'b111111111;
assign micromatrizz[31][375] = 9'b111111111;
assign micromatrizz[31][376] = 9'b111111111;
assign micromatrizz[31][377] = 9'b111111111;
assign micromatrizz[31][378] = 9'b111111111;
assign micromatrizz[31][379] = 9'b111111111;
assign micromatrizz[31][380] = 9'b111111111;
assign micromatrizz[31][381] = 9'b111111111;
assign micromatrizz[31][382] = 9'b111111111;
assign micromatrizz[31][383] = 9'b111111111;
assign micromatrizz[31][384] = 9'b111111111;
assign micromatrizz[31][385] = 9'b111111111;
assign micromatrizz[31][386] = 9'b111111111;
assign micromatrizz[31][387] = 9'b111111111;
assign micromatrizz[31][388] = 9'b111111111;
assign micromatrizz[31][389] = 9'b111111111;
assign micromatrizz[31][390] = 9'b111111111;
assign micromatrizz[31][391] = 9'b111111111;
assign micromatrizz[31][392] = 9'b111111111;
assign micromatrizz[31][393] = 9'b111111111;
assign micromatrizz[31][394] = 9'b111111111;
assign micromatrizz[31][395] = 9'b111111111;
assign micromatrizz[31][396] = 9'b111111111;
assign micromatrizz[31][397] = 9'b111111111;
assign micromatrizz[31][398] = 9'b111111111;
assign micromatrizz[31][399] = 9'b111111111;
assign micromatrizz[31][400] = 9'b111111111;
assign micromatrizz[31][401] = 9'b111111111;
assign micromatrizz[31][402] = 9'b111111111;
assign micromatrizz[31][403] = 9'b111111111;
assign micromatrizz[31][404] = 9'b111111111;
assign micromatrizz[31][405] = 9'b111111111;
assign micromatrizz[31][406] = 9'b111111111;
assign micromatrizz[31][407] = 9'b111111111;
assign micromatrizz[31][408] = 9'b111111111;
assign micromatrizz[31][409] = 9'b111111111;
assign micromatrizz[31][410] = 9'b111111111;
assign micromatrizz[31][411] = 9'b111111111;
assign micromatrizz[31][412] = 9'b111111111;
assign micromatrizz[31][413] = 9'b111111111;
assign micromatrizz[31][414] = 9'b111111111;
assign micromatrizz[31][415] = 9'b111111111;
assign micromatrizz[31][416] = 9'b111111111;
assign micromatrizz[31][417] = 9'b111111111;
assign micromatrizz[31][418] = 9'b111111111;
assign micromatrizz[31][419] = 9'b111111111;
assign micromatrizz[31][420] = 9'b111111111;
assign micromatrizz[31][421] = 9'b111111111;
assign micromatrizz[31][422] = 9'b111111111;
assign micromatrizz[31][423] = 9'b111111111;
assign micromatrizz[31][424] = 9'b111111111;
assign micromatrizz[31][425] = 9'b111111111;
assign micromatrizz[31][426] = 9'b111111111;
assign micromatrizz[31][427] = 9'b111111111;
assign micromatrizz[31][428] = 9'b111111111;
assign micromatrizz[31][429] = 9'b111111111;
assign micromatrizz[31][430] = 9'b111111111;
assign micromatrizz[31][431] = 9'b111111111;
assign micromatrizz[31][432] = 9'b111111111;
assign micromatrizz[31][433] = 9'b111111111;
assign micromatrizz[31][434] = 9'b111111111;
assign micromatrizz[31][435] = 9'b111111111;
assign micromatrizz[31][436] = 9'b111111111;
assign micromatrizz[31][437] = 9'b111111111;
assign micromatrizz[31][438] = 9'b111111111;
assign micromatrizz[31][439] = 9'b111111111;
assign micromatrizz[31][440] = 9'b111111111;
assign micromatrizz[31][441] = 9'b111111111;
assign micromatrizz[31][442] = 9'b111111111;
assign micromatrizz[31][443] = 9'b111111111;
assign micromatrizz[31][444] = 9'b111111111;
assign micromatrizz[31][445] = 9'b111111111;
assign micromatrizz[31][446] = 9'b111111111;
assign micromatrizz[31][447] = 9'b111111111;
assign micromatrizz[31][448] = 9'b111111111;
assign micromatrizz[31][449] = 9'b111111111;
assign micromatrizz[31][450] = 9'b111111111;
assign micromatrizz[31][451] = 9'b111111111;
assign micromatrizz[31][452] = 9'b111111111;
assign micromatrizz[31][453] = 9'b111111111;
assign micromatrizz[31][454] = 9'b111111111;
assign micromatrizz[31][455] = 9'b111111111;
assign micromatrizz[31][456] = 9'b111111111;
assign micromatrizz[31][457] = 9'b111111111;
assign micromatrizz[31][458] = 9'b111111111;
assign micromatrizz[31][459] = 9'b111111111;
assign micromatrizz[31][460] = 9'b111111111;
assign micromatrizz[31][461] = 9'b111111111;
assign micromatrizz[31][462] = 9'b111111111;
assign micromatrizz[31][463] = 9'b111111111;
assign micromatrizz[31][464] = 9'b111111111;
assign micromatrizz[31][465] = 9'b111111111;
assign micromatrizz[31][466] = 9'b111111111;
assign micromatrizz[31][467] = 9'b111111111;
assign micromatrizz[31][468] = 9'b111111111;
assign micromatrizz[31][469] = 9'b111111111;
assign micromatrizz[31][470] = 9'b111111111;
assign micromatrizz[31][471] = 9'b111111111;
assign micromatrizz[31][472] = 9'b111111111;
assign micromatrizz[31][473] = 9'b111111111;
assign micromatrizz[31][474] = 9'b111111111;
assign micromatrizz[31][475] = 9'b111111111;
assign micromatrizz[31][476] = 9'b111111111;
assign micromatrizz[31][477] = 9'b111111111;
assign micromatrizz[31][478] = 9'b111111111;
assign micromatrizz[31][479] = 9'b111111111;
assign micromatrizz[31][480] = 9'b111111111;
assign micromatrizz[31][481] = 9'b111111111;
assign micromatrizz[31][482] = 9'b111111111;
assign micromatrizz[31][483] = 9'b111111111;
assign micromatrizz[31][484] = 9'b111111111;
assign micromatrizz[31][485] = 9'b111111111;
assign micromatrizz[31][486] = 9'b111111111;
assign micromatrizz[31][487] = 9'b111111111;
assign micromatrizz[31][488] = 9'b111111111;
assign micromatrizz[31][489] = 9'b111111111;
assign micromatrizz[31][490] = 9'b111111111;
assign micromatrizz[31][491] = 9'b111111111;
assign micromatrizz[31][492] = 9'b111111111;
assign micromatrizz[31][493] = 9'b111111111;
assign micromatrizz[31][494] = 9'b111111111;
assign micromatrizz[31][495] = 9'b111111111;
assign micromatrizz[31][496] = 9'b111111111;
assign micromatrizz[31][497] = 9'b111111111;
assign micromatrizz[31][498] = 9'b111111111;
assign micromatrizz[31][499] = 9'b111111111;
assign micromatrizz[31][500] = 9'b111111111;
assign micromatrizz[31][501] = 9'b111111111;
assign micromatrizz[31][502] = 9'b111111111;
assign micromatrizz[31][503] = 9'b111111111;
assign micromatrizz[31][504] = 9'b111111111;
assign micromatrizz[31][505] = 9'b111111111;
assign micromatrizz[31][506] = 9'b111111111;
assign micromatrizz[31][507] = 9'b111111111;
assign micromatrizz[31][508] = 9'b111111111;
assign micromatrizz[31][509] = 9'b111111111;
assign micromatrizz[31][510] = 9'b111111111;
assign micromatrizz[31][511] = 9'b111111111;
assign micromatrizz[31][512] = 9'b111111111;
assign micromatrizz[31][513] = 9'b111111111;
assign micromatrizz[31][514] = 9'b111111111;
assign micromatrizz[31][515] = 9'b111111111;
assign micromatrizz[31][516] = 9'b111111111;
assign micromatrizz[31][517] = 9'b111111111;
assign micromatrizz[31][518] = 9'b111111111;
assign micromatrizz[31][519] = 9'b111111111;
assign micromatrizz[31][520] = 9'b111111111;
assign micromatrizz[31][521] = 9'b111111111;
assign micromatrizz[31][522] = 9'b111111111;
assign micromatrizz[31][523] = 9'b111111111;
assign micromatrizz[31][524] = 9'b111111111;
assign micromatrizz[31][525] = 9'b111111111;
assign micromatrizz[31][526] = 9'b111111111;
assign micromatrizz[31][527] = 9'b111111111;
assign micromatrizz[31][528] = 9'b111111111;
assign micromatrizz[31][529] = 9'b111111111;
assign micromatrizz[31][530] = 9'b111111111;
assign micromatrizz[31][531] = 9'b111111111;
assign micromatrizz[31][532] = 9'b111111111;
assign micromatrizz[31][533] = 9'b111111111;
assign micromatrizz[31][534] = 9'b111111111;
assign micromatrizz[31][535] = 9'b111111111;
assign micromatrizz[31][536] = 9'b111111111;
assign micromatrizz[31][537] = 9'b111111111;
assign micromatrizz[31][538] = 9'b111111111;
assign micromatrizz[31][539] = 9'b111111111;
assign micromatrizz[31][540] = 9'b111111111;
assign micromatrizz[31][541] = 9'b111111111;
assign micromatrizz[31][542] = 9'b111111111;
assign micromatrizz[31][543] = 9'b111111111;
assign micromatrizz[31][544] = 9'b111111111;
assign micromatrizz[31][545] = 9'b111111111;
assign micromatrizz[31][546] = 9'b111111111;
assign micromatrizz[31][547] = 9'b111111111;
assign micromatrizz[31][548] = 9'b111111111;
assign micromatrizz[31][549] = 9'b111111111;
assign micromatrizz[31][550] = 9'b111111111;
assign micromatrizz[31][551] = 9'b111111111;
assign micromatrizz[31][552] = 9'b111111111;
assign micromatrizz[31][553] = 9'b111111111;
assign micromatrizz[31][554] = 9'b111111111;
assign micromatrizz[31][555] = 9'b111111111;
assign micromatrizz[31][556] = 9'b111111111;
assign micromatrizz[31][557] = 9'b111111111;
assign micromatrizz[31][558] = 9'b111111111;
assign micromatrizz[31][559] = 9'b111111111;
assign micromatrizz[31][560] = 9'b111111111;
assign micromatrizz[31][561] = 9'b111111111;
assign micromatrizz[31][562] = 9'b111111111;
assign micromatrizz[31][563] = 9'b111111111;
assign micromatrizz[31][564] = 9'b111111111;
assign micromatrizz[31][565] = 9'b111111111;
assign micromatrizz[31][566] = 9'b111111111;
assign micromatrizz[31][567] = 9'b111111111;
assign micromatrizz[31][568] = 9'b111111111;
assign micromatrizz[31][569] = 9'b111111111;
assign micromatrizz[31][570] = 9'b111111111;
assign micromatrizz[31][571] = 9'b111111111;
assign micromatrizz[31][572] = 9'b111111111;
assign micromatrizz[31][573] = 9'b111111111;
assign micromatrizz[31][574] = 9'b111111111;
assign micromatrizz[31][575] = 9'b111111111;
assign micromatrizz[31][576] = 9'b111111111;
assign micromatrizz[31][577] = 9'b111111111;
assign micromatrizz[31][578] = 9'b111111111;
assign micromatrizz[31][579] = 9'b111111111;
assign micromatrizz[31][580] = 9'b111111111;
assign micromatrizz[31][581] = 9'b111111111;
assign micromatrizz[31][582] = 9'b111111111;
assign micromatrizz[31][583] = 9'b111111111;
assign micromatrizz[31][584] = 9'b111111111;
assign micromatrizz[31][585] = 9'b111111111;
assign micromatrizz[31][586] = 9'b111111111;
assign micromatrizz[31][587] = 9'b111111111;
assign micromatrizz[31][588] = 9'b111111111;
assign micromatrizz[31][589] = 9'b111111111;
assign micromatrizz[31][590] = 9'b111111111;
assign micromatrizz[31][591] = 9'b111111111;
assign micromatrizz[31][592] = 9'b111111111;
assign micromatrizz[31][593] = 9'b111111111;
assign micromatrizz[31][594] = 9'b111111111;
assign micromatrizz[31][595] = 9'b111111111;
assign micromatrizz[31][596] = 9'b111111111;
assign micromatrizz[31][597] = 9'b111111111;
assign micromatrizz[31][598] = 9'b111111111;
assign micromatrizz[31][599] = 9'b111111111;
assign micromatrizz[31][600] = 9'b111111111;
assign micromatrizz[31][601] = 9'b111111111;
assign micromatrizz[31][602] = 9'b111111111;
assign micromatrizz[31][603] = 9'b111111111;
assign micromatrizz[31][604] = 9'b111111111;
assign micromatrizz[31][605] = 9'b111111111;
assign micromatrizz[31][606] = 9'b111111111;
assign micromatrizz[31][607] = 9'b111111111;
assign micromatrizz[31][608] = 9'b111111111;
assign micromatrizz[31][609] = 9'b111111111;
assign micromatrizz[31][610] = 9'b111111111;
assign micromatrizz[31][611] = 9'b111111111;
assign micromatrizz[31][612] = 9'b111111111;
assign micromatrizz[31][613] = 9'b111111111;
assign micromatrizz[31][614] = 9'b111111111;
assign micromatrizz[31][615] = 9'b111111111;
assign micromatrizz[31][616] = 9'b111111111;
assign micromatrizz[31][617] = 9'b111111111;
assign micromatrizz[31][618] = 9'b111111111;
assign micromatrizz[31][619] = 9'b111111111;
assign micromatrizz[31][620] = 9'b111111111;
assign micromatrizz[31][621] = 9'b111111111;
assign micromatrizz[31][622] = 9'b111111111;
assign micromatrizz[31][623] = 9'b111111111;
assign micromatrizz[31][624] = 9'b111111111;
assign micromatrizz[31][625] = 9'b111111111;
assign micromatrizz[31][626] = 9'b111111111;
assign micromatrizz[31][627] = 9'b111111111;
assign micromatrizz[31][628] = 9'b111111111;
assign micromatrizz[31][629] = 9'b111111111;
assign micromatrizz[31][630] = 9'b111111111;
assign micromatrizz[31][631] = 9'b111111111;
assign micromatrizz[31][632] = 9'b111111111;
assign micromatrizz[31][633] = 9'b111111111;
assign micromatrizz[31][634] = 9'b111111111;
assign micromatrizz[31][635] = 9'b111111111;
assign micromatrizz[31][636] = 9'b111111111;
assign micromatrizz[31][637] = 9'b111111111;
assign micromatrizz[31][638] = 9'b111111111;
assign micromatrizz[31][639] = 9'b111111111;
assign micromatrizz[32][0] = 9'b111111111;
assign micromatrizz[32][1] = 9'b111111111;
assign micromatrizz[32][2] = 9'b111111111;
assign micromatrizz[32][3] = 9'b111111111;
assign micromatrizz[32][4] = 9'b111111111;
assign micromatrizz[32][5] = 9'b111111111;
assign micromatrizz[32][6] = 9'b111111111;
assign micromatrizz[32][7] = 9'b111111111;
assign micromatrizz[32][8] = 9'b111111111;
assign micromatrizz[32][9] = 9'b111111111;
assign micromatrizz[32][10] = 9'b111111111;
assign micromatrizz[32][11] = 9'b111111111;
assign micromatrizz[32][12] = 9'b111111111;
assign micromatrizz[32][13] = 9'b111111111;
assign micromatrizz[32][14] = 9'b111111111;
assign micromatrizz[32][15] = 9'b111111111;
assign micromatrizz[32][16] = 9'b111111111;
assign micromatrizz[32][17] = 9'b111111111;
assign micromatrizz[32][18] = 9'b111111111;
assign micromatrizz[32][19] = 9'b111111111;
assign micromatrizz[32][20] = 9'b111111111;
assign micromatrizz[32][21] = 9'b111111111;
assign micromatrizz[32][22] = 9'b111111111;
assign micromatrizz[32][23] = 9'b111111111;
assign micromatrizz[32][24] = 9'b111111111;
assign micromatrizz[32][25] = 9'b111111111;
assign micromatrizz[32][26] = 9'b111111111;
assign micromatrizz[32][27] = 9'b111111111;
assign micromatrizz[32][28] = 9'b111111111;
assign micromatrizz[32][29] = 9'b111111111;
assign micromatrizz[32][30] = 9'b111111111;
assign micromatrizz[32][31] = 9'b111111111;
assign micromatrizz[32][32] = 9'b111111111;
assign micromatrizz[32][33] = 9'b111111111;
assign micromatrizz[32][34] = 9'b111111111;
assign micromatrizz[32][35] = 9'b111111111;
assign micromatrizz[32][36] = 9'b111111111;
assign micromatrizz[32][37] = 9'b111111111;
assign micromatrizz[32][38] = 9'b111111111;
assign micromatrizz[32][39] = 9'b111111111;
assign micromatrizz[32][40] = 9'b111111111;
assign micromatrizz[32][41] = 9'b111111111;
assign micromatrizz[32][42] = 9'b111111111;
assign micromatrizz[32][43] = 9'b111111111;
assign micromatrizz[32][44] = 9'b111111111;
assign micromatrizz[32][45] = 9'b111111111;
assign micromatrizz[32][46] = 9'b111111111;
assign micromatrizz[32][47] = 9'b111111111;
assign micromatrizz[32][48] = 9'b111111111;
assign micromatrizz[32][49] = 9'b111111111;
assign micromatrizz[32][50] = 9'b111111111;
assign micromatrizz[32][51] = 9'b111111111;
assign micromatrizz[32][52] = 9'b111111111;
assign micromatrizz[32][53] = 9'b111111111;
assign micromatrizz[32][54] = 9'b111111111;
assign micromatrizz[32][55] = 9'b111111111;
assign micromatrizz[32][56] = 9'b111111111;
assign micromatrizz[32][57] = 9'b111111111;
assign micromatrizz[32][58] = 9'b111111111;
assign micromatrizz[32][59] = 9'b111111111;
assign micromatrizz[32][60] = 9'b111111111;
assign micromatrizz[32][61] = 9'b111111111;
assign micromatrizz[32][62] = 9'b111111111;
assign micromatrizz[32][63] = 9'b111111111;
assign micromatrizz[32][64] = 9'b111111111;
assign micromatrizz[32][65] = 9'b111111111;
assign micromatrizz[32][66] = 9'b111111111;
assign micromatrizz[32][67] = 9'b111111111;
assign micromatrizz[32][68] = 9'b111111111;
assign micromatrizz[32][69] = 9'b111111111;
assign micromatrizz[32][70] = 9'b111111111;
assign micromatrizz[32][71] = 9'b111111111;
assign micromatrizz[32][72] = 9'b111111111;
assign micromatrizz[32][73] = 9'b111111111;
assign micromatrizz[32][74] = 9'b111111111;
assign micromatrizz[32][75] = 9'b111111111;
assign micromatrizz[32][76] = 9'b111111111;
assign micromatrizz[32][77] = 9'b111111111;
assign micromatrizz[32][78] = 9'b111111111;
assign micromatrizz[32][79] = 9'b111111111;
assign micromatrizz[32][80] = 9'b111111111;
assign micromatrizz[32][81] = 9'b111111111;
assign micromatrizz[32][82] = 9'b111111111;
assign micromatrizz[32][83] = 9'b111111111;
assign micromatrizz[32][84] = 9'b111111111;
assign micromatrizz[32][85] = 9'b111111111;
assign micromatrizz[32][86] = 9'b111111111;
assign micromatrizz[32][87] = 9'b111111111;
assign micromatrizz[32][88] = 9'b111111111;
assign micromatrizz[32][89] = 9'b111111111;
assign micromatrizz[32][90] = 9'b111111111;
assign micromatrizz[32][91] = 9'b111111111;
assign micromatrizz[32][92] = 9'b111111111;
assign micromatrizz[32][93] = 9'b111111111;
assign micromatrizz[32][94] = 9'b111111111;
assign micromatrizz[32][95] = 9'b111111111;
assign micromatrizz[32][96] = 9'b111111111;
assign micromatrizz[32][97] = 9'b111111111;
assign micromatrizz[32][98] = 9'b111111111;
assign micromatrizz[32][99] = 9'b111111111;
assign micromatrizz[32][100] = 9'b111111111;
assign micromatrizz[32][101] = 9'b111111111;
assign micromatrizz[32][102] = 9'b111111111;
assign micromatrizz[32][103] = 9'b111111111;
assign micromatrizz[32][104] = 9'b111111111;
assign micromatrizz[32][105] = 9'b111111111;
assign micromatrizz[32][106] = 9'b111111111;
assign micromatrizz[32][107] = 9'b111111111;
assign micromatrizz[32][108] = 9'b111111111;
assign micromatrizz[32][109] = 9'b111111111;
assign micromatrizz[32][110] = 9'b111111111;
assign micromatrizz[32][111] = 9'b111111111;
assign micromatrizz[32][112] = 9'b111111111;
assign micromatrizz[32][113] = 9'b111111111;
assign micromatrizz[32][114] = 9'b111111111;
assign micromatrizz[32][115] = 9'b111111111;
assign micromatrizz[32][116] = 9'b111111111;
assign micromatrizz[32][117] = 9'b111111111;
assign micromatrizz[32][118] = 9'b111111111;
assign micromatrizz[32][119] = 9'b111111111;
assign micromatrizz[32][120] = 9'b111111111;
assign micromatrizz[32][121] = 9'b111111111;
assign micromatrizz[32][122] = 9'b111111111;
assign micromatrizz[32][123] = 9'b111111111;
assign micromatrizz[32][124] = 9'b111111111;
assign micromatrizz[32][125] = 9'b111111111;
assign micromatrizz[32][126] = 9'b111111111;
assign micromatrizz[32][127] = 9'b111111111;
assign micromatrizz[32][128] = 9'b111111111;
assign micromatrizz[32][129] = 9'b111111111;
assign micromatrizz[32][130] = 9'b111111111;
assign micromatrizz[32][131] = 9'b111111111;
assign micromatrizz[32][132] = 9'b111111111;
assign micromatrizz[32][133] = 9'b111111111;
assign micromatrizz[32][134] = 9'b111111111;
assign micromatrizz[32][135] = 9'b111111111;
assign micromatrizz[32][136] = 9'b111111111;
assign micromatrizz[32][137] = 9'b111111111;
assign micromatrizz[32][138] = 9'b111111111;
assign micromatrizz[32][139] = 9'b111111111;
assign micromatrizz[32][140] = 9'b111111111;
assign micromatrizz[32][141] = 9'b111111111;
assign micromatrizz[32][142] = 9'b111111111;
assign micromatrizz[32][143] = 9'b111111111;
assign micromatrizz[32][144] = 9'b111111111;
assign micromatrizz[32][145] = 9'b111111111;
assign micromatrizz[32][146] = 9'b111111111;
assign micromatrizz[32][147] = 9'b111111111;
assign micromatrizz[32][148] = 9'b111111111;
assign micromatrizz[32][149] = 9'b111111111;
assign micromatrizz[32][150] = 9'b111111111;
assign micromatrizz[32][151] = 9'b111111111;
assign micromatrizz[32][152] = 9'b111111111;
assign micromatrizz[32][153] = 9'b111111111;
assign micromatrizz[32][154] = 9'b111111111;
assign micromatrizz[32][155] = 9'b111111111;
assign micromatrizz[32][156] = 9'b111111111;
assign micromatrizz[32][157] = 9'b111111111;
assign micromatrizz[32][158] = 9'b111111111;
assign micromatrizz[32][159] = 9'b111111111;
assign micromatrizz[32][160] = 9'b111111111;
assign micromatrizz[32][161] = 9'b111111111;
assign micromatrizz[32][162] = 9'b111111111;
assign micromatrizz[32][163] = 9'b111111111;
assign micromatrizz[32][164] = 9'b111111111;
assign micromatrizz[32][165] = 9'b111111111;
assign micromatrizz[32][166] = 9'b111111111;
assign micromatrizz[32][167] = 9'b111111111;
assign micromatrizz[32][168] = 9'b111111111;
assign micromatrizz[32][169] = 9'b111111111;
assign micromatrizz[32][170] = 9'b111111111;
assign micromatrizz[32][171] = 9'b111111111;
assign micromatrizz[32][172] = 9'b111111111;
assign micromatrizz[32][173] = 9'b111111111;
assign micromatrizz[32][174] = 9'b111111111;
assign micromatrizz[32][175] = 9'b111111111;
assign micromatrizz[32][176] = 9'b111111111;
assign micromatrizz[32][177] = 9'b111111111;
assign micromatrizz[32][178] = 9'b111111111;
assign micromatrizz[32][179] = 9'b111111111;
assign micromatrizz[32][180] = 9'b111111111;
assign micromatrizz[32][181] = 9'b111111111;
assign micromatrizz[32][182] = 9'b111111111;
assign micromatrizz[32][183] = 9'b111111111;
assign micromatrizz[32][184] = 9'b111111111;
assign micromatrizz[32][185] = 9'b111111111;
assign micromatrizz[32][186] = 9'b111111111;
assign micromatrizz[32][187] = 9'b111111111;
assign micromatrizz[32][188] = 9'b111111111;
assign micromatrizz[32][189] = 9'b111111111;
assign micromatrizz[32][190] = 9'b111111111;
assign micromatrizz[32][191] = 9'b111111111;
assign micromatrizz[32][192] = 9'b111111111;
assign micromatrizz[32][193] = 9'b111111111;
assign micromatrizz[32][194] = 9'b111111111;
assign micromatrizz[32][195] = 9'b111111111;
assign micromatrizz[32][196] = 9'b111111111;
assign micromatrizz[32][197] = 9'b111111111;
assign micromatrizz[32][198] = 9'b111111111;
assign micromatrizz[32][199] = 9'b111111111;
assign micromatrizz[32][200] = 9'b111111111;
assign micromatrizz[32][201] = 9'b111111111;
assign micromatrizz[32][202] = 9'b111111111;
assign micromatrizz[32][203] = 9'b111111111;
assign micromatrizz[32][204] = 9'b111111111;
assign micromatrizz[32][205] = 9'b111111111;
assign micromatrizz[32][206] = 9'b111111111;
assign micromatrizz[32][207] = 9'b111111111;
assign micromatrizz[32][208] = 9'b111111111;
assign micromatrizz[32][209] = 9'b111111111;
assign micromatrizz[32][210] = 9'b111111111;
assign micromatrizz[32][211] = 9'b111111111;
assign micromatrizz[32][212] = 9'b111111111;
assign micromatrizz[32][213] = 9'b111111111;
assign micromatrizz[32][214] = 9'b111111111;
assign micromatrizz[32][215] = 9'b111111111;
assign micromatrizz[32][216] = 9'b111111111;
assign micromatrizz[32][217] = 9'b111111111;
assign micromatrizz[32][218] = 9'b111111111;
assign micromatrizz[32][219] = 9'b111111111;
assign micromatrizz[32][220] = 9'b111111111;
assign micromatrizz[32][221] = 9'b111111111;
assign micromatrizz[32][222] = 9'b111111111;
assign micromatrizz[32][223] = 9'b111111111;
assign micromatrizz[32][224] = 9'b111111111;
assign micromatrizz[32][225] = 9'b111111111;
assign micromatrizz[32][226] = 9'b111111111;
assign micromatrizz[32][227] = 9'b111111111;
assign micromatrizz[32][228] = 9'b111111111;
assign micromatrizz[32][229] = 9'b111111111;
assign micromatrizz[32][230] = 9'b111111111;
assign micromatrizz[32][231] = 9'b111111111;
assign micromatrizz[32][232] = 9'b111111111;
assign micromatrizz[32][233] = 9'b111111111;
assign micromatrizz[32][234] = 9'b111111111;
assign micromatrizz[32][235] = 9'b111111111;
assign micromatrizz[32][236] = 9'b111111111;
assign micromatrizz[32][237] = 9'b111111111;
assign micromatrizz[32][238] = 9'b111111111;
assign micromatrizz[32][239] = 9'b111111111;
assign micromatrizz[32][240] = 9'b111111111;
assign micromatrizz[32][241] = 9'b111111111;
assign micromatrizz[32][242] = 9'b111111111;
assign micromatrizz[32][243] = 9'b111111111;
assign micromatrizz[32][244] = 9'b111111111;
assign micromatrizz[32][245] = 9'b111111111;
assign micromatrizz[32][246] = 9'b111111111;
assign micromatrizz[32][247] = 9'b111111111;
assign micromatrizz[32][248] = 9'b111111111;
assign micromatrizz[32][249] = 9'b111111111;
assign micromatrizz[32][250] = 9'b111111111;
assign micromatrizz[32][251] = 9'b111111111;
assign micromatrizz[32][252] = 9'b111111111;
assign micromatrizz[32][253] = 9'b111111111;
assign micromatrizz[32][254] = 9'b111111111;
assign micromatrizz[32][255] = 9'b111111111;
assign micromatrizz[32][256] = 9'b111111111;
assign micromatrizz[32][257] = 9'b111111111;
assign micromatrizz[32][258] = 9'b111111111;
assign micromatrizz[32][259] = 9'b111111111;
assign micromatrizz[32][260] = 9'b111111111;
assign micromatrizz[32][261] = 9'b111111111;
assign micromatrizz[32][262] = 9'b111111111;
assign micromatrizz[32][263] = 9'b111111111;
assign micromatrizz[32][264] = 9'b111111111;
assign micromatrizz[32][265] = 9'b111111111;
assign micromatrizz[32][266] = 9'b111111111;
assign micromatrizz[32][267] = 9'b111111111;
assign micromatrizz[32][268] = 9'b111111111;
assign micromatrizz[32][269] = 9'b111111111;
assign micromatrizz[32][270] = 9'b111110010;
assign micromatrizz[32][271] = 9'b111110010;
assign micromatrizz[32][272] = 9'b111110010;
assign micromatrizz[32][273] = 9'b111110010;
assign micromatrizz[32][274] = 9'b111110010;
assign micromatrizz[32][275] = 9'b111110011;
assign micromatrizz[32][276] = 9'b111110011;
assign micromatrizz[32][277] = 9'b111110011;
assign micromatrizz[32][278] = 9'b111110011;
assign micromatrizz[32][279] = 9'b111111111;
assign micromatrizz[32][280] = 9'b111111111;
assign micromatrizz[32][281] = 9'b111111111;
assign micromatrizz[32][282] = 9'b111111111;
assign micromatrizz[32][283] = 9'b111111111;
assign micromatrizz[32][284] = 9'b111111111;
assign micromatrizz[32][285] = 9'b111111111;
assign micromatrizz[32][286] = 9'b111111111;
assign micromatrizz[32][287] = 9'b111111111;
assign micromatrizz[32][288] = 9'b111111111;
assign micromatrizz[32][289] = 9'b111111111;
assign micromatrizz[32][290] = 9'b111110110;
assign micromatrizz[32][291] = 9'b111110010;
assign micromatrizz[32][292] = 9'b111110011;
assign micromatrizz[32][293] = 9'b111110010;
assign micromatrizz[32][294] = 9'b111110011;
assign micromatrizz[32][295] = 9'b111110011;
assign micromatrizz[32][296] = 9'b111110011;
assign micromatrizz[32][297] = 9'b111110111;
assign micromatrizz[32][298] = 9'b111111111;
assign micromatrizz[32][299] = 9'b111111111;
assign micromatrizz[32][300] = 9'b111111111;
assign micromatrizz[32][301] = 9'b111111111;
assign micromatrizz[32][302] = 9'b111111111;
assign micromatrizz[32][303] = 9'b111111111;
assign micromatrizz[32][304] = 9'b111111111;
assign micromatrizz[32][305] = 9'b111110010;
assign micromatrizz[32][306] = 9'b111111111;
assign micromatrizz[32][307] = 9'b111111111;
assign micromatrizz[32][308] = 9'b111111111;
assign micromatrizz[32][309] = 9'b111111111;
assign micromatrizz[32][310] = 9'b111111111;
assign micromatrizz[32][311] = 9'b111111111;
assign micromatrizz[32][312] = 9'b111110110;
assign micromatrizz[32][313] = 9'b111110010;
assign micromatrizz[32][314] = 9'b111110010;
assign micromatrizz[32][315] = 9'b111110010;
assign micromatrizz[32][316] = 9'b111110010;
assign micromatrizz[32][317] = 9'b111110010;
assign micromatrizz[32][318] = 9'b111110010;
assign micromatrizz[32][319] = 9'b111110011;
assign micromatrizz[32][320] = 9'b111110010;
assign micromatrizz[32][321] = 9'b111111111;
assign micromatrizz[32][322] = 9'b111111111;
assign micromatrizz[32][323] = 9'b111111111;
assign micromatrizz[32][324] = 9'b111111111;
assign micromatrizz[32][325] = 9'b111111111;
assign micromatrizz[32][326] = 9'b111111111;
assign micromatrizz[32][327] = 9'b111111111;
assign micromatrizz[32][328] = 9'b111111111;
assign micromatrizz[32][329] = 9'b111111111;
assign micromatrizz[32][330] = 9'b111111111;
assign micromatrizz[32][331] = 9'b111111111;
assign micromatrizz[32][332] = 9'b111111111;
assign micromatrizz[32][333] = 9'b111111111;
assign micromatrizz[32][334] = 9'b111111111;
assign micromatrizz[32][335] = 9'b111111111;
assign micromatrizz[32][336] = 9'b111111111;
assign micromatrizz[32][337] = 9'b111111111;
assign micromatrizz[32][338] = 9'b111111111;
assign micromatrizz[32][339] = 9'b111111111;
assign micromatrizz[32][340] = 9'b111111111;
assign micromatrizz[32][341] = 9'b111111111;
assign micromatrizz[32][342] = 9'b111111111;
assign micromatrizz[32][343] = 9'b111111111;
assign micromatrizz[32][344] = 9'b111111111;
assign micromatrizz[32][345] = 9'b111111111;
assign micromatrizz[32][346] = 9'b111111111;
assign micromatrizz[32][347] = 9'b111111111;
assign micromatrizz[32][348] = 9'b111111111;
assign micromatrizz[32][349] = 9'b111111111;
assign micromatrizz[32][350] = 9'b111111111;
assign micromatrizz[32][351] = 9'b111111111;
assign micromatrizz[32][352] = 9'b111111111;
assign micromatrizz[32][353] = 9'b111111111;
assign micromatrizz[32][354] = 9'b111111111;
assign micromatrizz[32][355] = 9'b111111111;
assign micromatrizz[32][356] = 9'b111111111;
assign micromatrizz[32][357] = 9'b111111111;
assign micromatrizz[32][358] = 9'b111111111;
assign micromatrizz[32][359] = 9'b111111111;
assign micromatrizz[32][360] = 9'b111111111;
assign micromatrizz[32][361] = 9'b111111111;
assign micromatrizz[32][362] = 9'b111111111;
assign micromatrizz[32][363] = 9'b111111111;
assign micromatrizz[32][364] = 9'b111111111;
assign micromatrizz[32][365] = 9'b111111111;
assign micromatrizz[32][366] = 9'b111111111;
assign micromatrizz[32][367] = 9'b111111111;
assign micromatrizz[32][368] = 9'b111111111;
assign micromatrizz[32][369] = 9'b111111111;
assign micromatrizz[32][370] = 9'b111111111;
assign micromatrizz[32][371] = 9'b111111111;
assign micromatrizz[32][372] = 9'b111111111;
assign micromatrizz[32][373] = 9'b111111111;
assign micromatrizz[32][374] = 9'b111111111;
assign micromatrizz[32][375] = 9'b111111111;
assign micromatrizz[32][376] = 9'b111111111;
assign micromatrizz[32][377] = 9'b111111111;
assign micromatrizz[32][378] = 9'b111111111;
assign micromatrizz[32][379] = 9'b111111111;
assign micromatrizz[32][380] = 9'b111111111;
assign micromatrizz[32][381] = 9'b111111111;
assign micromatrizz[32][382] = 9'b111111111;
assign micromatrizz[32][383] = 9'b111111111;
assign micromatrizz[32][384] = 9'b111111111;
assign micromatrizz[32][385] = 9'b111111111;
assign micromatrizz[32][386] = 9'b111111111;
assign micromatrizz[32][387] = 9'b111111111;
assign micromatrizz[32][388] = 9'b111111111;
assign micromatrizz[32][389] = 9'b111111111;
assign micromatrizz[32][390] = 9'b111111111;
assign micromatrizz[32][391] = 9'b111111111;
assign micromatrizz[32][392] = 9'b111111111;
assign micromatrizz[32][393] = 9'b111111111;
assign micromatrizz[32][394] = 9'b111111111;
assign micromatrizz[32][395] = 9'b111111111;
assign micromatrizz[32][396] = 9'b111111111;
assign micromatrizz[32][397] = 9'b111111111;
assign micromatrizz[32][398] = 9'b111111111;
assign micromatrizz[32][399] = 9'b111111111;
assign micromatrizz[32][400] = 9'b111111111;
assign micromatrizz[32][401] = 9'b111111111;
assign micromatrizz[32][402] = 9'b111111111;
assign micromatrizz[32][403] = 9'b111111111;
assign micromatrizz[32][404] = 9'b111111111;
assign micromatrizz[32][405] = 9'b111111111;
assign micromatrizz[32][406] = 9'b111111111;
assign micromatrizz[32][407] = 9'b111111111;
assign micromatrizz[32][408] = 9'b111111111;
assign micromatrizz[32][409] = 9'b111111111;
assign micromatrizz[32][410] = 9'b111111111;
assign micromatrizz[32][411] = 9'b111111111;
assign micromatrizz[32][412] = 9'b111111111;
assign micromatrizz[32][413] = 9'b111111111;
assign micromatrizz[32][414] = 9'b111111111;
assign micromatrizz[32][415] = 9'b111111111;
assign micromatrizz[32][416] = 9'b111111111;
assign micromatrizz[32][417] = 9'b111111111;
assign micromatrizz[32][418] = 9'b111111111;
assign micromatrizz[32][419] = 9'b111111111;
assign micromatrizz[32][420] = 9'b111111111;
assign micromatrizz[32][421] = 9'b111111111;
assign micromatrizz[32][422] = 9'b111111111;
assign micromatrizz[32][423] = 9'b111111111;
assign micromatrizz[32][424] = 9'b111111111;
assign micromatrizz[32][425] = 9'b111111111;
assign micromatrizz[32][426] = 9'b111111111;
assign micromatrizz[32][427] = 9'b111111111;
assign micromatrizz[32][428] = 9'b111111111;
assign micromatrizz[32][429] = 9'b111111111;
assign micromatrizz[32][430] = 9'b111111111;
assign micromatrizz[32][431] = 9'b111111111;
assign micromatrizz[32][432] = 9'b111111111;
assign micromatrizz[32][433] = 9'b111111111;
assign micromatrizz[32][434] = 9'b111111111;
assign micromatrizz[32][435] = 9'b111111111;
assign micromatrizz[32][436] = 9'b111111111;
assign micromatrizz[32][437] = 9'b111111111;
assign micromatrizz[32][438] = 9'b111111111;
assign micromatrizz[32][439] = 9'b111111111;
assign micromatrizz[32][440] = 9'b111111111;
assign micromatrizz[32][441] = 9'b111111111;
assign micromatrizz[32][442] = 9'b111111111;
assign micromatrizz[32][443] = 9'b111111111;
assign micromatrizz[32][444] = 9'b111111111;
assign micromatrizz[32][445] = 9'b111111111;
assign micromatrizz[32][446] = 9'b111111111;
assign micromatrizz[32][447] = 9'b111111111;
assign micromatrizz[32][448] = 9'b111111111;
assign micromatrizz[32][449] = 9'b111111111;
assign micromatrizz[32][450] = 9'b111111111;
assign micromatrizz[32][451] = 9'b111111111;
assign micromatrizz[32][452] = 9'b111111111;
assign micromatrizz[32][453] = 9'b111111111;
assign micromatrizz[32][454] = 9'b111111111;
assign micromatrizz[32][455] = 9'b111111111;
assign micromatrizz[32][456] = 9'b111111111;
assign micromatrizz[32][457] = 9'b111111111;
assign micromatrizz[32][458] = 9'b111111111;
assign micromatrizz[32][459] = 9'b111111111;
assign micromatrizz[32][460] = 9'b111111111;
assign micromatrizz[32][461] = 9'b111111111;
assign micromatrizz[32][462] = 9'b111111111;
assign micromatrizz[32][463] = 9'b111111111;
assign micromatrizz[32][464] = 9'b111111111;
assign micromatrizz[32][465] = 9'b111111111;
assign micromatrizz[32][466] = 9'b111111111;
assign micromatrizz[32][467] = 9'b111111111;
assign micromatrizz[32][468] = 9'b111111111;
assign micromatrizz[32][469] = 9'b111111111;
assign micromatrizz[32][470] = 9'b111111111;
assign micromatrizz[32][471] = 9'b111111111;
assign micromatrizz[32][472] = 9'b111111111;
assign micromatrizz[32][473] = 9'b111111111;
assign micromatrizz[32][474] = 9'b111111111;
assign micromatrizz[32][475] = 9'b111111111;
assign micromatrizz[32][476] = 9'b111111111;
assign micromatrizz[32][477] = 9'b111111111;
assign micromatrizz[32][478] = 9'b111111111;
assign micromatrizz[32][479] = 9'b111111111;
assign micromatrizz[32][480] = 9'b111111111;
assign micromatrizz[32][481] = 9'b111111111;
assign micromatrizz[32][482] = 9'b111111111;
assign micromatrizz[32][483] = 9'b111111111;
assign micromatrizz[32][484] = 9'b111111111;
assign micromatrizz[32][485] = 9'b111111111;
assign micromatrizz[32][486] = 9'b111111111;
assign micromatrizz[32][487] = 9'b111111111;
assign micromatrizz[32][488] = 9'b111111111;
assign micromatrizz[32][489] = 9'b111111111;
assign micromatrizz[32][490] = 9'b111111111;
assign micromatrizz[32][491] = 9'b111111111;
assign micromatrizz[32][492] = 9'b111111111;
assign micromatrizz[32][493] = 9'b111111111;
assign micromatrizz[32][494] = 9'b111111111;
assign micromatrizz[32][495] = 9'b111111111;
assign micromatrizz[32][496] = 9'b111111111;
assign micromatrizz[32][497] = 9'b111111111;
assign micromatrizz[32][498] = 9'b111111111;
assign micromatrizz[32][499] = 9'b111111111;
assign micromatrizz[32][500] = 9'b111111111;
assign micromatrizz[32][501] = 9'b111111111;
assign micromatrizz[32][502] = 9'b111111111;
assign micromatrizz[32][503] = 9'b111111111;
assign micromatrizz[32][504] = 9'b111111111;
assign micromatrizz[32][505] = 9'b111111111;
assign micromatrizz[32][506] = 9'b111111111;
assign micromatrizz[32][507] = 9'b111111111;
assign micromatrizz[32][508] = 9'b111111111;
assign micromatrizz[32][509] = 9'b111111111;
assign micromatrizz[32][510] = 9'b111111111;
assign micromatrizz[32][511] = 9'b111111111;
assign micromatrizz[32][512] = 9'b111111111;
assign micromatrizz[32][513] = 9'b111111111;
assign micromatrizz[32][514] = 9'b111111111;
assign micromatrizz[32][515] = 9'b111111111;
assign micromatrizz[32][516] = 9'b111111111;
assign micromatrizz[32][517] = 9'b111111111;
assign micromatrizz[32][518] = 9'b111111111;
assign micromatrizz[32][519] = 9'b111111111;
assign micromatrizz[32][520] = 9'b111111111;
assign micromatrizz[32][521] = 9'b111111111;
assign micromatrizz[32][522] = 9'b111111111;
assign micromatrizz[32][523] = 9'b111111111;
assign micromatrizz[32][524] = 9'b111111111;
assign micromatrizz[32][525] = 9'b111111111;
assign micromatrizz[32][526] = 9'b111111111;
assign micromatrizz[32][527] = 9'b111111111;
assign micromatrizz[32][528] = 9'b111111111;
assign micromatrizz[32][529] = 9'b111111111;
assign micromatrizz[32][530] = 9'b111111111;
assign micromatrizz[32][531] = 9'b111111111;
assign micromatrizz[32][532] = 9'b111111111;
assign micromatrizz[32][533] = 9'b111111111;
assign micromatrizz[32][534] = 9'b111111111;
assign micromatrizz[32][535] = 9'b111111111;
assign micromatrizz[32][536] = 9'b111111111;
assign micromatrizz[32][537] = 9'b111111111;
assign micromatrizz[32][538] = 9'b111111111;
assign micromatrizz[32][539] = 9'b111111111;
assign micromatrizz[32][540] = 9'b111111111;
assign micromatrizz[32][541] = 9'b111111111;
assign micromatrizz[32][542] = 9'b111111111;
assign micromatrizz[32][543] = 9'b111111111;
assign micromatrizz[32][544] = 9'b111111111;
assign micromatrizz[32][545] = 9'b111111111;
assign micromatrizz[32][546] = 9'b111111111;
assign micromatrizz[32][547] = 9'b111111111;
assign micromatrizz[32][548] = 9'b111111111;
assign micromatrizz[32][549] = 9'b111111111;
assign micromatrizz[32][550] = 9'b111111111;
assign micromatrizz[32][551] = 9'b111111111;
assign micromatrizz[32][552] = 9'b111111111;
assign micromatrizz[32][553] = 9'b111111111;
assign micromatrizz[32][554] = 9'b111111111;
assign micromatrizz[32][555] = 9'b111111111;
assign micromatrizz[32][556] = 9'b111111111;
assign micromatrizz[32][557] = 9'b111111111;
assign micromatrizz[32][558] = 9'b111111111;
assign micromatrizz[32][559] = 9'b111111111;
assign micromatrizz[32][560] = 9'b111111111;
assign micromatrizz[32][561] = 9'b111111111;
assign micromatrizz[32][562] = 9'b111111111;
assign micromatrizz[32][563] = 9'b111111111;
assign micromatrizz[32][564] = 9'b111111111;
assign micromatrizz[32][565] = 9'b111111111;
assign micromatrizz[32][566] = 9'b111111111;
assign micromatrizz[32][567] = 9'b111111111;
assign micromatrizz[32][568] = 9'b111111111;
assign micromatrizz[32][569] = 9'b111111111;
assign micromatrizz[32][570] = 9'b111111111;
assign micromatrizz[32][571] = 9'b111111111;
assign micromatrizz[32][572] = 9'b111111111;
assign micromatrizz[32][573] = 9'b111111111;
assign micromatrizz[32][574] = 9'b111111111;
assign micromatrizz[32][575] = 9'b111111111;
assign micromatrizz[32][576] = 9'b111111111;
assign micromatrizz[32][577] = 9'b111111111;
assign micromatrizz[32][578] = 9'b111111111;
assign micromatrizz[32][579] = 9'b111111111;
assign micromatrizz[32][580] = 9'b111111111;
assign micromatrizz[32][581] = 9'b111111111;
assign micromatrizz[32][582] = 9'b111111111;
assign micromatrizz[32][583] = 9'b111111111;
assign micromatrizz[32][584] = 9'b111111111;
assign micromatrizz[32][585] = 9'b111111111;
assign micromatrizz[32][586] = 9'b111111111;
assign micromatrizz[32][587] = 9'b111111111;
assign micromatrizz[32][588] = 9'b111111111;
assign micromatrizz[32][589] = 9'b111111111;
assign micromatrizz[32][590] = 9'b111111111;
assign micromatrizz[32][591] = 9'b111111111;
assign micromatrizz[32][592] = 9'b111111111;
assign micromatrizz[32][593] = 9'b111111111;
assign micromatrizz[32][594] = 9'b111111111;
assign micromatrizz[32][595] = 9'b111111111;
assign micromatrizz[32][596] = 9'b111111111;
assign micromatrizz[32][597] = 9'b111111111;
assign micromatrizz[32][598] = 9'b111111111;
assign micromatrizz[32][599] = 9'b111111111;
assign micromatrizz[32][600] = 9'b111111111;
assign micromatrizz[32][601] = 9'b111111111;
assign micromatrizz[32][602] = 9'b111111111;
assign micromatrizz[32][603] = 9'b111111111;
assign micromatrizz[32][604] = 9'b111111111;
assign micromatrizz[32][605] = 9'b111111111;
assign micromatrizz[32][606] = 9'b111111111;
assign micromatrizz[32][607] = 9'b111111111;
assign micromatrizz[32][608] = 9'b111111111;
assign micromatrizz[32][609] = 9'b111111111;
assign micromatrizz[32][610] = 9'b111111111;
assign micromatrizz[32][611] = 9'b111111111;
assign micromatrizz[32][612] = 9'b111111111;
assign micromatrizz[32][613] = 9'b111111111;
assign micromatrizz[32][614] = 9'b111111111;
assign micromatrizz[32][615] = 9'b111111111;
assign micromatrizz[32][616] = 9'b111111111;
assign micromatrizz[32][617] = 9'b111111111;
assign micromatrizz[32][618] = 9'b111111111;
assign micromatrizz[32][619] = 9'b111111111;
assign micromatrizz[32][620] = 9'b111111111;
assign micromatrizz[32][621] = 9'b111111111;
assign micromatrizz[32][622] = 9'b111111111;
assign micromatrizz[32][623] = 9'b111111111;
assign micromatrizz[32][624] = 9'b111111111;
assign micromatrizz[32][625] = 9'b111111111;
assign micromatrizz[32][626] = 9'b111111111;
assign micromatrizz[32][627] = 9'b111111111;
assign micromatrizz[32][628] = 9'b111111111;
assign micromatrizz[32][629] = 9'b111111111;
assign micromatrizz[32][630] = 9'b111111111;
assign micromatrizz[32][631] = 9'b111111111;
assign micromatrizz[32][632] = 9'b111111111;
assign micromatrizz[32][633] = 9'b111111111;
assign micromatrizz[32][634] = 9'b111111111;
assign micromatrizz[32][635] = 9'b111111111;
assign micromatrizz[32][636] = 9'b111111111;
assign micromatrizz[32][637] = 9'b111111111;
assign micromatrizz[32][638] = 9'b111111111;
assign micromatrizz[32][639] = 9'b111111111;
assign micromatrizz[33][0] = 9'b111111111;
assign micromatrizz[33][1] = 9'b111111111;
assign micromatrizz[33][2] = 9'b111111111;
assign micromatrizz[33][3] = 9'b111111111;
assign micromatrizz[33][4] = 9'b111111111;
assign micromatrizz[33][5] = 9'b111111111;
assign micromatrizz[33][6] = 9'b111111111;
assign micromatrizz[33][7] = 9'b111111111;
assign micromatrizz[33][8] = 9'b111111111;
assign micromatrizz[33][9] = 9'b111111111;
assign micromatrizz[33][10] = 9'b111111111;
assign micromatrizz[33][11] = 9'b111111111;
assign micromatrizz[33][12] = 9'b111111111;
assign micromatrizz[33][13] = 9'b111111111;
assign micromatrizz[33][14] = 9'b111111111;
assign micromatrizz[33][15] = 9'b111111111;
assign micromatrizz[33][16] = 9'b111111111;
assign micromatrizz[33][17] = 9'b111111111;
assign micromatrizz[33][18] = 9'b111111111;
assign micromatrizz[33][19] = 9'b111111111;
assign micromatrizz[33][20] = 9'b111111111;
assign micromatrizz[33][21] = 9'b111111111;
assign micromatrizz[33][22] = 9'b111111111;
assign micromatrizz[33][23] = 9'b111111111;
assign micromatrizz[33][24] = 9'b111111111;
assign micromatrizz[33][25] = 9'b111111111;
assign micromatrizz[33][26] = 9'b111111111;
assign micromatrizz[33][27] = 9'b111111111;
assign micromatrizz[33][28] = 9'b111111111;
assign micromatrizz[33][29] = 9'b111111111;
assign micromatrizz[33][30] = 9'b111111111;
assign micromatrizz[33][31] = 9'b111111111;
assign micromatrizz[33][32] = 9'b111111111;
assign micromatrizz[33][33] = 9'b111111111;
assign micromatrizz[33][34] = 9'b111111111;
assign micromatrizz[33][35] = 9'b111111111;
assign micromatrizz[33][36] = 9'b111111111;
assign micromatrizz[33][37] = 9'b111111111;
assign micromatrizz[33][38] = 9'b111111111;
assign micromatrizz[33][39] = 9'b111111111;
assign micromatrizz[33][40] = 9'b111111111;
assign micromatrizz[33][41] = 9'b111111111;
assign micromatrizz[33][42] = 9'b111111111;
assign micromatrizz[33][43] = 9'b111111111;
assign micromatrizz[33][44] = 9'b111111111;
assign micromatrizz[33][45] = 9'b111111111;
assign micromatrizz[33][46] = 9'b111111111;
assign micromatrizz[33][47] = 9'b111111111;
assign micromatrizz[33][48] = 9'b111111111;
assign micromatrizz[33][49] = 9'b111111111;
assign micromatrizz[33][50] = 9'b111111111;
assign micromatrizz[33][51] = 9'b111111111;
assign micromatrizz[33][52] = 9'b111111111;
assign micromatrizz[33][53] = 9'b111111111;
assign micromatrizz[33][54] = 9'b111111111;
assign micromatrizz[33][55] = 9'b111111111;
assign micromatrizz[33][56] = 9'b111111111;
assign micromatrizz[33][57] = 9'b111111111;
assign micromatrizz[33][58] = 9'b111111111;
assign micromatrizz[33][59] = 9'b111111111;
assign micromatrizz[33][60] = 9'b111111111;
assign micromatrizz[33][61] = 9'b111111111;
assign micromatrizz[33][62] = 9'b111111111;
assign micromatrizz[33][63] = 9'b111111111;
assign micromatrizz[33][64] = 9'b111111111;
assign micromatrizz[33][65] = 9'b111111111;
assign micromatrizz[33][66] = 9'b111111111;
assign micromatrizz[33][67] = 9'b111111111;
assign micromatrizz[33][68] = 9'b111111111;
assign micromatrizz[33][69] = 9'b111111111;
assign micromatrizz[33][70] = 9'b111111111;
assign micromatrizz[33][71] = 9'b111111111;
assign micromatrizz[33][72] = 9'b111111111;
assign micromatrizz[33][73] = 9'b111111111;
assign micromatrizz[33][74] = 9'b111111111;
assign micromatrizz[33][75] = 9'b111111111;
assign micromatrizz[33][76] = 9'b111111111;
assign micromatrizz[33][77] = 9'b111111111;
assign micromatrizz[33][78] = 9'b111111111;
assign micromatrizz[33][79] = 9'b111111111;
assign micromatrizz[33][80] = 9'b111111111;
assign micromatrizz[33][81] = 9'b111111111;
assign micromatrizz[33][82] = 9'b111111111;
assign micromatrizz[33][83] = 9'b111111111;
assign micromatrizz[33][84] = 9'b111111111;
assign micromatrizz[33][85] = 9'b111111111;
assign micromatrizz[33][86] = 9'b111111111;
assign micromatrizz[33][87] = 9'b111111111;
assign micromatrizz[33][88] = 9'b111111111;
assign micromatrizz[33][89] = 9'b111111111;
assign micromatrizz[33][90] = 9'b111111111;
assign micromatrizz[33][91] = 9'b111111111;
assign micromatrizz[33][92] = 9'b111111111;
assign micromatrizz[33][93] = 9'b111111111;
assign micromatrizz[33][94] = 9'b111111111;
assign micromatrizz[33][95] = 9'b111111111;
assign micromatrizz[33][96] = 9'b111111111;
assign micromatrizz[33][97] = 9'b111111111;
assign micromatrizz[33][98] = 9'b111111111;
assign micromatrizz[33][99] = 9'b111111111;
assign micromatrizz[33][100] = 9'b111111111;
assign micromatrizz[33][101] = 9'b111111111;
assign micromatrizz[33][102] = 9'b111111111;
assign micromatrizz[33][103] = 9'b111111111;
assign micromatrizz[33][104] = 9'b111111111;
assign micromatrizz[33][105] = 9'b111111111;
assign micromatrizz[33][106] = 9'b111111111;
assign micromatrizz[33][107] = 9'b111111111;
assign micromatrizz[33][108] = 9'b111111111;
assign micromatrizz[33][109] = 9'b111111111;
assign micromatrizz[33][110] = 9'b111111111;
assign micromatrizz[33][111] = 9'b111111111;
assign micromatrizz[33][112] = 9'b111111111;
assign micromatrizz[33][113] = 9'b111111111;
assign micromatrizz[33][114] = 9'b111111111;
assign micromatrizz[33][115] = 9'b111111111;
assign micromatrizz[33][116] = 9'b111111111;
assign micromatrizz[33][117] = 9'b111111111;
assign micromatrizz[33][118] = 9'b111111111;
assign micromatrizz[33][119] = 9'b111111111;
assign micromatrizz[33][120] = 9'b111111111;
assign micromatrizz[33][121] = 9'b111111111;
assign micromatrizz[33][122] = 9'b111111111;
assign micromatrizz[33][123] = 9'b111111111;
assign micromatrizz[33][124] = 9'b111111111;
assign micromatrizz[33][125] = 9'b111111111;
assign micromatrizz[33][126] = 9'b111111111;
assign micromatrizz[33][127] = 9'b111111111;
assign micromatrizz[33][128] = 9'b111111111;
assign micromatrizz[33][129] = 9'b111111111;
assign micromatrizz[33][130] = 9'b111111111;
assign micromatrizz[33][131] = 9'b111111111;
assign micromatrizz[33][132] = 9'b111111111;
assign micromatrizz[33][133] = 9'b111111111;
assign micromatrizz[33][134] = 9'b111111111;
assign micromatrizz[33][135] = 9'b111111111;
assign micromatrizz[33][136] = 9'b111111111;
assign micromatrizz[33][137] = 9'b111111111;
assign micromatrizz[33][138] = 9'b111111111;
assign micromatrizz[33][139] = 9'b111111111;
assign micromatrizz[33][140] = 9'b111111111;
assign micromatrizz[33][141] = 9'b111111111;
assign micromatrizz[33][142] = 9'b111111111;
assign micromatrizz[33][143] = 9'b111111111;
assign micromatrizz[33][144] = 9'b111111111;
assign micromatrizz[33][145] = 9'b111111111;
assign micromatrizz[33][146] = 9'b111111111;
assign micromatrizz[33][147] = 9'b111111111;
assign micromatrizz[33][148] = 9'b111111111;
assign micromatrizz[33][149] = 9'b111111111;
assign micromatrizz[33][150] = 9'b111111111;
assign micromatrizz[33][151] = 9'b111111111;
assign micromatrizz[33][152] = 9'b111111111;
assign micromatrizz[33][153] = 9'b111111111;
assign micromatrizz[33][154] = 9'b111111111;
assign micromatrizz[33][155] = 9'b111111111;
assign micromatrizz[33][156] = 9'b111111111;
assign micromatrizz[33][157] = 9'b111111111;
assign micromatrizz[33][158] = 9'b111111111;
assign micromatrizz[33][159] = 9'b111111111;
assign micromatrizz[33][160] = 9'b111111111;
assign micromatrizz[33][161] = 9'b111111111;
assign micromatrizz[33][162] = 9'b111111111;
assign micromatrizz[33][163] = 9'b111111111;
assign micromatrizz[33][164] = 9'b111111111;
assign micromatrizz[33][165] = 9'b111111111;
assign micromatrizz[33][166] = 9'b111111111;
assign micromatrizz[33][167] = 9'b111111111;
assign micromatrizz[33][168] = 9'b111111111;
assign micromatrizz[33][169] = 9'b111111111;
assign micromatrizz[33][170] = 9'b111111111;
assign micromatrizz[33][171] = 9'b111111111;
assign micromatrizz[33][172] = 9'b111111111;
assign micromatrizz[33][173] = 9'b111111111;
assign micromatrizz[33][174] = 9'b111111111;
assign micromatrizz[33][175] = 9'b111111111;
assign micromatrizz[33][176] = 9'b111111111;
assign micromatrizz[33][177] = 9'b111111111;
assign micromatrizz[33][178] = 9'b111111111;
assign micromatrizz[33][179] = 9'b111111111;
assign micromatrizz[33][180] = 9'b111111111;
assign micromatrizz[33][181] = 9'b111111111;
assign micromatrizz[33][182] = 9'b111111111;
assign micromatrizz[33][183] = 9'b111111111;
assign micromatrizz[33][184] = 9'b111111111;
assign micromatrizz[33][185] = 9'b111111111;
assign micromatrizz[33][186] = 9'b111111111;
assign micromatrizz[33][187] = 9'b111111111;
assign micromatrizz[33][188] = 9'b111111111;
assign micromatrizz[33][189] = 9'b111111111;
assign micromatrizz[33][190] = 9'b111111111;
assign micromatrizz[33][191] = 9'b111111111;
assign micromatrizz[33][192] = 9'b111111111;
assign micromatrizz[33][193] = 9'b111111111;
assign micromatrizz[33][194] = 9'b111111111;
assign micromatrizz[33][195] = 9'b111111111;
assign micromatrizz[33][196] = 9'b111111111;
assign micromatrizz[33][197] = 9'b111111111;
assign micromatrizz[33][198] = 9'b111111111;
assign micromatrizz[33][199] = 9'b111111111;
assign micromatrizz[33][200] = 9'b111111111;
assign micromatrizz[33][201] = 9'b111111111;
assign micromatrizz[33][202] = 9'b111111111;
assign micromatrizz[33][203] = 9'b111111111;
assign micromatrizz[33][204] = 9'b111111111;
assign micromatrizz[33][205] = 9'b111111111;
assign micromatrizz[33][206] = 9'b111111111;
assign micromatrizz[33][207] = 9'b111111111;
assign micromatrizz[33][208] = 9'b111111111;
assign micromatrizz[33][209] = 9'b111111111;
assign micromatrizz[33][210] = 9'b111111111;
assign micromatrizz[33][211] = 9'b111111111;
assign micromatrizz[33][212] = 9'b111111111;
assign micromatrizz[33][213] = 9'b111111111;
assign micromatrizz[33][214] = 9'b111111111;
assign micromatrizz[33][215] = 9'b111111111;
assign micromatrizz[33][216] = 9'b111111111;
assign micromatrizz[33][217] = 9'b111111111;
assign micromatrizz[33][218] = 9'b111111111;
assign micromatrizz[33][219] = 9'b111111111;
assign micromatrizz[33][220] = 9'b111111111;
assign micromatrizz[33][221] = 9'b111111111;
assign micromatrizz[33][222] = 9'b111111111;
assign micromatrizz[33][223] = 9'b111111111;
assign micromatrizz[33][224] = 9'b111111111;
assign micromatrizz[33][225] = 9'b111111111;
assign micromatrizz[33][226] = 9'b111111111;
assign micromatrizz[33][227] = 9'b111111111;
assign micromatrizz[33][228] = 9'b111111111;
assign micromatrizz[33][229] = 9'b111111111;
assign micromatrizz[33][230] = 9'b111111111;
assign micromatrizz[33][231] = 9'b111111111;
assign micromatrizz[33][232] = 9'b111111111;
assign micromatrizz[33][233] = 9'b111111111;
assign micromatrizz[33][234] = 9'b111111111;
assign micromatrizz[33][235] = 9'b111111111;
assign micromatrizz[33][236] = 9'b111111111;
assign micromatrizz[33][237] = 9'b111111111;
assign micromatrizz[33][238] = 9'b111111111;
assign micromatrizz[33][239] = 9'b111111111;
assign micromatrizz[33][240] = 9'b111111111;
assign micromatrizz[33][241] = 9'b111111111;
assign micromatrizz[33][242] = 9'b111111111;
assign micromatrizz[33][243] = 9'b111111111;
assign micromatrizz[33][244] = 9'b111111111;
assign micromatrizz[33][245] = 9'b111111111;
assign micromatrizz[33][246] = 9'b111111111;
assign micromatrizz[33][247] = 9'b111111111;
assign micromatrizz[33][248] = 9'b111111111;
assign micromatrizz[33][249] = 9'b111111111;
assign micromatrizz[33][250] = 9'b111111111;
assign micromatrizz[33][251] = 9'b111111111;
assign micromatrizz[33][252] = 9'b111111111;
assign micromatrizz[33][253] = 9'b111111111;
assign micromatrizz[33][254] = 9'b111111111;
assign micromatrizz[33][255] = 9'b111111111;
assign micromatrizz[33][256] = 9'b111111111;
assign micromatrizz[33][257] = 9'b111111111;
assign micromatrizz[33][258] = 9'b111111111;
assign micromatrizz[33][259] = 9'b111111111;
assign micromatrizz[33][260] = 9'b111111111;
assign micromatrizz[33][261] = 9'b111111111;
assign micromatrizz[33][262] = 9'b111111111;
assign micromatrizz[33][263] = 9'b111111111;
assign micromatrizz[33][264] = 9'b111111111;
assign micromatrizz[33][265] = 9'b111111111;
assign micromatrizz[33][266] = 9'b111111111;
assign micromatrizz[33][267] = 9'b111111111;
assign micromatrizz[33][268] = 9'b111111111;
assign micromatrizz[33][269] = 9'b111111111;
assign micromatrizz[33][270] = 9'b111110110;
assign micromatrizz[33][271] = 9'b111110010;
assign micromatrizz[33][272] = 9'b111110010;
assign micromatrizz[33][273] = 9'b111110010;
assign micromatrizz[33][274] = 9'b111110011;
assign micromatrizz[33][275] = 9'b111110011;
assign micromatrizz[33][276] = 9'b111110011;
assign micromatrizz[33][277] = 9'b111110011;
assign micromatrizz[33][278] = 9'b111110011;
assign micromatrizz[33][279] = 9'b111111111;
assign micromatrizz[33][280] = 9'b111111111;
assign micromatrizz[33][281] = 9'b111111111;
assign micromatrizz[33][282] = 9'b111111111;
assign micromatrizz[33][283] = 9'b111111111;
assign micromatrizz[33][284] = 9'b111111111;
assign micromatrizz[33][285] = 9'b111111111;
assign micromatrizz[33][286] = 9'b111111111;
assign micromatrizz[33][287] = 9'b111111111;
assign micromatrizz[33][288] = 9'b111111111;
assign micromatrizz[33][289] = 9'b111111111;
assign micromatrizz[33][290] = 9'b111110111;
assign micromatrizz[33][291] = 9'b111110010;
assign micromatrizz[33][292] = 9'b111110011;
assign micromatrizz[33][293] = 9'b111110011;
assign micromatrizz[33][294] = 9'b111110011;
assign micromatrizz[33][295] = 9'b111110011;
assign micromatrizz[33][296] = 9'b111110011;
assign micromatrizz[33][297] = 9'b111110111;
assign micromatrizz[33][298] = 9'b111111111;
assign micromatrizz[33][299] = 9'b111111111;
assign micromatrizz[33][300] = 9'b111111111;
assign micromatrizz[33][301] = 9'b111111111;
assign micromatrizz[33][302] = 9'b111111111;
assign micromatrizz[33][303] = 9'b111111111;
assign micromatrizz[33][304] = 9'b111111111;
assign micromatrizz[33][305] = 9'b111110111;
assign micromatrizz[33][306] = 9'b111111111;
assign micromatrizz[33][307] = 9'b111111111;
assign micromatrizz[33][308] = 9'b111111111;
assign micromatrizz[33][309] = 9'b111111111;
assign micromatrizz[33][310] = 9'b111111111;
assign micromatrizz[33][311] = 9'b111111111;
assign micromatrizz[33][312] = 9'b111111111;
assign micromatrizz[33][313] = 9'b111110010;
assign micromatrizz[33][314] = 9'b111110010;
assign micromatrizz[33][315] = 9'b111110010;
assign micromatrizz[33][316] = 9'b111110010;
assign micromatrizz[33][317] = 9'b111110011;
assign micromatrizz[33][318] = 9'b111110011;
assign micromatrizz[33][319] = 9'b111110011;
assign micromatrizz[33][320] = 9'b111110011;
assign micromatrizz[33][321] = 9'b111111111;
assign micromatrizz[33][322] = 9'b111111111;
assign micromatrizz[33][323] = 9'b111111111;
assign micromatrizz[33][324] = 9'b111111111;
assign micromatrizz[33][325] = 9'b111111111;
assign micromatrizz[33][326] = 9'b111111111;
assign micromatrizz[33][327] = 9'b111111111;
assign micromatrizz[33][328] = 9'b111111111;
assign micromatrizz[33][329] = 9'b111111111;
assign micromatrizz[33][330] = 9'b111111111;
assign micromatrizz[33][331] = 9'b111111111;
assign micromatrizz[33][332] = 9'b111111111;
assign micromatrizz[33][333] = 9'b111111111;
assign micromatrizz[33][334] = 9'b111111111;
assign micromatrizz[33][335] = 9'b111111111;
assign micromatrizz[33][336] = 9'b111111111;
assign micromatrizz[33][337] = 9'b111111111;
assign micromatrizz[33][338] = 9'b111111111;
assign micromatrizz[33][339] = 9'b111111111;
assign micromatrizz[33][340] = 9'b111111111;
assign micromatrizz[33][341] = 9'b111111111;
assign micromatrizz[33][342] = 9'b111111111;
assign micromatrizz[33][343] = 9'b111111111;
assign micromatrizz[33][344] = 9'b111111111;
assign micromatrizz[33][345] = 9'b111111111;
assign micromatrizz[33][346] = 9'b111111111;
assign micromatrizz[33][347] = 9'b111111111;
assign micromatrizz[33][348] = 9'b111111111;
assign micromatrizz[33][349] = 9'b111111111;
assign micromatrizz[33][350] = 9'b111111111;
assign micromatrizz[33][351] = 9'b111111111;
assign micromatrizz[33][352] = 9'b111111111;
assign micromatrizz[33][353] = 9'b111111111;
assign micromatrizz[33][354] = 9'b111111111;
assign micromatrizz[33][355] = 9'b111111111;
assign micromatrizz[33][356] = 9'b111111111;
assign micromatrizz[33][357] = 9'b111111111;
assign micromatrizz[33][358] = 9'b111111111;
assign micromatrizz[33][359] = 9'b111111111;
assign micromatrizz[33][360] = 9'b111111111;
assign micromatrizz[33][361] = 9'b111111111;
assign micromatrizz[33][362] = 9'b111111111;
assign micromatrizz[33][363] = 9'b111111111;
assign micromatrizz[33][364] = 9'b111111111;
assign micromatrizz[33][365] = 9'b111111111;
assign micromatrizz[33][366] = 9'b111111111;
assign micromatrizz[33][367] = 9'b111111111;
assign micromatrizz[33][368] = 9'b111111111;
assign micromatrizz[33][369] = 9'b111111111;
assign micromatrizz[33][370] = 9'b111111111;
assign micromatrizz[33][371] = 9'b111111111;
assign micromatrizz[33][372] = 9'b111111111;
assign micromatrizz[33][373] = 9'b111111111;
assign micromatrizz[33][374] = 9'b111111111;
assign micromatrizz[33][375] = 9'b111111111;
assign micromatrizz[33][376] = 9'b111111111;
assign micromatrizz[33][377] = 9'b111111111;
assign micromatrizz[33][378] = 9'b111111111;
assign micromatrizz[33][379] = 9'b111111111;
assign micromatrizz[33][380] = 9'b111111111;
assign micromatrizz[33][381] = 9'b111111111;
assign micromatrizz[33][382] = 9'b111111111;
assign micromatrizz[33][383] = 9'b111111111;
assign micromatrizz[33][384] = 9'b111111111;
assign micromatrizz[33][385] = 9'b111111111;
assign micromatrizz[33][386] = 9'b111111111;
assign micromatrizz[33][387] = 9'b111111111;
assign micromatrizz[33][388] = 9'b111111111;
assign micromatrizz[33][389] = 9'b111111111;
assign micromatrizz[33][390] = 9'b111111111;
assign micromatrizz[33][391] = 9'b111111111;
assign micromatrizz[33][392] = 9'b111111111;
assign micromatrizz[33][393] = 9'b111111111;
assign micromatrizz[33][394] = 9'b111111111;
assign micromatrizz[33][395] = 9'b111111111;
assign micromatrizz[33][396] = 9'b111111111;
assign micromatrizz[33][397] = 9'b111111111;
assign micromatrizz[33][398] = 9'b111111111;
assign micromatrizz[33][399] = 9'b111111111;
assign micromatrizz[33][400] = 9'b111111111;
assign micromatrizz[33][401] = 9'b111111111;
assign micromatrizz[33][402] = 9'b111111111;
assign micromatrizz[33][403] = 9'b111111111;
assign micromatrizz[33][404] = 9'b111111111;
assign micromatrizz[33][405] = 9'b111111111;
assign micromatrizz[33][406] = 9'b111111111;
assign micromatrizz[33][407] = 9'b111111111;
assign micromatrizz[33][408] = 9'b111111111;
assign micromatrizz[33][409] = 9'b111111111;
assign micromatrizz[33][410] = 9'b111111111;
assign micromatrizz[33][411] = 9'b111111111;
assign micromatrizz[33][412] = 9'b111111111;
assign micromatrizz[33][413] = 9'b111111111;
assign micromatrizz[33][414] = 9'b111111111;
assign micromatrizz[33][415] = 9'b111111111;
assign micromatrizz[33][416] = 9'b111111111;
assign micromatrizz[33][417] = 9'b111111111;
assign micromatrizz[33][418] = 9'b111111111;
assign micromatrizz[33][419] = 9'b111111111;
assign micromatrizz[33][420] = 9'b111111111;
assign micromatrizz[33][421] = 9'b111111111;
assign micromatrizz[33][422] = 9'b111111111;
assign micromatrizz[33][423] = 9'b111111111;
assign micromatrizz[33][424] = 9'b111111111;
assign micromatrizz[33][425] = 9'b111111111;
assign micromatrizz[33][426] = 9'b111111111;
assign micromatrizz[33][427] = 9'b111111111;
assign micromatrizz[33][428] = 9'b111111111;
assign micromatrizz[33][429] = 9'b111111111;
assign micromatrizz[33][430] = 9'b111111111;
assign micromatrizz[33][431] = 9'b111111111;
assign micromatrizz[33][432] = 9'b111111111;
assign micromatrizz[33][433] = 9'b111111111;
assign micromatrizz[33][434] = 9'b111111111;
assign micromatrizz[33][435] = 9'b111111111;
assign micromatrizz[33][436] = 9'b111111111;
assign micromatrizz[33][437] = 9'b111111111;
assign micromatrizz[33][438] = 9'b111111111;
assign micromatrizz[33][439] = 9'b111111111;
assign micromatrizz[33][440] = 9'b111111111;
assign micromatrizz[33][441] = 9'b111111111;
assign micromatrizz[33][442] = 9'b111111111;
assign micromatrizz[33][443] = 9'b111111111;
assign micromatrizz[33][444] = 9'b111111111;
assign micromatrizz[33][445] = 9'b111111111;
assign micromatrizz[33][446] = 9'b111111111;
assign micromatrizz[33][447] = 9'b111111111;
assign micromatrizz[33][448] = 9'b111111111;
assign micromatrizz[33][449] = 9'b111111111;
assign micromatrizz[33][450] = 9'b111111111;
assign micromatrizz[33][451] = 9'b111111111;
assign micromatrizz[33][452] = 9'b111111111;
assign micromatrizz[33][453] = 9'b111111111;
assign micromatrizz[33][454] = 9'b111111111;
assign micromatrizz[33][455] = 9'b111111111;
assign micromatrizz[33][456] = 9'b111111111;
assign micromatrizz[33][457] = 9'b111111111;
assign micromatrizz[33][458] = 9'b111111111;
assign micromatrizz[33][459] = 9'b111111111;
assign micromatrizz[33][460] = 9'b111111111;
assign micromatrizz[33][461] = 9'b111111111;
assign micromatrizz[33][462] = 9'b111111111;
assign micromatrizz[33][463] = 9'b111111111;
assign micromatrizz[33][464] = 9'b111111111;
assign micromatrizz[33][465] = 9'b111111111;
assign micromatrizz[33][466] = 9'b111111111;
assign micromatrizz[33][467] = 9'b111111111;
assign micromatrizz[33][468] = 9'b111111111;
assign micromatrizz[33][469] = 9'b111111111;
assign micromatrizz[33][470] = 9'b111111111;
assign micromatrizz[33][471] = 9'b111111111;
assign micromatrizz[33][472] = 9'b111111111;
assign micromatrizz[33][473] = 9'b111111111;
assign micromatrizz[33][474] = 9'b111111111;
assign micromatrizz[33][475] = 9'b111111111;
assign micromatrizz[33][476] = 9'b111111111;
assign micromatrizz[33][477] = 9'b111111111;
assign micromatrizz[33][478] = 9'b111111111;
assign micromatrizz[33][479] = 9'b111111111;
assign micromatrizz[33][480] = 9'b111111111;
assign micromatrizz[33][481] = 9'b111111111;
assign micromatrizz[33][482] = 9'b111111111;
assign micromatrizz[33][483] = 9'b111111111;
assign micromatrizz[33][484] = 9'b111111111;
assign micromatrizz[33][485] = 9'b111111111;
assign micromatrizz[33][486] = 9'b111111111;
assign micromatrizz[33][487] = 9'b111111111;
assign micromatrizz[33][488] = 9'b111111111;
assign micromatrizz[33][489] = 9'b111111111;
assign micromatrizz[33][490] = 9'b111111111;
assign micromatrizz[33][491] = 9'b111111111;
assign micromatrizz[33][492] = 9'b111111111;
assign micromatrizz[33][493] = 9'b111111111;
assign micromatrizz[33][494] = 9'b111111111;
assign micromatrizz[33][495] = 9'b111111111;
assign micromatrizz[33][496] = 9'b111111111;
assign micromatrizz[33][497] = 9'b111111111;
assign micromatrizz[33][498] = 9'b111111111;
assign micromatrizz[33][499] = 9'b111111111;
assign micromatrizz[33][500] = 9'b111111111;
assign micromatrizz[33][501] = 9'b111111111;
assign micromatrizz[33][502] = 9'b111111111;
assign micromatrizz[33][503] = 9'b111111111;
assign micromatrizz[33][504] = 9'b111111111;
assign micromatrizz[33][505] = 9'b111111111;
assign micromatrizz[33][506] = 9'b111111111;
assign micromatrizz[33][507] = 9'b111111111;
assign micromatrizz[33][508] = 9'b111111111;
assign micromatrizz[33][509] = 9'b111111111;
assign micromatrizz[33][510] = 9'b111111111;
assign micromatrizz[33][511] = 9'b111111111;
assign micromatrizz[33][512] = 9'b111111111;
assign micromatrizz[33][513] = 9'b111111111;
assign micromatrizz[33][514] = 9'b111111111;
assign micromatrizz[33][515] = 9'b111111111;
assign micromatrizz[33][516] = 9'b111111111;
assign micromatrizz[33][517] = 9'b111111111;
assign micromatrizz[33][518] = 9'b111111111;
assign micromatrizz[33][519] = 9'b111111111;
assign micromatrizz[33][520] = 9'b111111111;
assign micromatrizz[33][521] = 9'b111111111;
assign micromatrizz[33][522] = 9'b111111111;
assign micromatrizz[33][523] = 9'b111111111;
assign micromatrizz[33][524] = 9'b111111111;
assign micromatrizz[33][525] = 9'b111111111;
assign micromatrizz[33][526] = 9'b111111111;
assign micromatrizz[33][527] = 9'b111111111;
assign micromatrizz[33][528] = 9'b111111111;
assign micromatrizz[33][529] = 9'b111111111;
assign micromatrizz[33][530] = 9'b111111111;
assign micromatrizz[33][531] = 9'b111111111;
assign micromatrizz[33][532] = 9'b111111111;
assign micromatrizz[33][533] = 9'b111111111;
assign micromatrizz[33][534] = 9'b111111111;
assign micromatrizz[33][535] = 9'b111111111;
assign micromatrizz[33][536] = 9'b111111111;
assign micromatrizz[33][537] = 9'b111111111;
assign micromatrizz[33][538] = 9'b111111111;
assign micromatrizz[33][539] = 9'b111111111;
assign micromatrizz[33][540] = 9'b111111111;
assign micromatrizz[33][541] = 9'b111111111;
assign micromatrizz[33][542] = 9'b111111111;
assign micromatrizz[33][543] = 9'b111111111;
assign micromatrizz[33][544] = 9'b111111111;
assign micromatrizz[33][545] = 9'b111111111;
assign micromatrizz[33][546] = 9'b111111111;
assign micromatrizz[33][547] = 9'b111111111;
assign micromatrizz[33][548] = 9'b111111111;
assign micromatrizz[33][549] = 9'b111111111;
assign micromatrizz[33][550] = 9'b111111111;
assign micromatrizz[33][551] = 9'b111111111;
assign micromatrizz[33][552] = 9'b111111111;
assign micromatrizz[33][553] = 9'b111111111;
assign micromatrizz[33][554] = 9'b111111111;
assign micromatrizz[33][555] = 9'b111111111;
assign micromatrizz[33][556] = 9'b111111111;
assign micromatrizz[33][557] = 9'b111111111;
assign micromatrizz[33][558] = 9'b111111111;
assign micromatrizz[33][559] = 9'b111111111;
assign micromatrizz[33][560] = 9'b111111111;
assign micromatrizz[33][561] = 9'b111111111;
assign micromatrizz[33][562] = 9'b111111111;
assign micromatrizz[33][563] = 9'b111111111;
assign micromatrizz[33][564] = 9'b111111111;
assign micromatrizz[33][565] = 9'b111111111;
assign micromatrizz[33][566] = 9'b111111111;
assign micromatrizz[33][567] = 9'b111111111;
assign micromatrizz[33][568] = 9'b111111111;
assign micromatrizz[33][569] = 9'b111111111;
assign micromatrizz[33][570] = 9'b111111111;
assign micromatrizz[33][571] = 9'b111111111;
assign micromatrizz[33][572] = 9'b111111111;
assign micromatrizz[33][573] = 9'b111111111;
assign micromatrizz[33][574] = 9'b111111111;
assign micromatrizz[33][575] = 9'b111111111;
assign micromatrizz[33][576] = 9'b111111111;
assign micromatrizz[33][577] = 9'b111111111;
assign micromatrizz[33][578] = 9'b111111111;
assign micromatrizz[33][579] = 9'b111111111;
assign micromatrizz[33][580] = 9'b111111111;
assign micromatrizz[33][581] = 9'b111111111;
assign micromatrizz[33][582] = 9'b111111111;
assign micromatrizz[33][583] = 9'b111111111;
assign micromatrizz[33][584] = 9'b111111111;
assign micromatrizz[33][585] = 9'b111111111;
assign micromatrizz[33][586] = 9'b111111111;
assign micromatrizz[33][587] = 9'b111111111;
assign micromatrizz[33][588] = 9'b111111111;
assign micromatrizz[33][589] = 9'b111111111;
assign micromatrizz[33][590] = 9'b111111111;
assign micromatrizz[33][591] = 9'b111111111;
assign micromatrizz[33][592] = 9'b111111111;
assign micromatrizz[33][593] = 9'b111111111;
assign micromatrizz[33][594] = 9'b111111111;
assign micromatrizz[33][595] = 9'b111111111;
assign micromatrizz[33][596] = 9'b111111111;
assign micromatrizz[33][597] = 9'b111111111;
assign micromatrizz[33][598] = 9'b111111111;
assign micromatrizz[33][599] = 9'b111111111;
assign micromatrizz[33][600] = 9'b111111111;
assign micromatrizz[33][601] = 9'b111111111;
assign micromatrizz[33][602] = 9'b111111111;
assign micromatrizz[33][603] = 9'b111111111;
assign micromatrizz[33][604] = 9'b111111111;
assign micromatrizz[33][605] = 9'b111111111;
assign micromatrizz[33][606] = 9'b111111111;
assign micromatrizz[33][607] = 9'b111111111;
assign micromatrizz[33][608] = 9'b111111111;
assign micromatrizz[33][609] = 9'b111111111;
assign micromatrizz[33][610] = 9'b111111111;
assign micromatrizz[33][611] = 9'b111111111;
assign micromatrizz[33][612] = 9'b111111111;
assign micromatrizz[33][613] = 9'b111111111;
assign micromatrizz[33][614] = 9'b111111111;
assign micromatrizz[33][615] = 9'b111111111;
assign micromatrizz[33][616] = 9'b111111111;
assign micromatrizz[33][617] = 9'b111111111;
assign micromatrizz[33][618] = 9'b111111111;
assign micromatrizz[33][619] = 9'b111111111;
assign micromatrizz[33][620] = 9'b111111111;
assign micromatrizz[33][621] = 9'b111111111;
assign micromatrizz[33][622] = 9'b111111111;
assign micromatrizz[33][623] = 9'b111111111;
assign micromatrizz[33][624] = 9'b111111111;
assign micromatrizz[33][625] = 9'b111111111;
assign micromatrizz[33][626] = 9'b111111111;
assign micromatrizz[33][627] = 9'b111111111;
assign micromatrizz[33][628] = 9'b111111111;
assign micromatrizz[33][629] = 9'b111111111;
assign micromatrizz[33][630] = 9'b111111111;
assign micromatrizz[33][631] = 9'b111111111;
assign micromatrizz[33][632] = 9'b111111111;
assign micromatrizz[33][633] = 9'b111111111;
assign micromatrizz[33][634] = 9'b111111111;
assign micromatrizz[33][635] = 9'b111111111;
assign micromatrizz[33][636] = 9'b111111111;
assign micromatrizz[33][637] = 9'b111111111;
assign micromatrizz[33][638] = 9'b111111111;
assign micromatrizz[33][639] = 9'b111111111;
assign micromatrizz[34][0] = 9'b111111111;
assign micromatrizz[34][1] = 9'b111111111;
assign micromatrizz[34][2] = 9'b111111111;
assign micromatrizz[34][3] = 9'b111111111;
assign micromatrizz[34][4] = 9'b111111111;
assign micromatrizz[34][5] = 9'b111111111;
assign micromatrizz[34][6] = 9'b111111111;
assign micromatrizz[34][7] = 9'b111111111;
assign micromatrizz[34][8] = 9'b111111111;
assign micromatrizz[34][9] = 9'b111111111;
assign micromatrizz[34][10] = 9'b111111111;
assign micromatrizz[34][11] = 9'b111111111;
assign micromatrizz[34][12] = 9'b111111111;
assign micromatrizz[34][13] = 9'b111111111;
assign micromatrizz[34][14] = 9'b111111111;
assign micromatrizz[34][15] = 9'b111111111;
assign micromatrizz[34][16] = 9'b111111111;
assign micromatrizz[34][17] = 9'b111111111;
assign micromatrizz[34][18] = 9'b111111111;
assign micromatrizz[34][19] = 9'b111111111;
assign micromatrizz[34][20] = 9'b111111111;
assign micromatrizz[34][21] = 9'b111111111;
assign micromatrizz[34][22] = 9'b111111111;
assign micromatrizz[34][23] = 9'b111111111;
assign micromatrizz[34][24] = 9'b111111111;
assign micromatrizz[34][25] = 9'b111111111;
assign micromatrizz[34][26] = 9'b111111111;
assign micromatrizz[34][27] = 9'b111111111;
assign micromatrizz[34][28] = 9'b111111111;
assign micromatrizz[34][29] = 9'b111111111;
assign micromatrizz[34][30] = 9'b111111111;
assign micromatrizz[34][31] = 9'b111111111;
assign micromatrizz[34][32] = 9'b111111111;
assign micromatrizz[34][33] = 9'b111111111;
assign micromatrizz[34][34] = 9'b111111111;
assign micromatrizz[34][35] = 9'b111111111;
assign micromatrizz[34][36] = 9'b111111111;
assign micromatrizz[34][37] = 9'b111111111;
assign micromatrizz[34][38] = 9'b111111111;
assign micromatrizz[34][39] = 9'b111111111;
assign micromatrizz[34][40] = 9'b111111111;
assign micromatrizz[34][41] = 9'b111111111;
assign micromatrizz[34][42] = 9'b111111111;
assign micromatrizz[34][43] = 9'b111111111;
assign micromatrizz[34][44] = 9'b111111111;
assign micromatrizz[34][45] = 9'b111111111;
assign micromatrizz[34][46] = 9'b111111111;
assign micromatrizz[34][47] = 9'b111111111;
assign micromatrizz[34][48] = 9'b111111111;
assign micromatrizz[34][49] = 9'b111111111;
assign micromatrizz[34][50] = 9'b111111111;
assign micromatrizz[34][51] = 9'b111111111;
assign micromatrizz[34][52] = 9'b111111111;
assign micromatrizz[34][53] = 9'b111111111;
assign micromatrizz[34][54] = 9'b111111111;
assign micromatrizz[34][55] = 9'b111111111;
assign micromatrizz[34][56] = 9'b111111111;
assign micromatrizz[34][57] = 9'b111111111;
assign micromatrizz[34][58] = 9'b111111111;
assign micromatrizz[34][59] = 9'b111111111;
assign micromatrizz[34][60] = 9'b111111111;
assign micromatrizz[34][61] = 9'b111111111;
assign micromatrizz[34][62] = 9'b111111111;
assign micromatrizz[34][63] = 9'b111111111;
assign micromatrizz[34][64] = 9'b111111111;
assign micromatrizz[34][65] = 9'b111111111;
assign micromatrizz[34][66] = 9'b111111111;
assign micromatrizz[34][67] = 9'b111111111;
assign micromatrizz[34][68] = 9'b111111111;
assign micromatrizz[34][69] = 9'b111111111;
assign micromatrizz[34][70] = 9'b111111111;
assign micromatrizz[34][71] = 9'b111111111;
assign micromatrizz[34][72] = 9'b111111111;
assign micromatrizz[34][73] = 9'b111111111;
assign micromatrizz[34][74] = 9'b111111111;
assign micromatrizz[34][75] = 9'b111111111;
assign micromatrizz[34][76] = 9'b111111111;
assign micromatrizz[34][77] = 9'b111111111;
assign micromatrizz[34][78] = 9'b111111111;
assign micromatrizz[34][79] = 9'b111111111;
assign micromatrizz[34][80] = 9'b111111111;
assign micromatrizz[34][81] = 9'b111111111;
assign micromatrizz[34][82] = 9'b111111111;
assign micromatrizz[34][83] = 9'b111111111;
assign micromatrizz[34][84] = 9'b111111111;
assign micromatrizz[34][85] = 9'b111111111;
assign micromatrizz[34][86] = 9'b111111111;
assign micromatrizz[34][87] = 9'b111111111;
assign micromatrizz[34][88] = 9'b111111111;
assign micromatrizz[34][89] = 9'b111111111;
assign micromatrizz[34][90] = 9'b111111111;
assign micromatrizz[34][91] = 9'b111111111;
assign micromatrizz[34][92] = 9'b111111111;
assign micromatrizz[34][93] = 9'b111111111;
assign micromatrizz[34][94] = 9'b111111111;
assign micromatrizz[34][95] = 9'b111111111;
assign micromatrizz[34][96] = 9'b111111111;
assign micromatrizz[34][97] = 9'b111111111;
assign micromatrizz[34][98] = 9'b111111111;
assign micromatrizz[34][99] = 9'b111111111;
assign micromatrizz[34][100] = 9'b111111111;
assign micromatrizz[34][101] = 9'b111111111;
assign micromatrizz[34][102] = 9'b111111111;
assign micromatrizz[34][103] = 9'b111111111;
assign micromatrizz[34][104] = 9'b111111111;
assign micromatrizz[34][105] = 9'b111111111;
assign micromatrizz[34][106] = 9'b111111111;
assign micromatrizz[34][107] = 9'b111111111;
assign micromatrizz[34][108] = 9'b111111111;
assign micromatrizz[34][109] = 9'b111111111;
assign micromatrizz[34][110] = 9'b111111111;
assign micromatrizz[34][111] = 9'b111111111;
assign micromatrizz[34][112] = 9'b111111111;
assign micromatrizz[34][113] = 9'b111111111;
assign micromatrizz[34][114] = 9'b111111111;
assign micromatrizz[34][115] = 9'b111111111;
assign micromatrizz[34][116] = 9'b111111111;
assign micromatrizz[34][117] = 9'b111111111;
assign micromatrizz[34][118] = 9'b111111111;
assign micromatrizz[34][119] = 9'b111111111;
assign micromatrizz[34][120] = 9'b111111111;
assign micromatrizz[34][121] = 9'b111111111;
assign micromatrizz[34][122] = 9'b111111111;
assign micromatrizz[34][123] = 9'b111111111;
assign micromatrizz[34][124] = 9'b111111111;
assign micromatrizz[34][125] = 9'b111111111;
assign micromatrizz[34][126] = 9'b111111111;
assign micromatrizz[34][127] = 9'b111111111;
assign micromatrizz[34][128] = 9'b111111111;
assign micromatrizz[34][129] = 9'b111111111;
assign micromatrizz[34][130] = 9'b111111111;
assign micromatrizz[34][131] = 9'b111111111;
assign micromatrizz[34][132] = 9'b111111111;
assign micromatrizz[34][133] = 9'b111111111;
assign micromatrizz[34][134] = 9'b111111111;
assign micromatrizz[34][135] = 9'b111111111;
assign micromatrizz[34][136] = 9'b111111111;
assign micromatrizz[34][137] = 9'b111111111;
assign micromatrizz[34][138] = 9'b111111111;
assign micromatrizz[34][139] = 9'b111111111;
assign micromatrizz[34][140] = 9'b111111111;
assign micromatrizz[34][141] = 9'b111111111;
assign micromatrizz[34][142] = 9'b111111111;
assign micromatrizz[34][143] = 9'b111111111;
assign micromatrizz[34][144] = 9'b111111111;
assign micromatrizz[34][145] = 9'b111111111;
assign micromatrizz[34][146] = 9'b111111111;
assign micromatrizz[34][147] = 9'b111111111;
assign micromatrizz[34][148] = 9'b111111111;
assign micromatrizz[34][149] = 9'b111111111;
assign micromatrizz[34][150] = 9'b111111111;
assign micromatrizz[34][151] = 9'b111111111;
assign micromatrizz[34][152] = 9'b111111111;
assign micromatrizz[34][153] = 9'b111111111;
assign micromatrizz[34][154] = 9'b111111111;
assign micromatrizz[34][155] = 9'b111111111;
assign micromatrizz[34][156] = 9'b111111111;
assign micromatrizz[34][157] = 9'b111111111;
assign micromatrizz[34][158] = 9'b111111111;
assign micromatrizz[34][159] = 9'b111111111;
assign micromatrizz[34][160] = 9'b111111111;
assign micromatrizz[34][161] = 9'b111111111;
assign micromatrizz[34][162] = 9'b111111111;
assign micromatrizz[34][163] = 9'b111111111;
assign micromatrizz[34][164] = 9'b111111111;
assign micromatrizz[34][165] = 9'b111111111;
assign micromatrizz[34][166] = 9'b111111111;
assign micromatrizz[34][167] = 9'b111111111;
assign micromatrizz[34][168] = 9'b111111111;
assign micromatrizz[34][169] = 9'b111111111;
assign micromatrizz[34][170] = 9'b111111111;
assign micromatrizz[34][171] = 9'b111111111;
assign micromatrizz[34][172] = 9'b111111111;
assign micromatrizz[34][173] = 9'b111111111;
assign micromatrizz[34][174] = 9'b111111111;
assign micromatrizz[34][175] = 9'b111111111;
assign micromatrizz[34][176] = 9'b111111111;
assign micromatrizz[34][177] = 9'b111111111;
assign micromatrizz[34][178] = 9'b111111111;
assign micromatrizz[34][179] = 9'b111111111;
assign micromatrizz[34][180] = 9'b111111111;
assign micromatrizz[34][181] = 9'b111111111;
assign micromatrizz[34][182] = 9'b111111111;
assign micromatrizz[34][183] = 9'b111111111;
assign micromatrizz[34][184] = 9'b111111111;
assign micromatrizz[34][185] = 9'b111111111;
assign micromatrizz[34][186] = 9'b111111111;
assign micromatrizz[34][187] = 9'b111111111;
assign micromatrizz[34][188] = 9'b111111111;
assign micromatrizz[34][189] = 9'b111111111;
assign micromatrizz[34][190] = 9'b111111111;
assign micromatrizz[34][191] = 9'b111111111;
assign micromatrizz[34][192] = 9'b111111111;
assign micromatrizz[34][193] = 9'b111111111;
assign micromatrizz[34][194] = 9'b111111111;
assign micromatrizz[34][195] = 9'b111111111;
assign micromatrizz[34][196] = 9'b111111111;
assign micromatrizz[34][197] = 9'b111111111;
assign micromatrizz[34][198] = 9'b111111111;
assign micromatrizz[34][199] = 9'b111111111;
assign micromatrizz[34][200] = 9'b111111111;
assign micromatrizz[34][201] = 9'b111111111;
assign micromatrizz[34][202] = 9'b111111111;
assign micromatrizz[34][203] = 9'b111111111;
assign micromatrizz[34][204] = 9'b111111111;
assign micromatrizz[34][205] = 9'b111111111;
assign micromatrizz[34][206] = 9'b111111111;
assign micromatrizz[34][207] = 9'b111111111;
assign micromatrizz[34][208] = 9'b111111111;
assign micromatrizz[34][209] = 9'b111111111;
assign micromatrizz[34][210] = 9'b111111111;
assign micromatrizz[34][211] = 9'b111111111;
assign micromatrizz[34][212] = 9'b111111111;
assign micromatrizz[34][213] = 9'b111111111;
assign micromatrizz[34][214] = 9'b111111111;
assign micromatrizz[34][215] = 9'b111111111;
assign micromatrizz[34][216] = 9'b111111111;
assign micromatrizz[34][217] = 9'b111111111;
assign micromatrizz[34][218] = 9'b111111111;
assign micromatrizz[34][219] = 9'b111111111;
assign micromatrizz[34][220] = 9'b111111111;
assign micromatrizz[34][221] = 9'b111111111;
assign micromatrizz[34][222] = 9'b111111111;
assign micromatrizz[34][223] = 9'b111111111;
assign micromatrizz[34][224] = 9'b111111111;
assign micromatrizz[34][225] = 9'b111111111;
assign micromatrizz[34][226] = 9'b111111111;
assign micromatrizz[34][227] = 9'b111111111;
assign micromatrizz[34][228] = 9'b111111111;
assign micromatrizz[34][229] = 9'b111111111;
assign micromatrizz[34][230] = 9'b111111111;
assign micromatrizz[34][231] = 9'b111111111;
assign micromatrizz[34][232] = 9'b111111111;
assign micromatrizz[34][233] = 9'b111111111;
assign micromatrizz[34][234] = 9'b111111111;
assign micromatrizz[34][235] = 9'b111111111;
assign micromatrizz[34][236] = 9'b111111111;
assign micromatrizz[34][237] = 9'b111111111;
assign micromatrizz[34][238] = 9'b111111111;
assign micromatrizz[34][239] = 9'b111111111;
assign micromatrizz[34][240] = 9'b111111111;
assign micromatrizz[34][241] = 9'b111111111;
assign micromatrizz[34][242] = 9'b111111111;
assign micromatrizz[34][243] = 9'b111111111;
assign micromatrizz[34][244] = 9'b111111111;
assign micromatrizz[34][245] = 9'b111111111;
assign micromatrizz[34][246] = 9'b111111111;
assign micromatrizz[34][247] = 9'b111111111;
assign micromatrizz[34][248] = 9'b111111111;
assign micromatrizz[34][249] = 9'b111111111;
assign micromatrizz[34][250] = 9'b111111111;
assign micromatrizz[34][251] = 9'b111111111;
assign micromatrizz[34][252] = 9'b111111111;
assign micromatrizz[34][253] = 9'b111111111;
assign micromatrizz[34][254] = 9'b111111111;
assign micromatrizz[34][255] = 9'b111111111;
assign micromatrizz[34][256] = 9'b111111111;
assign micromatrizz[34][257] = 9'b111111111;
assign micromatrizz[34][258] = 9'b111111111;
assign micromatrizz[34][259] = 9'b111111111;
assign micromatrizz[34][260] = 9'b111111111;
assign micromatrizz[34][261] = 9'b111111111;
assign micromatrizz[34][262] = 9'b111111111;
assign micromatrizz[34][263] = 9'b111111111;
assign micromatrizz[34][264] = 9'b111111111;
assign micromatrizz[34][265] = 9'b111111111;
assign micromatrizz[34][266] = 9'b111111111;
assign micromatrizz[34][267] = 9'b111111111;
assign micromatrizz[34][268] = 9'b111111111;
assign micromatrizz[34][269] = 9'b111111111;
assign micromatrizz[34][270] = 9'b111110010;
assign micromatrizz[34][271] = 9'b111110010;
assign micromatrizz[34][272] = 9'b111110010;
assign micromatrizz[34][273] = 9'b111110010;
assign micromatrizz[34][274] = 9'b111110011;
assign micromatrizz[34][275] = 9'b111110011;
assign micromatrizz[34][276] = 9'b111110011;
assign micromatrizz[34][277] = 9'b111110011;
assign micromatrizz[34][278] = 9'b111110011;
assign micromatrizz[34][279] = 9'b111111111;
assign micromatrizz[34][280] = 9'b111111111;
assign micromatrizz[34][281] = 9'b111111111;
assign micromatrizz[34][282] = 9'b111111111;
assign micromatrizz[34][283] = 9'b111111111;
assign micromatrizz[34][284] = 9'b111111111;
assign micromatrizz[34][285] = 9'b111111111;
assign micromatrizz[34][286] = 9'b111111111;
assign micromatrizz[34][287] = 9'b111111111;
assign micromatrizz[34][288] = 9'b111111111;
assign micromatrizz[34][289] = 9'b111111111;
assign micromatrizz[34][290] = 9'b111111111;
assign micromatrizz[34][291] = 9'b111110111;
assign micromatrizz[34][292] = 9'b111110010;
assign micromatrizz[34][293] = 9'b111110011;
assign micromatrizz[34][294] = 9'b111110011;
assign micromatrizz[34][295] = 9'b111110011;
assign micromatrizz[34][296] = 9'b111110011;
assign micromatrizz[34][297] = 9'b111110111;
assign micromatrizz[34][298] = 9'b111111111;
assign micromatrizz[34][299] = 9'b111111111;
assign micromatrizz[34][300] = 9'b111111111;
assign micromatrizz[34][301] = 9'b111111111;
assign micromatrizz[34][302] = 9'b111111111;
assign micromatrizz[34][303] = 9'b111111111;
assign micromatrizz[34][304] = 9'b111110111;
assign micromatrizz[34][305] = 9'b111111111;
assign micromatrizz[34][306] = 9'b111111111;
assign micromatrizz[34][307] = 9'b111111111;
assign micromatrizz[34][308] = 9'b111111111;
assign micromatrizz[34][309] = 9'b111111111;
assign micromatrizz[34][310] = 9'b111111111;
assign micromatrizz[34][311] = 9'b111111111;
assign micromatrizz[34][312] = 9'b111111111;
assign micromatrizz[34][313] = 9'b111111111;
assign micromatrizz[34][314] = 9'b111110011;
assign micromatrizz[34][315] = 9'b111110010;
assign micromatrizz[34][316] = 9'b111110011;
assign micromatrizz[34][317] = 9'b111110011;
assign micromatrizz[34][318] = 9'b111110011;
assign micromatrizz[34][319] = 9'b111110011;
assign micromatrizz[34][320] = 9'b111110010;
assign micromatrizz[34][321] = 9'b111111111;
assign micromatrizz[34][322] = 9'b111111111;
assign micromatrizz[34][323] = 9'b111111111;
assign micromatrizz[34][324] = 9'b111111111;
assign micromatrizz[34][325] = 9'b111111111;
assign micromatrizz[34][326] = 9'b111111111;
assign micromatrizz[34][327] = 9'b111111111;
assign micromatrizz[34][328] = 9'b111111111;
assign micromatrizz[34][329] = 9'b111111111;
assign micromatrizz[34][330] = 9'b111111111;
assign micromatrizz[34][331] = 9'b111111111;
assign micromatrizz[34][332] = 9'b111111111;
assign micromatrizz[34][333] = 9'b111111111;
assign micromatrizz[34][334] = 9'b111111111;
assign micromatrizz[34][335] = 9'b111111111;
assign micromatrizz[34][336] = 9'b111111111;
assign micromatrizz[34][337] = 9'b111111111;
assign micromatrizz[34][338] = 9'b111111111;
assign micromatrizz[34][339] = 9'b111111111;
assign micromatrizz[34][340] = 9'b111111111;
assign micromatrizz[34][341] = 9'b111111111;
assign micromatrizz[34][342] = 9'b111111111;
assign micromatrizz[34][343] = 9'b111111111;
assign micromatrizz[34][344] = 9'b111111111;
assign micromatrizz[34][345] = 9'b111111111;
assign micromatrizz[34][346] = 9'b111111111;
assign micromatrizz[34][347] = 9'b111111111;
assign micromatrizz[34][348] = 9'b111111111;
assign micromatrizz[34][349] = 9'b111111111;
assign micromatrizz[34][350] = 9'b111111111;
assign micromatrizz[34][351] = 9'b111111111;
assign micromatrizz[34][352] = 9'b111111111;
assign micromatrizz[34][353] = 9'b111111111;
assign micromatrizz[34][354] = 9'b111111111;
assign micromatrizz[34][355] = 9'b111111111;
assign micromatrizz[34][356] = 9'b111111111;
assign micromatrizz[34][357] = 9'b111111111;
assign micromatrizz[34][358] = 9'b111111111;
assign micromatrizz[34][359] = 9'b111111111;
assign micromatrizz[34][360] = 9'b111111111;
assign micromatrizz[34][361] = 9'b111111111;
assign micromatrizz[34][362] = 9'b111111111;
assign micromatrizz[34][363] = 9'b111111111;
assign micromatrizz[34][364] = 9'b111111111;
assign micromatrizz[34][365] = 9'b111111111;
assign micromatrizz[34][366] = 9'b111111111;
assign micromatrizz[34][367] = 9'b111111111;
assign micromatrizz[34][368] = 9'b111111111;
assign micromatrizz[34][369] = 9'b111111111;
assign micromatrizz[34][370] = 9'b111111111;
assign micromatrizz[34][371] = 9'b111111111;
assign micromatrizz[34][372] = 9'b111111111;
assign micromatrizz[34][373] = 9'b111111111;
assign micromatrizz[34][374] = 9'b111111111;
assign micromatrizz[34][375] = 9'b111111111;
assign micromatrizz[34][376] = 9'b111111111;
assign micromatrizz[34][377] = 9'b111111111;
assign micromatrizz[34][378] = 9'b111111111;
assign micromatrizz[34][379] = 9'b111111111;
assign micromatrizz[34][380] = 9'b111111111;
assign micromatrizz[34][381] = 9'b111111111;
assign micromatrizz[34][382] = 9'b111111111;
assign micromatrizz[34][383] = 9'b111111111;
assign micromatrizz[34][384] = 9'b111111111;
assign micromatrizz[34][385] = 9'b111111111;
assign micromatrizz[34][386] = 9'b111111111;
assign micromatrizz[34][387] = 9'b111111111;
assign micromatrizz[34][388] = 9'b111111111;
assign micromatrizz[34][389] = 9'b111111111;
assign micromatrizz[34][390] = 9'b111111111;
assign micromatrizz[34][391] = 9'b111111111;
assign micromatrizz[34][392] = 9'b111111111;
assign micromatrizz[34][393] = 9'b111111111;
assign micromatrizz[34][394] = 9'b111111111;
assign micromatrizz[34][395] = 9'b111111111;
assign micromatrizz[34][396] = 9'b111111111;
assign micromatrizz[34][397] = 9'b111111111;
assign micromatrizz[34][398] = 9'b111111111;
assign micromatrizz[34][399] = 9'b111111111;
assign micromatrizz[34][400] = 9'b111111111;
assign micromatrizz[34][401] = 9'b111111111;
assign micromatrizz[34][402] = 9'b111111111;
assign micromatrizz[34][403] = 9'b111111111;
assign micromatrizz[34][404] = 9'b111111111;
assign micromatrizz[34][405] = 9'b111111111;
assign micromatrizz[34][406] = 9'b111111111;
assign micromatrizz[34][407] = 9'b111111111;
assign micromatrizz[34][408] = 9'b111111111;
assign micromatrizz[34][409] = 9'b111111111;
assign micromatrizz[34][410] = 9'b111111111;
assign micromatrizz[34][411] = 9'b111111111;
assign micromatrizz[34][412] = 9'b111111111;
assign micromatrizz[34][413] = 9'b111111111;
assign micromatrizz[34][414] = 9'b111111111;
assign micromatrizz[34][415] = 9'b111111111;
assign micromatrizz[34][416] = 9'b111111111;
assign micromatrizz[34][417] = 9'b111111111;
assign micromatrizz[34][418] = 9'b111111111;
assign micromatrizz[34][419] = 9'b111111111;
assign micromatrizz[34][420] = 9'b111111111;
assign micromatrizz[34][421] = 9'b111111111;
assign micromatrizz[34][422] = 9'b111111111;
assign micromatrizz[34][423] = 9'b111111111;
assign micromatrizz[34][424] = 9'b111111111;
assign micromatrizz[34][425] = 9'b111111111;
assign micromatrizz[34][426] = 9'b111111111;
assign micromatrizz[34][427] = 9'b111111111;
assign micromatrizz[34][428] = 9'b111111111;
assign micromatrizz[34][429] = 9'b111111111;
assign micromatrizz[34][430] = 9'b111111111;
assign micromatrizz[34][431] = 9'b111111111;
assign micromatrizz[34][432] = 9'b111111111;
assign micromatrizz[34][433] = 9'b111111111;
assign micromatrizz[34][434] = 9'b111111111;
assign micromatrizz[34][435] = 9'b111111111;
assign micromatrizz[34][436] = 9'b111111111;
assign micromatrizz[34][437] = 9'b111111111;
assign micromatrizz[34][438] = 9'b111111111;
assign micromatrizz[34][439] = 9'b111111111;
assign micromatrizz[34][440] = 9'b111111111;
assign micromatrizz[34][441] = 9'b111111111;
assign micromatrizz[34][442] = 9'b111111111;
assign micromatrizz[34][443] = 9'b111111111;
assign micromatrizz[34][444] = 9'b111111111;
assign micromatrizz[34][445] = 9'b111111111;
assign micromatrizz[34][446] = 9'b111111111;
assign micromatrizz[34][447] = 9'b111111111;
assign micromatrizz[34][448] = 9'b111111111;
assign micromatrizz[34][449] = 9'b111111111;
assign micromatrizz[34][450] = 9'b111111111;
assign micromatrizz[34][451] = 9'b111111111;
assign micromatrizz[34][452] = 9'b111111111;
assign micromatrizz[34][453] = 9'b111111111;
assign micromatrizz[34][454] = 9'b111111111;
assign micromatrizz[34][455] = 9'b111111111;
assign micromatrizz[34][456] = 9'b111111111;
assign micromatrizz[34][457] = 9'b111111111;
assign micromatrizz[34][458] = 9'b111111111;
assign micromatrizz[34][459] = 9'b111111111;
assign micromatrizz[34][460] = 9'b111111111;
assign micromatrizz[34][461] = 9'b111111111;
assign micromatrizz[34][462] = 9'b111111111;
assign micromatrizz[34][463] = 9'b111111111;
assign micromatrizz[34][464] = 9'b111111111;
assign micromatrizz[34][465] = 9'b111111111;
assign micromatrizz[34][466] = 9'b111111111;
assign micromatrizz[34][467] = 9'b111111111;
assign micromatrizz[34][468] = 9'b111111111;
assign micromatrizz[34][469] = 9'b111111111;
assign micromatrizz[34][470] = 9'b111111111;
assign micromatrizz[34][471] = 9'b111111111;
assign micromatrizz[34][472] = 9'b111111111;
assign micromatrizz[34][473] = 9'b111111111;
assign micromatrizz[34][474] = 9'b111111111;
assign micromatrizz[34][475] = 9'b111111111;
assign micromatrizz[34][476] = 9'b111111111;
assign micromatrizz[34][477] = 9'b111111111;
assign micromatrizz[34][478] = 9'b111111111;
assign micromatrizz[34][479] = 9'b111111111;
assign micromatrizz[34][480] = 9'b111111111;
assign micromatrizz[34][481] = 9'b111111111;
assign micromatrizz[34][482] = 9'b111111111;
assign micromatrizz[34][483] = 9'b111111111;
assign micromatrizz[34][484] = 9'b111111111;
assign micromatrizz[34][485] = 9'b111111111;
assign micromatrizz[34][486] = 9'b111111111;
assign micromatrizz[34][487] = 9'b111111111;
assign micromatrizz[34][488] = 9'b111111111;
assign micromatrizz[34][489] = 9'b111111111;
assign micromatrizz[34][490] = 9'b111111111;
assign micromatrizz[34][491] = 9'b111111111;
assign micromatrizz[34][492] = 9'b111111111;
assign micromatrizz[34][493] = 9'b111111111;
assign micromatrizz[34][494] = 9'b111111111;
assign micromatrizz[34][495] = 9'b111111111;
assign micromatrizz[34][496] = 9'b111111111;
assign micromatrizz[34][497] = 9'b111111111;
assign micromatrizz[34][498] = 9'b111111111;
assign micromatrizz[34][499] = 9'b111111111;
assign micromatrizz[34][500] = 9'b111111111;
assign micromatrizz[34][501] = 9'b111111111;
assign micromatrizz[34][502] = 9'b111111111;
assign micromatrizz[34][503] = 9'b111111111;
assign micromatrizz[34][504] = 9'b111111111;
assign micromatrizz[34][505] = 9'b111111111;
assign micromatrizz[34][506] = 9'b111111111;
assign micromatrizz[34][507] = 9'b111111111;
assign micromatrizz[34][508] = 9'b111111111;
assign micromatrizz[34][509] = 9'b111111111;
assign micromatrizz[34][510] = 9'b111111111;
assign micromatrizz[34][511] = 9'b111111111;
assign micromatrizz[34][512] = 9'b111111111;
assign micromatrizz[34][513] = 9'b111111111;
assign micromatrizz[34][514] = 9'b111111111;
assign micromatrizz[34][515] = 9'b111111111;
assign micromatrizz[34][516] = 9'b111111111;
assign micromatrizz[34][517] = 9'b111111111;
assign micromatrizz[34][518] = 9'b111111111;
assign micromatrizz[34][519] = 9'b111111111;
assign micromatrizz[34][520] = 9'b111111111;
assign micromatrizz[34][521] = 9'b111111111;
assign micromatrizz[34][522] = 9'b111111111;
assign micromatrizz[34][523] = 9'b111111111;
assign micromatrizz[34][524] = 9'b111111111;
assign micromatrizz[34][525] = 9'b111111111;
assign micromatrizz[34][526] = 9'b111111111;
assign micromatrizz[34][527] = 9'b111111111;
assign micromatrizz[34][528] = 9'b111111111;
assign micromatrizz[34][529] = 9'b111111111;
assign micromatrizz[34][530] = 9'b111111111;
assign micromatrizz[34][531] = 9'b111111111;
assign micromatrizz[34][532] = 9'b111111111;
assign micromatrizz[34][533] = 9'b111111111;
assign micromatrizz[34][534] = 9'b111111111;
assign micromatrizz[34][535] = 9'b111111111;
assign micromatrizz[34][536] = 9'b111111111;
assign micromatrizz[34][537] = 9'b111111111;
assign micromatrizz[34][538] = 9'b111111111;
assign micromatrizz[34][539] = 9'b111111111;
assign micromatrizz[34][540] = 9'b111111111;
assign micromatrizz[34][541] = 9'b111111111;
assign micromatrizz[34][542] = 9'b111111111;
assign micromatrizz[34][543] = 9'b111111111;
assign micromatrizz[34][544] = 9'b111111111;
assign micromatrizz[34][545] = 9'b111111111;
assign micromatrizz[34][546] = 9'b111111111;
assign micromatrizz[34][547] = 9'b111111111;
assign micromatrizz[34][548] = 9'b111111111;
assign micromatrizz[34][549] = 9'b111111111;
assign micromatrizz[34][550] = 9'b111111111;
assign micromatrizz[34][551] = 9'b111111111;
assign micromatrizz[34][552] = 9'b111111111;
assign micromatrizz[34][553] = 9'b111111111;
assign micromatrizz[34][554] = 9'b111111111;
assign micromatrizz[34][555] = 9'b111111111;
assign micromatrizz[34][556] = 9'b111111111;
assign micromatrizz[34][557] = 9'b111111111;
assign micromatrizz[34][558] = 9'b111111111;
assign micromatrizz[34][559] = 9'b111111111;
assign micromatrizz[34][560] = 9'b111111111;
assign micromatrizz[34][561] = 9'b111111111;
assign micromatrizz[34][562] = 9'b111111111;
assign micromatrizz[34][563] = 9'b111111111;
assign micromatrizz[34][564] = 9'b111111111;
assign micromatrizz[34][565] = 9'b111111111;
assign micromatrizz[34][566] = 9'b111111111;
assign micromatrizz[34][567] = 9'b111111111;
assign micromatrizz[34][568] = 9'b111111111;
assign micromatrizz[34][569] = 9'b111111111;
assign micromatrizz[34][570] = 9'b111111111;
assign micromatrizz[34][571] = 9'b111111111;
assign micromatrizz[34][572] = 9'b111111111;
assign micromatrizz[34][573] = 9'b111111111;
assign micromatrizz[34][574] = 9'b111111111;
assign micromatrizz[34][575] = 9'b111111111;
assign micromatrizz[34][576] = 9'b111111111;
assign micromatrizz[34][577] = 9'b111111111;
assign micromatrizz[34][578] = 9'b111111111;
assign micromatrizz[34][579] = 9'b111111111;
assign micromatrizz[34][580] = 9'b111111111;
assign micromatrizz[34][581] = 9'b111111111;
assign micromatrizz[34][582] = 9'b111111111;
assign micromatrizz[34][583] = 9'b111111111;
assign micromatrizz[34][584] = 9'b111111111;
assign micromatrizz[34][585] = 9'b111111111;
assign micromatrizz[34][586] = 9'b111111111;
assign micromatrizz[34][587] = 9'b111111111;
assign micromatrizz[34][588] = 9'b111111111;
assign micromatrizz[34][589] = 9'b111111111;
assign micromatrizz[34][590] = 9'b111111111;
assign micromatrizz[34][591] = 9'b111111111;
assign micromatrizz[34][592] = 9'b111111111;
assign micromatrizz[34][593] = 9'b111111111;
assign micromatrizz[34][594] = 9'b111111111;
assign micromatrizz[34][595] = 9'b111111111;
assign micromatrizz[34][596] = 9'b111111111;
assign micromatrizz[34][597] = 9'b111111111;
assign micromatrizz[34][598] = 9'b111111111;
assign micromatrizz[34][599] = 9'b111111111;
assign micromatrizz[34][600] = 9'b111111111;
assign micromatrizz[34][601] = 9'b111111111;
assign micromatrizz[34][602] = 9'b111111111;
assign micromatrizz[34][603] = 9'b111111111;
assign micromatrizz[34][604] = 9'b111111111;
assign micromatrizz[34][605] = 9'b111111111;
assign micromatrizz[34][606] = 9'b111111111;
assign micromatrizz[34][607] = 9'b111111111;
assign micromatrizz[34][608] = 9'b111111111;
assign micromatrizz[34][609] = 9'b111111111;
assign micromatrizz[34][610] = 9'b111111111;
assign micromatrizz[34][611] = 9'b111111111;
assign micromatrizz[34][612] = 9'b111111111;
assign micromatrizz[34][613] = 9'b111111111;
assign micromatrizz[34][614] = 9'b111111111;
assign micromatrizz[34][615] = 9'b111111111;
assign micromatrizz[34][616] = 9'b111111111;
assign micromatrizz[34][617] = 9'b111111111;
assign micromatrizz[34][618] = 9'b111111111;
assign micromatrizz[34][619] = 9'b111111111;
assign micromatrizz[34][620] = 9'b111111111;
assign micromatrizz[34][621] = 9'b111111111;
assign micromatrizz[34][622] = 9'b111111111;
assign micromatrizz[34][623] = 9'b111111111;
assign micromatrizz[34][624] = 9'b111111111;
assign micromatrizz[34][625] = 9'b111111111;
assign micromatrizz[34][626] = 9'b111111111;
assign micromatrizz[34][627] = 9'b111111111;
assign micromatrizz[34][628] = 9'b111111111;
assign micromatrizz[34][629] = 9'b111111111;
assign micromatrizz[34][630] = 9'b111111111;
assign micromatrizz[34][631] = 9'b111111111;
assign micromatrizz[34][632] = 9'b111111111;
assign micromatrizz[34][633] = 9'b111111111;
assign micromatrizz[34][634] = 9'b111111111;
assign micromatrizz[34][635] = 9'b111111111;
assign micromatrizz[34][636] = 9'b111111111;
assign micromatrizz[34][637] = 9'b111111111;
assign micromatrizz[34][638] = 9'b111111111;
assign micromatrizz[34][639] = 9'b111111111;
assign micromatrizz[35][0] = 9'b111111111;
assign micromatrizz[35][1] = 9'b111111111;
assign micromatrizz[35][2] = 9'b111111111;
assign micromatrizz[35][3] = 9'b111111111;
assign micromatrizz[35][4] = 9'b111111111;
assign micromatrizz[35][5] = 9'b111111111;
assign micromatrizz[35][6] = 9'b111111111;
assign micromatrizz[35][7] = 9'b111111111;
assign micromatrizz[35][8] = 9'b111111111;
assign micromatrizz[35][9] = 9'b111111111;
assign micromatrizz[35][10] = 9'b111111111;
assign micromatrizz[35][11] = 9'b111111111;
assign micromatrizz[35][12] = 9'b111111111;
assign micromatrizz[35][13] = 9'b111111111;
assign micromatrizz[35][14] = 9'b111111111;
assign micromatrizz[35][15] = 9'b111111111;
assign micromatrizz[35][16] = 9'b111111111;
assign micromatrizz[35][17] = 9'b111111111;
assign micromatrizz[35][18] = 9'b111111111;
assign micromatrizz[35][19] = 9'b111111111;
assign micromatrizz[35][20] = 9'b111111111;
assign micromatrizz[35][21] = 9'b111111111;
assign micromatrizz[35][22] = 9'b111111111;
assign micromatrizz[35][23] = 9'b111111111;
assign micromatrizz[35][24] = 9'b111111111;
assign micromatrizz[35][25] = 9'b111111111;
assign micromatrizz[35][26] = 9'b111111111;
assign micromatrizz[35][27] = 9'b111111111;
assign micromatrizz[35][28] = 9'b111111111;
assign micromatrizz[35][29] = 9'b111111111;
assign micromatrizz[35][30] = 9'b111111111;
assign micromatrizz[35][31] = 9'b111111111;
assign micromatrizz[35][32] = 9'b111111111;
assign micromatrizz[35][33] = 9'b111111111;
assign micromatrizz[35][34] = 9'b111111111;
assign micromatrizz[35][35] = 9'b111111111;
assign micromatrizz[35][36] = 9'b111111111;
assign micromatrizz[35][37] = 9'b111111111;
assign micromatrizz[35][38] = 9'b111111111;
assign micromatrizz[35][39] = 9'b111111111;
assign micromatrizz[35][40] = 9'b111111111;
assign micromatrizz[35][41] = 9'b111111111;
assign micromatrizz[35][42] = 9'b111111111;
assign micromatrizz[35][43] = 9'b111111111;
assign micromatrizz[35][44] = 9'b111111111;
assign micromatrizz[35][45] = 9'b111111111;
assign micromatrizz[35][46] = 9'b111111111;
assign micromatrizz[35][47] = 9'b111111111;
assign micromatrizz[35][48] = 9'b111111111;
assign micromatrizz[35][49] = 9'b111111111;
assign micromatrizz[35][50] = 9'b111111111;
assign micromatrizz[35][51] = 9'b111111111;
assign micromatrizz[35][52] = 9'b111111111;
assign micromatrizz[35][53] = 9'b111111111;
assign micromatrizz[35][54] = 9'b111111111;
assign micromatrizz[35][55] = 9'b111111111;
assign micromatrizz[35][56] = 9'b111111111;
assign micromatrizz[35][57] = 9'b111111111;
assign micromatrizz[35][58] = 9'b111111111;
assign micromatrizz[35][59] = 9'b111111111;
assign micromatrizz[35][60] = 9'b111111111;
assign micromatrizz[35][61] = 9'b111111111;
assign micromatrizz[35][62] = 9'b111111111;
assign micromatrizz[35][63] = 9'b111111111;
assign micromatrizz[35][64] = 9'b111111111;
assign micromatrizz[35][65] = 9'b111111111;
assign micromatrizz[35][66] = 9'b111111111;
assign micromatrizz[35][67] = 9'b111111111;
assign micromatrizz[35][68] = 9'b111111111;
assign micromatrizz[35][69] = 9'b111111111;
assign micromatrizz[35][70] = 9'b111111111;
assign micromatrizz[35][71] = 9'b111111111;
assign micromatrizz[35][72] = 9'b111111111;
assign micromatrizz[35][73] = 9'b111111111;
assign micromatrizz[35][74] = 9'b111111111;
assign micromatrizz[35][75] = 9'b111111111;
assign micromatrizz[35][76] = 9'b111111111;
assign micromatrizz[35][77] = 9'b111111111;
assign micromatrizz[35][78] = 9'b111111111;
assign micromatrizz[35][79] = 9'b111111111;
assign micromatrizz[35][80] = 9'b111111111;
assign micromatrizz[35][81] = 9'b111111111;
assign micromatrizz[35][82] = 9'b111111111;
assign micromatrizz[35][83] = 9'b111111111;
assign micromatrizz[35][84] = 9'b111111111;
assign micromatrizz[35][85] = 9'b111111111;
assign micromatrizz[35][86] = 9'b111111111;
assign micromatrizz[35][87] = 9'b111111111;
assign micromatrizz[35][88] = 9'b111111111;
assign micromatrizz[35][89] = 9'b111111111;
assign micromatrizz[35][90] = 9'b111111111;
assign micromatrizz[35][91] = 9'b111111111;
assign micromatrizz[35][92] = 9'b111111111;
assign micromatrizz[35][93] = 9'b111111111;
assign micromatrizz[35][94] = 9'b111111111;
assign micromatrizz[35][95] = 9'b111111111;
assign micromatrizz[35][96] = 9'b111111111;
assign micromatrizz[35][97] = 9'b111111111;
assign micromatrizz[35][98] = 9'b111111111;
assign micromatrizz[35][99] = 9'b111111111;
assign micromatrizz[35][100] = 9'b111111111;
assign micromatrizz[35][101] = 9'b111111111;
assign micromatrizz[35][102] = 9'b111111111;
assign micromatrizz[35][103] = 9'b111111111;
assign micromatrizz[35][104] = 9'b111111111;
assign micromatrizz[35][105] = 9'b111111111;
assign micromatrizz[35][106] = 9'b111111111;
assign micromatrizz[35][107] = 9'b111111111;
assign micromatrizz[35][108] = 9'b111111111;
assign micromatrizz[35][109] = 9'b111111111;
assign micromatrizz[35][110] = 9'b111111111;
assign micromatrizz[35][111] = 9'b111111111;
assign micromatrizz[35][112] = 9'b111111111;
assign micromatrizz[35][113] = 9'b111111111;
assign micromatrizz[35][114] = 9'b111111111;
assign micromatrizz[35][115] = 9'b111111111;
assign micromatrizz[35][116] = 9'b111111111;
assign micromatrizz[35][117] = 9'b111111111;
assign micromatrizz[35][118] = 9'b111111111;
assign micromatrizz[35][119] = 9'b111111111;
assign micromatrizz[35][120] = 9'b111111111;
assign micromatrizz[35][121] = 9'b111111111;
assign micromatrizz[35][122] = 9'b111111111;
assign micromatrizz[35][123] = 9'b111111111;
assign micromatrizz[35][124] = 9'b111111111;
assign micromatrizz[35][125] = 9'b111111111;
assign micromatrizz[35][126] = 9'b111111111;
assign micromatrizz[35][127] = 9'b111111111;
assign micromatrizz[35][128] = 9'b111111111;
assign micromatrizz[35][129] = 9'b111111111;
assign micromatrizz[35][130] = 9'b111111111;
assign micromatrizz[35][131] = 9'b111111111;
assign micromatrizz[35][132] = 9'b111111111;
assign micromatrizz[35][133] = 9'b111111111;
assign micromatrizz[35][134] = 9'b111111111;
assign micromatrizz[35][135] = 9'b111111111;
assign micromatrizz[35][136] = 9'b111111111;
assign micromatrizz[35][137] = 9'b111111111;
assign micromatrizz[35][138] = 9'b111111111;
assign micromatrizz[35][139] = 9'b111111111;
assign micromatrizz[35][140] = 9'b111111111;
assign micromatrizz[35][141] = 9'b111111111;
assign micromatrizz[35][142] = 9'b111111111;
assign micromatrizz[35][143] = 9'b111111111;
assign micromatrizz[35][144] = 9'b111111111;
assign micromatrizz[35][145] = 9'b111111111;
assign micromatrizz[35][146] = 9'b111111111;
assign micromatrizz[35][147] = 9'b111111111;
assign micromatrizz[35][148] = 9'b111111111;
assign micromatrizz[35][149] = 9'b111111111;
assign micromatrizz[35][150] = 9'b111111111;
assign micromatrizz[35][151] = 9'b111111111;
assign micromatrizz[35][152] = 9'b111111111;
assign micromatrizz[35][153] = 9'b111111111;
assign micromatrizz[35][154] = 9'b111111111;
assign micromatrizz[35][155] = 9'b111111111;
assign micromatrizz[35][156] = 9'b111111111;
assign micromatrizz[35][157] = 9'b111111111;
assign micromatrizz[35][158] = 9'b111111111;
assign micromatrizz[35][159] = 9'b111111111;
assign micromatrizz[35][160] = 9'b111111111;
assign micromatrizz[35][161] = 9'b111111111;
assign micromatrizz[35][162] = 9'b111111111;
assign micromatrizz[35][163] = 9'b111111111;
assign micromatrizz[35][164] = 9'b111111111;
assign micromatrizz[35][165] = 9'b111111111;
assign micromatrizz[35][166] = 9'b111111111;
assign micromatrizz[35][167] = 9'b111111111;
assign micromatrizz[35][168] = 9'b111111111;
assign micromatrizz[35][169] = 9'b111111111;
assign micromatrizz[35][170] = 9'b111111111;
assign micromatrizz[35][171] = 9'b111111111;
assign micromatrizz[35][172] = 9'b111111111;
assign micromatrizz[35][173] = 9'b111111111;
assign micromatrizz[35][174] = 9'b111111111;
assign micromatrizz[35][175] = 9'b111111111;
assign micromatrizz[35][176] = 9'b111111111;
assign micromatrizz[35][177] = 9'b111111111;
assign micromatrizz[35][178] = 9'b111111111;
assign micromatrizz[35][179] = 9'b111111111;
assign micromatrizz[35][180] = 9'b111111111;
assign micromatrizz[35][181] = 9'b111111111;
assign micromatrizz[35][182] = 9'b111111111;
assign micromatrizz[35][183] = 9'b111111111;
assign micromatrizz[35][184] = 9'b111111111;
assign micromatrizz[35][185] = 9'b111111111;
assign micromatrizz[35][186] = 9'b111111111;
assign micromatrizz[35][187] = 9'b111111111;
assign micromatrizz[35][188] = 9'b111111111;
assign micromatrizz[35][189] = 9'b111111111;
assign micromatrizz[35][190] = 9'b111111111;
assign micromatrizz[35][191] = 9'b111111111;
assign micromatrizz[35][192] = 9'b111111111;
assign micromatrizz[35][193] = 9'b111111111;
assign micromatrizz[35][194] = 9'b111111111;
assign micromatrizz[35][195] = 9'b111111111;
assign micromatrizz[35][196] = 9'b111111111;
assign micromatrizz[35][197] = 9'b111111111;
assign micromatrizz[35][198] = 9'b111111111;
assign micromatrizz[35][199] = 9'b111111111;
assign micromatrizz[35][200] = 9'b111111111;
assign micromatrizz[35][201] = 9'b111111111;
assign micromatrizz[35][202] = 9'b111111111;
assign micromatrizz[35][203] = 9'b111111111;
assign micromatrizz[35][204] = 9'b111111111;
assign micromatrizz[35][205] = 9'b111111111;
assign micromatrizz[35][206] = 9'b111111111;
assign micromatrizz[35][207] = 9'b111111111;
assign micromatrizz[35][208] = 9'b111111111;
assign micromatrizz[35][209] = 9'b111111111;
assign micromatrizz[35][210] = 9'b111111111;
assign micromatrizz[35][211] = 9'b111111111;
assign micromatrizz[35][212] = 9'b111111111;
assign micromatrizz[35][213] = 9'b111111111;
assign micromatrizz[35][214] = 9'b111111111;
assign micromatrizz[35][215] = 9'b111111111;
assign micromatrizz[35][216] = 9'b111111111;
assign micromatrizz[35][217] = 9'b111111111;
assign micromatrizz[35][218] = 9'b111111111;
assign micromatrizz[35][219] = 9'b111111111;
assign micromatrizz[35][220] = 9'b111111111;
assign micromatrizz[35][221] = 9'b111111111;
assign micromatrizz[35][222] = 9'b111111111;
assign micromatrizz[35][223] = 9'b111111111;
assign micromatrizz[35][224] = 9'b111111111;
assign micromatrizz[35][225] = 9'b111111111;
assign micromatrizz[35][226] = 9'b111111111;
assign micromatrizz[35][227] = 9'b111111111;
assign micromatrizz[35][228] = 9'b111111111;
assign micromatrizz[35][229] = 9'b111111111;
assign micromatrizz[35][230] = 9'b111111111;
assign micromatrizz[35][231] = 9'b111111111;
assign micromatrizz[35][232] = 9'b111111111;
assign micromatrizz[35][233] = 9'b111111111;
assign micromatrizz[35][234] = 9'b111111111;
assign micromatrizz[35][235] = 9'b111111111;
assign micromatrizz[35][236] = 9'b111111111;
assign micromatrizz[35][237] = 9'b111111111;
assign micromatrizz[35][238] = 9'b111111111;
assign micromatrizz[35][239] = 9'b111111111;
assign micromatrizz[35][240] = 9'b111111111;
assign micromatrizz[35][241] = 9'b111111111;
assign micromatrizz[35][242] = 9'b111111111;
assign micromatrizz[35][243] = 9'b111111111;
assign micromatrizz[35][244] = 9'b111111111;
assign micromatrizz[35][245] = 9'b111111111;
assign micromatrizz[35][246] = 9'b111111111;
assign micromatrizz[35][247] = 9'b111111111;
assign micromatrizz[35][248] = 9'b111111111;
assign micromatrizz[35][249] = 9'b111111111;
assign micromatrizz[35][250] = 9'b111111111;
assign micromatrizz[35][251] = 9'b111111111;
assign micromatrizz[35][252] = 9'b111111111;
assign micromatrizz[35][253] = 9'b111111111;
assign micromatrizz[35][254] = 9'b111111111;
assign micromatrizz[35][255] = 9'b111111111;
assign micromatrizz[35][256] = 9'b111111111;
assign micromatrizz[35][257] = 9'b111111111;
assign micromatrizz[35][258] = 9'b111111111;
assign micromatrizz[35][259] = 9'b111111111;
assign micromatrizz[35][260] = 9'b111111111;
assign micromatrizz[35][261] = 9'b111111111;
assign micromatrizz[35][262] = 9'b111111111;
assign micromatrizz[35][263] = 9'b111111111;
assign micromatrizz[35][264] = 9'b111111111;
assign micromatrizz[35][265] = 9'b111111111;
assign micromatrizz[35][266] = 9'b111111111;
assign micromatrizz[35][267] = 9'b111111111;
assign micromatrizz[35][268] = 9'b111111111;
assign micromatrizz[35][269] = 9'b111111111;
assign micromatrizz[35][270] = 9'b111110010;
assign micromatrizz[35][271] = 9'b111110010;
assign micromatrizz[35][272] = 9'b111110010;
assign micromatrizz[35][273] = 9'b111110010;
assign micromatrizz[35][274] = 9'b111110010;
assign micromatrizz[35][275] = 9'b111110011;
assign micromatrizz[35][276] = 9'b111110011;
assign micromatrizz[35][277] = 9'b111110011;
assign micromatrizz[35][278] = 9'b111110011;
assign micromatrizz[35][279] = 9'b111111111;
assign micromatrizz[35][280] = 9'b111111111;
assign micromatrizz[35][281] = 9'b111111111;
assign micromatrizz[35][282] = 9'b111111111;
assign micromatrizz[35][283] = 9'b111111111;
assign micromatrizz[35][284] = 9'b111111111;
assign micromatrizz[35][285] = 9'b111111111;
assign micromatrizz[35][286] = 9'b111111111;
assign micromatrizz[35][287] = 9'b111111111;
assign micromatrizz[35][288] = 9'b111111111;
assign micromatrizz[35][289] = 9'b111111111;
assign micromatrizz[35][290] = 9'b111111111;
assign micromatrizz[35][291] = 9'b111111111;
assign micromatrizz[35][292] = 9'b111110011;
assign micromatrizz[35][293] = 9'b111110010;
assign micromatrizz[35][294] = 9'b111110011;
assign micromatrizz[35][295] = 9'b111110011;
assign micromatrizz[35][296] = 9'b111110011;
assign micromatrizz[35][297] = 9'b111110111;
assign micromatrizz[35][298] = 9'b111111111;
assign micromatrizz[35][299] = 9'b111111111;
assign micromatrizz[35][300] = 9'b111111111;
assign micromatrizz[35][301] = 9'b111111111;
assign micromatrizz[35][302] = 9'b111111111;
assign micromatrizz[35][303] = 9'b111110111;
assign micromatrizz[35][304] = 9'b111110111;
assign micromatrizz[35][305] = 9'b111111111;
assign micromatrizz[35][306] = 9'b111111111;
assign micromatrizz[35][307] = 9'b111111111;
assign micromatrizz[35][308] = 9'b111111111;
assign micromatrizz[35][309] = 9'b111111111;
assign micromatrizz[35][310] = 9'b111111111;
assign micromatrizz[35][311] = 9'b111111111;
assign micromatrizz[35][312] = 9'b111111111;
assign micromatrizz[35][313] = 9'b111111111;
assign micromatrizz[35][314] = 9'b111111111;
assign micromatrizz[35][315] = 9'b111110111;
assign micromatrizz[35][316] = 9'b111110010;
assign micromatrizz[35][317] = 9'b111110011;
assign micromatrizz[35][318] = 9'b111110010;
assign micromatrizz[35][319] = 9'b111110010;
assign micromatrizz[35][320] = 9'b111110111;
assign micromatrizz[35][321] = 9'b111111111;
assign micromatrizz[35][322] = 9'b111111111;
assign micromatrizz[35][323] = 9'b111111111;
assign micromatrizz[35][324] = 9'b111111111;
assign micromatrizz[35][325] = 9'b111111111;
assign micromatrizz[35][326] = 9'b111111111;
assign micromatrizz[35][327] = 9'b111111111;
assign micromatrizz[35][328] = 9'b111111111;
assign micromatrizz[35][329] = 9'b111111111;
assign micromatrizz[35][330] = 9'b111111111;
assign micromatrizz[35][331] = 9'b111111111;
assign micromatrizz[35][332] = 9'b111111111;
assign micromatrizz[35][333] = 9'b111111111;
assign micromatrizz[35][334] = 9'b111111111;
assign micromatrizz[35][335] = 9'b111111111;
assign micromatrizz[35][336] = 9'b111111111;
assign micromatrizz[35][337] = 9'b111111111;
assign micromatrizz[35][338] = 9'b111111111;
assign micromatrizz[35][339] = 9'b111111111;
assign micromatrizz[35][340] = 9'b111111111;
assign micromatrizz[35][341] = 9'b111111111;
assign micromatrizz[35][342] = 9'b111111111;
assign micromatrizz[35][343] = 9'b111111111;
assign micromatrizz[35][344] = 9'b111111111;
assign micromatrizz[35][345] = 9'b111111111;
assign micromatrizz[35][346] = 9'b111111111;
assign micromatrizz[35][347] = 9'b111111111;
assign micromatrizz[35][348] = 9'b111111111;
assign micromatrizz[35][349] = 9'b111111111;
assign micromatrizz[35][350] = 9'b111111111;
assign micromatrizz[35][351] = 9'b111111111;
assign micromatrizz[35][352] = 9'b111111111;
assign micromatrizz[35][353] = 9'b111111111;
assign micromatrizz[35][354] = 9'b111111111;
assign micromatrizz[35][355] = 9'b111111111;
assign micromatrizz[35][356] = 9'b111111111;
assign micromatrizz[35][357] = 9'b111111111;
assign micromatrizz[35][358] = 9'b111111111;
assign micromatrizz[35][359] = 9'b111111111;
assign micromatrizz[35][360] = 9'b111111111;
assign micromatrizz[35][361] = 9'b111111111;
assign micromatrizz[35][362] = 9'b111111111;
assign micromatrizz[35][363] = 9'b111111111;
assign micromatrizz[35][364] = 9'b111111111;
assign micromatrizz[35][365] = 9'b111111111;
assign micromatrizz[35][366] = 9'b111111111;
assign micromatrizz[35][367] = 9'b111111111;
assign micromatrizz[35][368] = 9'b111111111;
assign micromatrizz[35][369] = 9'b111111111;
assign micromatrizz[35][370] = 9'b111111111;
assign micromatrizz[35][371] = 9'b111111111;
assign micromatrizz[35][372] = 9'b111111111;
assign micromatrizz[35][373] = 9'b111111111;
assign micromatrizz[35][374] = 9'b111111111;
assign micromatrizz[35][375] = 9'b111111111;
assign micromatrizz[35][376] = 9'b111111111;
assign micromatrizz[35][377] = 9'b111111111;
assign micromatrizz[35][378] = 9'b111111111;
assign micromatrizz[35][379] = 9'b111111111;
assign micromatrizz[35][380] = 9'b111111111;
assign micromatrizz[35][381] = 9'b111111111;
assign micromatrizz[35][382] = 9'b111111111;
assign micromatrizz[35][383] = 9'b111111111;
assign micromatrizz[35][384] = 9'b111111111;
assign micromatrizz[35][385] = 9'b111111111;
assign micromatrizz[35][386] = 9'b111111111;
assign micromatrizz[35][387] = 9'b111111111;
assign micromatrizz[35][388] = 9'b111111111;
assign micromatrizz[35][389] = 9'b111111111;
assign micromatrizz[35][390] = 9'b111111111;
assign micromatrizz[35][391] = 9'b111111111;
assign micromatrizz[35][392] = 9'b111111111;
assign micromatrizz[35][393] = 9'b111111111;
assign micromatrizz[35][394] = 9'b111111111;
assign micromatrizz[35][395] = 9'b111111111;
assign micromatrizz[35][396] = 9'b111111111;
assign micromatrizz[35][397] = 9'b111111111;
assign micromatrizz[35][398] = 9'b111111111;
assign micromatrizz[35][399] = 9'b111111111;
assign micromatrizz[35][400] = 9'b111111111;
assign micromatrizz[35][401] = 9'b111111111;
assign micromatrizz[35][402] = 9'b111111111;
assign micromatrizz[35][403] = 9'b111111111;
assign micromatrizz[35][404] = 9'b111111111;
assign micromatrizz[35][405] = 9'b111111111;
assign micromatrizz[35][406] = 9'b111111111;
assign micromatrizz[35][407] = 9'b111111111;
assign micromatrizz[35][408] = 9'b111111111;
assign micromatrizz[35][409] = 9'b111111111;
assign micromatrizz[35][410] = 9'b111111111;
assign micromatrizz[35][411] = 9'b111111111;
assign micromatrizz[35][412] = 9'b111111111;
assign micromatrizz[35][413] = 9'b111111111;
assign micromatrizz[35][414] = 9'b111111111;
assign micromatrizz[35][415] = 9'b111111111;
assign micromatrizz[35][416] = 9'b111111111;
assign micromatrizz[35][417] = 9'b111111111;
assign micromatrizz[35][418] = 9'b111111111;
assign micromatrizz[35][419] = 9'b111111111;
assign micromatrizz[35][420] = 9'b111111111;
assign micromatrizz[35][421] = 9'b111111111;
assign micromatrizz[35][422] = 9'b111111111;
assign micromatrizz[35][423] = 9'b111111111;
assign micromatrizz[35][424] = 9'b111111111;
assign micromatrizz[35][425] = 9'b111111111;
assign micromatrizz[35][426] = 9'b111111111;
assign micromatrizz[35][427] = 9'b111111111;
assign micromatrizz[35][428] = 9'b111111111;
assign micromatrizz[35][429] = 9'b111111111;
assign micromatrizz[35][430] = 9'b111111111;
assign micromatrizz[35][431] = 9'b111111111;
assign micromatrizz[35][432] = 9'b111111111;
assign micromatrizz[35][433] = 9'b111111111;
assign micromatrizz[35][434] = 9'b111111111;
assign micromatrizz[35][435] = 9'b111111111;
assign micromatrizz[35][436] = 9'b111111111;
assign micromatrizz[35][437] = 9'b111111111;
assign micromatrizz[35][438] = 9'b111111111;
assign micromatrizz[35][439] = 9'b111111111;
assign micromatrizz[35][440] = 9'b111111111;
assign micromatrizz[35][441] = 9'b111111111;
assign micromatrizz[35][442] = 9'b111111111;
assign micromatrizz[35][443] = 9'b111111111;
assign micromatrizz[35][444] = 9'b111111111;
assign micromatrizz[35][445] = 9'b111111111;
assign micromatrizz[35][446] = 9'b111111111;
assign micromatrizz[35][447] = 9'b111111111;
assign micromatrizz[35][448] = 9'b111111111;
assign micromatrizz[35][449] = 9'b111111111;
assign micromatrizz[35][450] = 9'b111111111;
assign micromatrizz[35][451] = 9'b111111111;
assign micromatrizz[35][452] = 9'b111111111;
assign micromatrizz[35][453] = 9'b111111111;
assign micromatrizz[35][454] = 9'b111111111;
assign micromatrizz[35][455] = 9'b111111111;
assign micromatrizz[35][456] = 9'b111111111;
assign micromatrizz[35][457] = 9'b111111111;
assign micromatrizz[35][458] = 9'b111111111;
assign micromatrizz[35][459] = 9'b111111111;
assign micromatrizz[35][460] = 9'b111111111;
assign micromatrizz[35][461] = 9'b111111111;
assign micromatrizz[35][462] = 9'b111111111;
assign micromatrizz[35][463] = 9'b111111111;
assign micromatrizz[35][464] = 9'b111111111;
assign micromatrizz[35][465] = 9'b111111111;
assign micromatrizz[35][466] = 9'b111111111;
assign micromatrizz[35][467] = 9'b111111111;
assign micromatrizz[35][468] = 9'b111111111;
assign micromatrizz[35][469] = 9'b111111111;
assign micromatrizz[35][470] = 9'b111111111;
assign micromatrizz[35][471] = 9'b111111111;
assign micromatrizz[35][472] = 9'b111111111;
assign micromatrizz[35][473] = 9'b111111111;
assign micromatrizz[35][474] = 9'b111111111;
assign micromatrizz[35][475] = 9'b111111111;
assign micromatrizz[35][476] = 9'b111111111;
assign micromatrizz[35][477] = 9'b111111111;
assign micromatrizz[35][478] = 9'b111111111;
assign micromatrizz[35][479] = 9'b111111111;
assign micromatrizz[35][480] = 9'b111111111;
assign micromatrizz[35][481] = 9'b111111111;
assign micromatrizz[35][482] = 9'b111111111;
assign micromatrizz[35][483] = 9'b111111111;
assign micromatrizz[35][484] = 9'b111111111;
assign micromatrizz[35][485] = 9'b111111111;
assign micromatrizz[35][486] = 9'b111111111;
assign micromatrizz[35][487] = 9'b111111111;
assign micromatrizz[35][488] = 9'b111111111;
assign micromatrizz[35][489] = 9'b111111111;
assign micromatrizz[35][490] = 9'b111111111;
assign micromatrizz[35][491] = 9'b111111111;
assign micromatrizz[35][492] = 9'b111111111;
assign micromatrizz[35][493] = 9'b111111111;
assign micromatrizz[35][494] = 9'b111111111;
assign micromatrizz[35][495] = 9'b111111111;
assign micromatrizz[35][496] = 9'b111111111;
assign micromatrizz[35][497] = 9'b111111111;
assign micromatrizz[35][498] = 9'b111111111;
assign micromatrizz[35][499] = 9'b111111111;
assign micromatrizz[35][500] = 9'b111111111;
assign micromatrizz[35][501] = 9'b111111111;
assign micromatrizz[35][502] = 9'b111111111;
assign micromatrizz[35][503] = 9'b111111111;
assign micromatrizz[35][504] = 9'b111111111;
assign micromatrizz[35][505] = 9'b111111111;
assign micromatrizz[35][506] = 9'b111111111;
assign micromatrizz[35][507] = 9'b111111111;
assign micromatrizz[35][508] = 9'b111111111;
assign micromatrizz[35][509] = 9'b111111111;
assign micromatrizz[35][510] = 9'b111111111;
assign micromatrizz[35][511] = 9'b111111111;
assign micromatrizz[35][512] = 9'b111111111;
assign micromatrizz[35][513] = 9'b111111111;
assign micromatrizz[35][514] = 9'b111111111;
assign micromatrizz[35][515] = 9'b111111111;
assign micromatrizz[35][516] = 9'b111111111;
assign micromatrizz[35][517] = 9'b111111111;
assign micromatrizz[35][518] = 9'b111111111;
assign micromatrizz[35][519] = 9'b111111111;
assign micromatrizz[35][520] = 9'b111111111;
assign micromatrizz[35][521] = 9'b111111111;
assign micromatrizz[35][522] = 9'b111111111;
assign micromatrizz[35][523] = 9'b111111111;
assign micromatrizz[35][524] = 9'b111111111;
assign micromatrizz[35][525] = 9'b111111111;
assign micromatrizz[35][526] = 9'b111111111;
assign micromatrizz[35][527] = 9'b111111111;
assign micromatrizz[35][528] = 9'b111111111;
assign micromatrizz[35][529] = 9'b111111111;
assign micromatrizz[35][530] = 9'b111111111;
assign micromatrizz[35][531] = 9'b111111111;
assign micromatrizz[35][532] = 9'b111111111;
assign micromatrizz[35][533] = 9'b111111111;
assign micromatrizz[35][534] = 9'b111111111;
assign micromatrizz[35][535] = 9'b111111111;
assign micromatrizz[35][536] = 9'b111111111;
assign micromatrizz[35][537] = 9'b111111111;
assign micromatrizz[35][538] = 9'b111111111;
assign micromatrizz[35][539] = 9'b111111111;
assign micromatrizz[35][540] = 9'b111111111;
assign micromatrizz[35][541] = 9'b111111111;
assign micromatrizz[35][542] = 9'b111111111;
assign micromatrizz[35][543] = 9'b111111111;
assign micromatrizz[35][544] = 9'b111111111;
assign micromatrizz[35][545] = 9'b111111111;
assign micromatrizz[35][546] = 9'b111111111;
assign micromatrizz[35][547] = 9'b111111111;
assign micromatrizz[35][548] = 9'b111111111;
assign micromatrizz[35][549] = 9'b111111111;
assign micromatrizz[35][550] = 9'b111111111;
assign micromatrizz[35][551] = 9'b111111111;
assign micromatrizz[35][552] = 9'b111111111;
assign micromatrizz[35][553] = 9'b111111111;
assign micromatrizz[35][554] = 9'b111111111;
assign micromatrizz[35][555] = 9'b111111111;
assign micromatrizz[35][556] = 9'b111111111;
assign micromatrizz[35][557] = 9'b111111111;
assign micromatrizz[35][558] = 9'b111111111;
assign micromatrizz[35][559] = 9'b111111111;
assign micromatrizz[35][560] = 9'b111111111;
assign micromatrizz[35][561] = 9'b111111111;
assign micromatrizz[35][562] = 9'b111111111;
assign micromatrizz[35][563] = 9'b111111111;
assign micromatrizz[35][564] = 9'b111111111;
assign micromatrizz[35][565] = 9'b111111111;
assign micromatrizz[35][566] = 9'b111111111;
assign micromatrizz[35][567] = 9'b111111111;
assign micromatrizz[35][568] = 9'b111111111;
assign micromatrizz[35][569] = 9'b111111111;
assign micromatrizz[35][570] = 9'b111111111;
assign micromatrizz[35][571] = 9'b111111111;
assign micromatrizz[35][572] = 9'b111111111;
assign micromatrizz[35][573] = 9'b111111111;
assign micromatrizz[35][574] = 9'b111111111;
assign micromatrizz[35][575] = 9'b111111111;
assign micromatrizz[35][576] = 9'b111111111;
assign micromatrizz[35][577] = 9'b111111111;
assign micromatrizz[35][578] = 9'b111111111;
assign micromatrizz[35][579] = 9'b111111111;
assign micromatrizz[35][580] = 9'b111111111;
assign micromatrizz[35][581] = 9'b111111111;
assign micromatrizz[35][582] = 9'b111111111;
assign micromatrizz[35][583] = 9'b111111111;
assign micromatrizz[35][584] = 9'b111111111;
assign micromatrizz[35][585] = 9'b111111111;
assign micromatrizz[35][586] = 9'b111111111;
assign micromatrizz[35][587] = 9'b111111111;
assign micromatrizz[35][588] = 9'b111111111;
assign micromatrizz[35][589] = 9'b111111111;
assign micromatrizz[35][590] = 9'b111111111;
assign micromatrizz[35][591] = 9'b111111111;
assign micromatrizz[35][592] = 9'b111111111;
assign micromatrizz[35][593] = 9'b111111111;
assign micromatrizz[35][594] = 9'b111111111;
assign micromatrizz[35][595] = 9'b111111111;
assign micromatrizz[35][596] = 9'b111111111;
assign micromatrizz[35][597] = 9'b111111111;
assign micromatrizz[35][598] = 9'b111111111;
assign micromatrizz[35][599] = 9'b111111111;
assign micromatrizz[35][600] = 9'b111111111;
assign micromatrizz[35][601] = 9'b111111111;
assign micromatrizz[35][602] = 9'b111111111;
assign micromatrizz[35][603] = 9'b111111111;
assign micromatrizz[35][604] = 9'b111111111;
assign micromatrizz[35][605] = 9'b111111111;
assign micromatrizz[35][606] = 9'b111111111;
assign micromatrizz[35][607] = 9'b111111111;
assign micromatrizz[35][608] = 9'b111111111;
assign micromatrizz[35][609] = 9'b111111111;
assign micromatrizz[35][610] = 9'b111111111;
assign micromatrizz[35][611] = 9'b111111111;
assign micromatrizz[35][612] = 9'b111111111;
assign micromatrizz[35][613] = 9'b111111111;
assign micromatrizz[35][614] = 9'b111111111;
assign micromatrizz[35][615] = 9'b111111111;
assign micromatrizz[35][616] = 9'b111111111;
assign micromatrizz[35][617] = 9'b111111111;
assign micromatrizz[35][618] = 9'b111111111;
assign micromatrizz[35][619] = 9'b111111111;
assign micromatrizz[35][620] = 9'b111111111;
assign micromatrizz[35][621] = 9'b111111111;
assign micromatrizz[35][622] = 9'b111111111;
assign micromatrizz[35][623] = 9'b111111111;
assign micromatrizz[35][624] = 9'b111111111;
assign micromatrizz[35][625] = 9'b111111111;
assign micromatrizz[35][626] = 9'b111111111;
assign micromatrizz[35][627] = 9'b111111111;
assign micromatrizz[35][628] = 9'b111111111;
assign micromatrizz[35][629] = 9'b111111111;
assign micromatrizz[35][630] = 9'b111111111;
assign micromatrizz[35][631] = 9'b111111111;
assign micromatrizz[35][632] = 9'b111111111;
assign micromatrizz[35][633] = 9'b111111111;
assign micromatrizz[35][634] = 9'b111111111;
assign micromatrizz[35][635] = 9'b111111111;
assign micromatrizz[35][636] = 9'b111111111;
assign micromatrizz[35][637] = 9'b111111111;
assign micromatrizz[35][638] = 9'b111111111;
assign micromatrizz[35][639] = 9'b111111111;
assign micromatrizz[36][0] = 9'b111111111;
assign micromatrizz[36][1] = 9'b111111111;
assign micromatrizz[36][2] = 9'b111111111;
assign micromatrizz[36][3] = 9'b111111111;
assign micromatrizz[36][4] = 9'b111111111;
assign micromatrizz[36][5] = 9'b111111111;
assign micromatrizz[36][6] = 9'b111111111;
assign micromatrizz[36][7] = 9'b111111111;
assign micromatrizz[36][8] = 9'b111111111;
assign micromatrizz[36][9] = 9'b111111111;
assign micromatrizz[36][10] = 9'b111111111;
assign micromatrizz[36][11] = 9'b111111111;
assign micromatrizz[36][12] = 9'b111111111;
assign micromatrizz[36][13] = 9'b111111111;
assign micromatrizz[36][14] = 9'b111111111;
assign micromatrizz[36][15] = 9'b111111111;
assign micromatrizz[36][16] = 9'b111111111;
assign micromatrizz[36][17] = 9'b111111111;
assign micromatrizz[36][18] = 9'b111111111;
assign micromatrizz[36][19] = 9'b111111111;
assign micromatrizz[36][20] = 9'b111111111;
assign micromatrizz[36][21] = 9'b111111111;
assign micromatrizz[36][22] = 9'b111111111;
assign micromatrizz[36][23] = 9'b111111111;
assign micromatrizz[36][24] = 9'b111111111;
assign micromatrizz[36][25] = 9'b111111111;
assign micromatrizz[36][26] = 9'b111111111;
assign micromatrizz[36][27] = 9'b111111111;
assign micromatrizz[36][28] = 9'b111111111;
assign micromatrizz[36][29] = 9'b111111111;
assign micromatrizz[36][30] = 9'b111111111;
assign micromatrizz[36][31] = 9'b111111111;
assign micromatrizz[36][32] = 9'b111111111;
assign micromatrizz[36][33] = 9'b111111111;
assign micromatrizz[36][34] = 9'b111111111;
assign micromatrizz[36][35] = 9'b111111111;
assign micromatrizz[36][36] = 9'b111111111;
assign micromatrizz[36][37] = 9'b111111111;
assign micromatrizz[36][38] = 9'b111111111;
assign micromatrizz[36][39] = 9'b111111111;
assign micromatrizz[36][40] = 9'b111111111;
assign micromatrizz[36][41] = 9'b111111111;
assign micromatrizz[36][42] = 9'b111111111;
assign micromatrizz[36][43] = 9'b111111111;
assign micromatrizz[36][44] = 9'b111111111;
assign micromatrizz[36][45] = 9'b111111111;
assign micromatrizz[36][46] = 9'b111111111;
assign micromatrizz[36][47] = 9'b111111111;
assign micromatrizz[36][48] = 9'b111111111;
assign micromatrizz[36][49] = 9'b111111111;
assign micromatrizz[36][50] = 9'b111111111;
assign micromatrizz[36][51] = 9'b111111111;
assign micromatrizz[36][52] = 9'b111111111;
assign micromatrizz[36][53] = 9'b111111111;
assign micromatrizz[36][54] = 9'b111111111;
assign micromatrizz[36][55] = 9'b111111111;
assign micromatrizz[36][56] = 9'b111111111;
assign micromatrizz[36][57] = 9'b111111111;
assign micromatrizz[36][58] = 9'b111111111;
assign micromatrizz[36][59] = 9'b111111111;
assign micromatrizz[36][60] = 9'b111111111;
assign micromatrizz[36][61] = 9'b111111111;
assign micromatrizz[36][62] = 9'b111111111;
assign micromatrizz[36][63] = 9'b111111111;
assign micromatrizz[36][64] = 9'b111111111;
assign micromatrizz[36][65] = 9'b111111111;
assign micromatrizz[36][66] = 9'b111111111;
assign micromatrizz[36][67] = 9'b111111111;
assign micromatrizz[36][68] = 9'b111111111;
assign micromatrizz[36][69] = 9'b111111111;
assign micromatrizz[36][70] = 9'b111111111;
assign micromatrizz[36][71] = 9'b111111111;
assign micromatrizz[36][72] = 9'b111111111;
assign micromatrizz[36][73] = 9'b111111111;
assign micromatrizz[36][74] = 9'b111111111;
assign micromatrizz[36][75] = 9'b111111111;
assign micromatrizz[36][76] = 9'b111111111;
assign micromatrizz[36][77] = 9'b111111111;
assign micromatrizz[36][78] = 9'b111111111;
assign micromatrizz[36][79] = 9'b111111111;
assign micromatrizz[36][80] = 9'b111111111;
assign micromatrizz[36][81] = 9'b111111111;
assign micromatrizz[36][82] = 9'b111111111;
assign micromatrizz[36][83] = 9'b111111111;
assign micromatrizz[36][84] = 9'b111111111;
assign micromatrizz[36][85] = 9'b111111111;
assign micromatrizz[36][86] = 9'b111111111;
assign micromatrizz[36][87] = 9'b111111111;
assign micromatrizz[36][88] = 9'b111111111;
assign micromatrizz[36][89] = 9'b111111111;
assign micromatrizz[36][90] = 9'b111111111;
assign micromatrizz[36][91] = 9'b111111111;
assign micromatrizz[36][92] = 9'b111111111;
assign micromatrizz[36][93] = 9'b111111111;
assign micromatrizz[36][94] = 9'b111111111;
assign micromatrizz[36][95] = 9'b111111111;
assign micromatrizz[36][96] = 9'b111111111;
assign micromatrizz[36][97] = 9'b111111111;
assign micromatrizz[36][98] = 9'b111111111;
assign micromatrizz[36][99] = 9'b111111111;
assign micromatrizz[36][100] = 9'b111111111;
assign micromatrizz[36][101] = 9'b111111111;
assign micromatrizz[36][102] = 9'b111111111;
assign micromatrizz[36][103] = 9'b111111111;
assign micromatrizz[36][104] = 9'b111111111;
assign micromatrizz[36][105] = 9'b111111111;
assign micromatrizz[36][106] = 9'b111111111;
assign micromatrizz[36][107] = 9'b111111111;
assign micromatrizz[36][108] = 9'b111111111;
assign micromatrizz[36][109] = 9'b111111111;
assign micromatrizz[36][110] = 9'b111111111;
assign micromatrizz[36][111] = 9'b111111111;
assign micromatrizz[36][112] = 9'b111111111;
assign micromatrizz[36][113] = 9'b111111111;
assign micromatrizz[36][114] = 9'b111111111;
assign micromatrizz[36][115] = 9'b111111111;
assign micromatrizz[36][116] = 9'b111111111;
assign micromatrizz[36][117] = 9'b111111111;
assign micromatrizz[36][118] = 9'b111111111;
assign micromatrizz[36][119] = 9'b111111111;
assign micromatrizz[36][120] = 9'b111111111;
assign micromatrizz[36][121] = 9'b111111111;
assign micromatrizz[36][122] = 9'b111111111;
assign micromatrizz[36][123] = 9'b111111111;
assign micromatrizz[36][124] = 9'b111111111;
assign micromatrizz[36][125] = 9'b111111111;
assign micromatrizz[36][126] = 9'b111111111;
assign micromatrizz[36][127] = 9'b111111111;
assign micromatrizz[36][128] = 9'b111111111;
assign micromatrizz[36][129] = 9'b111111111;
assign micromatrizz[36][130] = 9'b111111111;
assign micromatrizz[36][131] = 9'b111111111;
assign micromatrizz[36][132] = 9'b111111111;
assign micromatrizz[36][133] = 9'b111111111;
assign micromatrizz[36][134] = 9'b111111111;
assign micromatrizz[36][135] = 9'b111111111;
assign micromatrizz[36][136] = 9'b111111111;
assign micromatrizz[36][137] = 9'b111111111;
assign micromatrizz[36][138] = 9'b111111111;
assign micromatrizz[36][139] = 9'b111111111;
assign micromatrizz[36][140] = 9'b111111111;
assign micromatrizz[36][141] = 9'b111111111;
assign micromatrizz[36][142] = 9'b111111111;
assign micromatrizz[36][143] = 9'b111111111;
assign micromatrizz[36][144] = 9'b111111111;
assign micromatrizz[36][145] = 9'b111111111;
assign micromatrizz[36][146] = 9'b111111111;
assign micromatrizz[36][147] = 9'b111111111;
assign micromatrizz[36][148] = 9'b111111111;
assign micromatrizz[36][149] = 9'b111111111;
assign micromatrizz[36][150] = 9'b111111111;
assign micromatrizz[36][151] = 9'b111111111;
assign micromatrizz[36][152] = 9'b111111111;
assign micromatrizz[36][153] = 9'b111111111;
assign micromatrizz[36][154] = 9'b111111111;
assign micromatrizz[36][155] = 9'b111111111;
assign micromatrizz[36][156] = 9'b111111111;
assign micromatrizz[36][157] = 9'b111111111;
assign micromatrizz[36][158] = 9'b111111111;
assign micromatrizz[36][159] = 9'b111111111;
assign micromatrizz[36][160] = 9'b111111111;
assign micromatrizz[36][161] = 9'b111111111;
assign micromatrizz[36][162] = 9'b111111111;
assign micromatrizz[36][163] = 9'b111111111;
assign micromatrizz[36][164] = 9'b111111111;
assign micromatrizz[36][165] = 9'b111111111;
assign micromatrizz[36][166] = 9'b111111111;
assign micromatrizz[36][167] = 9'b111111111;
assign micromatrizz[36][168] = 9'b111111111;
assign micromatrizz[36][169] = 9'b111111111;
assign micromatrizz[36][170] = 9'b111111111;
assign micromatrizz[36][171] = 9'b111111111;
assign micromatrizz[36][172] = 9'b111111111;
assign micromatrizz[36][173] = 9'b111111111;
assign micromatrizz[36][174] = 9'b111111111;
assign micromatrizz[36][175] = 9'b111111111;
assign micromatrizz[36][176] = 9'b111111111;
assign micromatrizz[36][177] = 9'b111111111;
assign micromatrizz[36][178] = 9'b111111111;
assign micromatrizz[36][179] = 9'b111111111;
assign micromatrizz[36][180] = 9'b111111111;
assign micromatrizz[36][181] = 9'b111111111;
assign micromatrizz[36][182] = 9'b111111111;
assign micromatrizz[36][183] = 9'b111111111;
assign micromatrizz[36][184] = 9'b111111111;
assign micromatrizz[36][185] = 9'b111111111;
assign micromatrizz[36][186] = 9'b111111111;
assign micromatrizz[36][187] = 9'b111111111;
assign micromatrizz[36][188] = 9'b111111111;
assign micromatrizz[36][189] = 9'b111111111;
assign micromatrizz[36][190] = 9'b111111111;
assign micromatrizz[36][191] = 9'b111111111;
assign micromatrizz[36][192] = 9'b111111111;
assign micromatrizz[36][193] = 9'b111111111;
assign micromatrizz[36][194] = 9'b111111111;
assign micromatrizz[36][195] = 9'b111111111;
assign micromatrizz[36][196] = 9'b111111111;
assign micromatrizz[36][197] = 9'b111111111;
assign micromatrizz[36][198] = 9'b111111111;
assign micromatrizz[36][199] = 9'b111111111;
assign micromatrizz[36][200] = 9'b111111111;
assign micromatrizz[36][201] = 9'b111111111;
assign micromatrizz[36][202] = 9'b111111111;
assign micromatrizz[36][203] = 9'b111111111;
assign micromatrizz[36][204] = 9'b111111111;
assign micromatrizz[36][205] = 9'b111111111;
assign micromatrizz[36][206] = 9'b111111111;
assign micromatrizz[36][207] = 9'b111111111;
assign micromatrizz[36][208] = 9'b111111111;
assign micromatrizz[36][209] = 9'b111111111;
assign micromatrizz[36][210] = 9'b111111111;
assign micromatrizz[36][211] = 9'b111111111;
assign micromatrizz[36][212] = 9'b111111111;
assign micromatrizz[36][213] = 9'b111111111;
assign micromatrizz[36][214] = 9'b111111111;
assign micromatrizz[36][215] = 9'b111111111;
assign micromatrizz[36][216] = 9'b111111111;
assign micromatrizz[36][217] = 9'b111111111;
assign micromatrizz[36][218] = 9'b111111111;
assign micromatrizz[36][219] = 9'b111111111;
assign micromatrizz[36][220] = 9'b111111111;
assign micromatrizz[36][221] = 9'b111111111;
assign micromatrizz[36][222] = 9'b111111111;
assign micromatrizz[36][223] = 9'b111111111;
assign micromatrizz[36][224] = 9'b111111111;
assign micromatrizz[36][225] = 9'b111111111;
assign micromatrizz[36][226] = 9'b111111111;
assign micromatrizz[36][227] = 9'b111111111;
assign micromatrizz[36][228] = 9'b111111111;
assign micromatrizz[36][229] = 9'b111111111;
assign micromatrizz[36][230] = 9'b111111111;
assign micromatrizz[36][231] = 9'b111111111;
assign micromatrizz[36][232] = 9'b111111111;
assign micromatrizz[36][233] = 9'b111111111;
assign micromatrizz[36][234] = 9'b111111111;
assign micromatrizz[36][235] = 9'b111111111;
assign micromatrizz[36][236] = 9'b111111111;
assign micromatrizz[36][237] = 9'b111111111;
assign micromatrizz[36][238] = 9'b111111111;
assign micromatrizz[36][239] = 9'b111111111;
assign micromatrizz[36][240] = 9'b111111111;
assign micromatrizz[36][241] = 9'b111111111;
assign micromatrizz[36][242] = 9'b111111111;
assign micromatrizz[36][243] = 9'b111111111;
assign micromatrizz[36][244] = 9'b111111111;
assign micromatrizz[36][245] = 9'b111111111;
assign micromatrizz[36][246] = 9'b111111111;
assign micromatrizz[36][247] = 9'b111111111;
assign micromatrizz[36][248] = 9'b111111111;
assign micromatrizz[36][249] = 9'b111111111;
assign micromatrizz[36][250] = 9'b111111111;
assign micromatrizz[36][251] = 9'b111111111;
assign micromatrizz[36][252] = 9'b111111111;
assign micromatrizz[36][253] = 9'b111111111;
assign micromatrizz[36][254] = 9'b111111111;
assign micromatrizz[36][255] = 9'b111111111;
assign micromatrizz[36][256] = 9'b111111111;
assign micromatrizz[36][257] = 9'b111111111;
assign micromatrizz[36][258] = 9'b111111111;
assign micromatrizz[36][259] = 9'b111111111;
assign micromatrizz[36][260] = 9'b111111111;
assign micromatrizz[36][261] = 9'b111111111;
assign micromatrizz[36][262] = 9'b111111111;
assign micromatrizz[36][263] = 9'b111111111;
assign micromatrizz[36][264] = 9'b111111111;
assign micromatrizz[36][265] = 9'b111111111;
assign micromatrizz[36][266] = 9'b111111111;
assign micromatrizz[36][267] = 9'b111111111;
assign micromatrizz[36][268] = 9'b111111111;
assign micromatrizz[36][269] = 9'b111111111;
assign micromatrizz[36][270] = 9'b111110010;
assign micromatrizz[36][271] = 9'b111110010;
assign micromatrizz[36][272] = 9'b111110010;
assign micromatrizz[36][273] = 9'b111110010;
assign micromatrizz[36][274] = 9'b111110010;
assign micromatrizz[36][275] = 9'b111110010;
assign micromatrizz[36][276] = 9'b111110011;
assign micromatrizz[36][277] = 9'b111110010;
assign micromatrizz[36][278] = 9'b111110010;
assign micromatrizz[36][279] = 9'b111111111;
assign micromatrizz[36][280] = 9'b111111111;
assign micromatrizz[36][281] = 9'b111111111;
assign micromatrizz[36][282] = 9'b111111111;
assign micromatrizz[36][283] = 9'b111111111;
assign micromatrizz[36][284] = 9'b111111111;
assign micromatrizz[36][285] = 9'b111111111;
assign micromatrizz[36][286] = 9'b111111111;
assign micromatrizz[36][287] = 9'b111111111;
assign micromatrizz[36][288] = 9'b111111111;
assign micromatrizz[36][289] = 9'b111111111;
assign micromatrizz[36][290] = 9'b111111111;
assign micromatrizz[36][291] = 9'b111111111;
assign micromatrizz[36][292] = 9'b111111111;
assign micromatrizz[36][293] = 9'b111111111;
assign micromatrizz[36][294] = 9'b111110111;
assign micromatrizz[36][295] = 9'b111110011;
assign micromatrizz[36][296] = 9'b111110010;
assign micromatrizz[36][297] = 9'b111110111;
assign micromatrizz[36][298] = 9'b111111111;
assign micromatrizz[36][299] = 9'b111111111;
assign micromatrizz[36][300] = 9'b111111111;
assign micromatrizz[36][301] = 9'b111111111;
assign micromatrizz[36][302] = 9'b111111111;
assign micromatrizz[36][303] = 9'b111111111;
assign micromatrizz[36][304] = 9'b111111111;
assign micromatrizz[36][305] = 9'b111111111;
assign micromatrizz[36][306] = 9'b111111111;
assign micromatrizz[36][307] = 9'b111111111;
assign micromatrizz[36][308] = 9'b111111111;
assign micromatrizz[36][309] = 9'b111111111;
assign micromatrizz[36][310] = 9'b111110111;
assign micromatrizz[36][311] = 9'b111110111;
assign micromatrizz[36][312] = 9'b111111111;
assign micromatrizz[36][313] = 9'b111111111;
assign micromatrizz[36][314] = 9'b111111111;
assign micromatrizz[36][315] = 9'b111111111;
assign micromatrizz[36][316] = 9'b111110010;
assign micromatrizz[36][317] = 9'b111110011;
assign micromatrizz[36][318] = 9'b111110011;
assign micromatrizz[36][319] = 9'b111110111;
assign micromatrizz[36][320] = 9'b111111111;
assign micromatrizz[36][321] = 9'b111111111;
assign micromatrizz[36][322] = 9'b111111111;
assign micromatrizz[36][323] = 9'b111111111;
assign micromatrizz[36][324] = 9'b111111111;
assign micromatrizz[36][325] = 9'b111111111;
assign micromatrizz[36][326] = 9'b111111111;
assign micromatrizz[36][327] = 9'b111111111;
assign micromatrizz[36][328] = 9'b111111111;
assign micromatrizz[36][329] = 9'b111111111;
assign micromatrizz[36][330] = 9'b111111111;
assign micromatrizz[36][331] = 9'b111111111;
assign micromatrizz[36][332] = 9'b111111111;
assign micromatrizz[36][333] = 9'b111111111;
assign micromatrizz[36][334] = 9'b111111111;
assign micromatrizz[36][335] = 9'b111111111;
assign micromatrizz[36][336] = 9'b111111111;
assign micromatrizz[36][337] = 9'b111111111;
assign micromatrizz[36][338] = 9'b111111111;
assign micromatrizz[36][339] = 9'b111111111;
assign micromatrizz[36][340] = 9'b111111111;
assign micromatrizz[36][341] = 9'b111111111;
assign micromatrizz[36][342] = 9'b111111111;
assign micromatrizz[36][343] = 9'b111111111;
assign micromatrizz[36][344] = 9'b111111111;
assign micromatrizz[36][345] = 9'b111111111;
assign micromatrizz[36][346] = 9'b111111111;
assign micromatrizz[36][347] = 9'b111111111;
assign micromatrizz[36][348] = 9'b111111111;
assign micromatrizz[36][349] = 9'b111111111;
assign micromatrizz[36][350] = 9'b111111111;
assign micromatrizz[36][351] = 9'b111111111;
assign micromatrizz[36][352] = 9'b111111111;
assign micromatrizz[36][353] = 9'b111111111;
assign micromatrizz[36][354] = 9'b111111111;
assign micromatrizz[36][355] = 9'b111111111;
assign micromatrizz[36][356] = 9'b111111111;
assign micromatrizz[36][357] = 9'b111111111;
assign micromatrizz[36][358] = 9'b111111111;
assign micromatrizz[36][359] = 9'b111111111;
assign micromatrizz[36][360] = 9'b111111111;
assign micromatrizz[36][361] = 9'b111111111;
assign micromatrizz[36][362] = 9'b111111111;
assign micromatrizz[36][363] = 9'b111111111;
assign micromatrizz[36][364] = 9'b111111111;
assign micromatrizz[36][365] = 9'b111111111;
assign micromatrizz[36][366] = 9'b111111111;
assign micromatrizz[36][367] = 9'b111111111;
assign micromatrizz[36][368] = 9'b111111111;
assign micromatrizz[36][369] = 9'b111111111;
assign micromatrizz[36][370] = 9'b111111111;
assign micromatrizz[36][371] = 9'b111111111;
assign micromatrizz[36][372] = 9'b111111111;
assign micromatrizz[36][373] = 9'b111111111;
assign micromatrizz[36][374] = 9'b111111111;
assign micromatrizz[36][375] = 9'b111111111;
assign micromatrizz[36][376] = 9'b111111111;
assign micromatrizz[36][377] = 9'b111111111;
assign micromatrizz[36][378] = 9'b111111111;
assign micromatrizz[36][379] = 9'b111111111;
assign micromatrizz[36][380] = 9'b111111111;
assign micromatrizz[36][381] = 9'b111111111;
assign micromatrizz[36][382] = 9'b111111111;
assign micromatrizz[36][383] = 9'b111111111;
assign micromatrizz[36][384] = 9'b111111111;
assign micromatrizz[36][385] = 9'b111111111;
assign micromatrizz[36][386] = 9'b111111111;
assign micromatrizz[36][387] = 9'b111111111;
assign micromatrizz[36][388] = 9'b111111111;
assign micromatrizz[36][389] = 9'b111111111;
assign micromatrizz[36][390] = 9'b111111111;
assign micromatrizz[36][391] = 9'b111111111;
assign micromatrizz[36][392] = 9'b111111111;
assign micromatrizz[36][393] = 9'b111111111;
assign micromatrizz[36][394] = 9'b111111111;
assign micromatrizz[36][395] = 9'b111111111;
assign micromatrizz[36][396] = 9'b111111111;
assign micromatrizz[36][397] = 9'b111111111;
assign micromatrizz[36][398] = 9'b111111111;
assign micromatrizz[36][399] = 9'b111111111;
assign micromatrizz[36][400] = 9'b111111111;
assign micromatrizz[36][401] = 9'b111111111;
assign micromatrizz[36][402] = 9'b111111111;
assign micromatrizz[36][403] = 9'b111111111;
assign micromatrizz[36][404] = 9'b111111111;
assign micromatrizz[36][405] = 9'b111111111;
assign micromatrizz[36][406] = 9'b111111111;
assign micromatrizz[36][407] = 9'b111111111;
assign micromatrizz[36][408] = 9'b111111111;
assign micromatrizz[36][409] = 9'b111111111;
assign micromatrizz[36][410] = 9'b111111111;
assign micromatrizz[36][411] = 9'b111111111;
assign micromatrizz[36][412] = 9'b111111111;
assign micromatrizz[36][413] = 9'b111111111;
assign micromatrizz[36][414] = 9'b111111111;
assign micromatrizz[36][415] = 9'b111111111;
assign micromatrizz[36][416] = 9'b111111111;
assign micromatrizz[36][417] = 9'b111111111;
assign micromatrizz[36][418] = 9'b111111111;
assign micromatrizz[36][419] = 9'b111111111;
assign micromatrizz[36][420] = 9'b111111111;
assign micromatrizz[36][421] = 9'b111111111;
assign micromatrizz[36][422] = 9'b111111111;
assign micromatrizz[36][423] = 9'b111111111;
assign micromatrizz[36][424] = 9'b111111111;
assign micromatrizz[36][425] = 9'b111111111;
assign micromatrizz[36][426] = 9'b111111111;
assign micromatrizz[36][427] = 9'b111111111;
assign micromatrizz[36][428] = 9'b111111111;
assign micromatrizz[36][429] = 9'b111111111;
assign micromatrizz[36][430] = 9'b111111111;
assign micromatrizz[36][431] = 9'b111111111;
assign micromatrizz[36][432] = 9'b111111111;
assign micromatrizz[36][433] = 9'b111111111;
assign micromatrizz[36][434] = 9'b111111111;
assign micromatrizz[36][435] = 9'b111111111;
assign micromatrizz[36][436] = 9'b111111111;
assign micromatrizz[36][437] = 9'b111111111;
assign micromatrizz[36][438] = 9'b111111111;
assign micromatrizz[36][439] = 9'b111111111;
assign micromatrizz[36][440] = 9'b111111111;
assign micromatrizz[36][441] = 9'b111111111;
assign micromatrizz[36][442] = 9'b111111111;
assign micromatrizz[36][443] = 9'b111111111;
assign micromatrizz[36][444] = 9'b111111111;
assign micromatrizz[36][445] = 9'b111111111;
assign micromatrizz[36][446] = 9'b111111111;
assign micromatrizz[36][447] = 9'b111111111;
assign micromatrizz[36][448] = 9'b111111111;
assign micromatrizz[36][449] = 9'b111111111;
assign micromatrizz[36][450] = 9'b111111111;
assign micromatrizz[36][451] = 9'b111111111;
assign micromatrizz[36][452] = 9'b111111111;
assign micromatrizz[36][453] = 9'b111111111;
assign micromatrizz[36][454] = 9'b111111111;
assign micromatrizz[36][455] = 9'b111111111;
assign micromatrizz[36][456] = 9'b111111111;
assign micromatrizz[36][457] = 9'b111111111;
assign micromatrizz[36][458] = 9'b111111111;
assign micromatrizz[36][459] = 9'b111111111;
assign micromatrizz[36][460] = 9'b111111111;
assign micromatrizz[36][461] = 9'b111111111;
assign micromatrizz[36][462] = 9'b111111111;
assign micromatrizz[36][463] = 9'b111111111;
assign micromatrizz[36][464] = 9'b111111111;
assign micromatrizz[36][465] = 9'b111111111;
assign micromatrizz[36][466] = 9'b111111111;
assign micromatrizz[36][467] = 9'b111111111;
assign micromatrizz[36][468] = 9'b111111111;
assign micromatrizz[36][469] = 9'b111111111;
assign micromatrizz[36][470] = 9'b111111111;
assign micromatrizz[36][471] = 9'b111111111;
assign micromatrizz[36][472] = 9'b111111111;
assign micromatrizz[36][473] = 9'b111111111;
assign micromatrizz[36][474] = 9'b111111111;
assign micromatrizz[36][475] = 9'b111111111;
assign micromatrizz[36][476] = 9'b111111111;
assign micromatrizz[36][477] = 9'b111111111;
assign micromatrizz[36][478] = 9'b111111111;
assign micromatrizz[36][479] = 9'b111111111;
assign micromatrizz[36][480] = 9'b111111111;
assign micromatrizz[36][481] = 9'b111111111;
assign micromatrizz[36][482] = 9'b111111111;
assign micromatrizz[36][483] = 9'b111111111;
assign micromatrizz[36][484] = 9'b111111111;
assign micromatrizz[36][485] = 9'b111111111;
assign micromatrizz[36][486] = 9'b111111111;
assign micromatrizz[36][487] = 9'b111111111;
assign micromatrizz[36][488] = 9'b111111111;
assign micromatrizz[36][489] = 9'b111111111;
assign micromatrizz[36][490] = 9'b111111111;
assign micromatrizz[36][491] = 9'b111111111;
assign micromatrizz[36][492] = 9'b111111111;
assign micromatrizz[36][493] = 9'b111111111;
assign micromatrizz[36][494] = 9'b111111111;
assign micromatrizz[36][495] = 9'b111111111;
assign micromatrizz[36][496] = 9'b111111111;
assign micromatrizz[36][497] = 9'b111111111;
assign micromatrizz[36][498] = 9'b111111111;
assign micromatrizz[36][499] = 9'b111111111;
assign micromatrizz[36][500] = 9'b111111111;
assign micromatrizz[36][501] = 9'b111111111;
assign micromatrizz[36][502] = 9'b111111111;
assign micromatrizz[36][503] = 9'b111111111;
assign micromatrizz[36][504] = 9'b111111111;
assign micromatrizz[36][505] = 9'b111111111;
assign micromatrizz[36][506] = 9'b111111111;
assign micromatrizz[36][507] = 9'b111111111;
assign micromatrizz[36][508] = 9'b111111111;
assign micromatrizz[36][509] = 9'b111111111;
assign micromatrizz[36][510] = 9'b111111111;
assign micromatrizz[36][511] = 9'b111111111;
assign micromatrizz[36][512] = 9'b111111111;
assign micromatrizz[36][513] = 9'b111111111;
assign micromatrizz[36][514] = 9'b111111111;
assign micromatrizz[36][515] = 9'b111111111;
assign micromatrizz[36][516] = 9'b111111111;
assign micromatrizz[36][517] = 9'b111111111;
assign micromatrizz[36][518] = 9'b111111111;
assign micromatrizz[36][519] = 9'b111111111;
assign micromatrizz[36][520] = 9'b111111111;
assign micromatrizz[36][521] = 9'b111111111;
assign micromatrizz[36][522] = 9'b111111111;
assign micromatrizz[36][523] = 9'b111111111;
assign micromatrizz[36][524] = 9'b111111111;
assign micromatrizz[36][525] = 9'b111111111;
assign micromatrizz[36][526] = 9'b111111111;
assign micromatrizz[36][527] = 9'b111111111;
assign micromatrizz[36][528] = 9'b111111111;
assign micromatrizz[36][529] = 9'b111111111;
assign micromatrizz[36][530] = 9'b111111111;
assign micromatrizz[36][531] = 9'b111111111;
assign micromatrizz[36][532] = 9'b111111111;
assign micromatrizz[36][533] = 9'b111111111;
assign micromatrizz[36][534] = 9'b111111111;
assign micromatrizz[36][535] = 9'b111111111;
assign micromatrizz[36][536] = 9'b111111111;
assign micromatrizz[36][537] = 9'b111111111;
assign micromatrizz[36][538] = 9'b111111111;
assign micromatrizz[36][539] = 9'b111111111;
assign micromatrizz[36][540] = 9'b111111111;
assign micromatrizz[36][541] = 9'b111111111;
assign micromatrizz[36][542] = 9'b111111111;
assign micromatrizz[36][543] = 9'b111111111;
assign micromatrizz[36][544] = 9'b111111111;
assign micromatrizz[36][545] = 9'b111111111;
assign micromatrizz[36][546] = 9'b111111111;
assign micromatrizz[36][547] = 9'b111111111;
assign micromatrizz[36][548] = 9'b111111111;
assign micromatrizz[36][549] = 9'b111111111;
assign micromatrizz[36][550] = 9'b111111111;
assign micromatrizz[36][551] = 9'b111111111;
assign micromatrizz[36][552] = 9'b111111111;
assign micromatrizz[36][553] = 9'b111111111;
assign micromatrizz[36][554] = 9'b111111111;
assign micromatrizz[36][555] = 9'b111111111;
assign micromatrizz[36][556] = 9'b111111111;
assign micromatrizz[36][557] = 9'b111111111;
assign micromatrizz[36][558] = 9'b111111111;
assign micromatrizz[36][559] = 9'b111111111;
assign micromatrizz[36][560] = 9'b111111111;
assign micromatrizz[36][561] = 9'b111111111;
assign micromatrizz[36][562] = 9'b111111111;
assign micromatrizz[36][563] = 9'b111111111;
assign micromatrizz[36][564] = 9'b111111111;
assign micromatrizz[36][565] = 9'b111111111;
assign micromatrizz[36][566] = 9'b111111111;
assign micromatrizz[36][567] = 9'b111111111;
assign micromatrizz[36][568] = 9'b111111111;
assign micromatrizz[36][569] = 9'b111111111;
assign micromatrizz[36][570] = 9'b111111111;
assign micromatrizz[36][571] = 9'b111111111;
assign micromatrizz[36][572] = 9'b111111111;
assign micromatrizz[36][573] = 9'b111111111;
assign micromatrizz[36][574] = 9'b111111111;
assign micromatrizz[36][575] = 9'b111111111;
assign micromatrizz[36][576] = 9'b111111111;
assign micromatrizz[36][577] = 9'b111111111;
assign micromatrizz[36][578] = 9'b111111111;
assign micromatrizz[36][579] = 9'b111111111;
assign micromatrizz[36][580] = 9'b111111111;
assign micromatrizz[36][581] = 9'b111111111;
assign micromatrizz[36][582] = 9'b111111111;
assign micromatrizz[36][583] = 9'b111111111;
assign micromatrizz[36][584] = 9'b111111111;
assign micromatrizz[36][585] = 9'b111111111;
assign micromatrizz[36][586] = 9'b111111111;
assign micromatrizz[36][587] = 9'b111111111;
assign micromatrizz[36][588] = 9'b111111111;
assign micromatrizz[36][589] = 9'b111111111;
assign micromatrizz[36][590] = 9'b111111111;
assign micromatrizz[36][591] = 9'b111111111;
assign micromatrizz[36][592] = 9'b111111111;
assign micromatrizz[36][593] = 9'b111111111;
assign micromatrizz[36][594] = 9'b111111111;
assign micromatrizz[36][595] = 9'b111111111;
assign micromatrizz[36][596] = 9'b111111111;
assign micromatrizz[36][597] = 9'b111111111;
assign micromatrizz[36][598] = 9'b111111111;
assign micromatrizz[36][599] = 9'b111111111;
assign micromatrizz[36][600] = 9'b111111111;
assign micromatrizz[36][601] = 9'b111111111;
assign micromatrizz[36][602] = 9'b111111111;
assign micromatrizz[36][603] = 9'b111111111;
assign micromatrizz[36][604] = 9'b111111111;
assign micromatrizz[36][605] = 9'b111111111;
assign micromatrizz[36][606] = 9'b111111111;
assign micromatrizz[36][607] = 9'b111111111;
assign micromatrizz[36][608] = 9'b111111111;
assign micromatrizz[36][609] = 9'b111111111;
assign micromatrizz[36][610] = 9'b111111111;
assign micromatrizz[36][611] = 9'b111111111;
assign micromatrizz[36][612] = 9'b111111111;
assign micromatrizz[36][613] = 9'b111111111;
assign micromatrizz[36][614] = 9'b111111111;
assign micromatrizz[36][615] = 9'b111111111;
assign micromatrizz[36][616] = 9'b111111111;
assign micromatrizz[36][617] = 9'b111111111;
assign micromatrizz[36][618] = 9'b111111111;
assign micromatrizz[36][619] = 9'b111111111;
assign micromatrizz[36][620] = 9'b111111111;
assign micromatrizz[36][621] = 9'b111111111;
assign micromatrizz[36][622] = 9'b111111111;
assign micromatrizz[36][623] = 9'b111111111;
assign micromatrizz[36][624] = 9'b111111111;
assign micromatrizz[36][625] = 9'b111111111;
assign micromatrizz[36][626] = 9'b111111111;
assign micromatrizz[36][627] = 9'b111111111;
assign micromatrizz[36][628] = 9'b111111111;
assign micromatrizz[36][629] = 9'b111111111;
assign micromatrizz[36][630] = 9'b111111111;
assign micromatrizz[36][631] = 9'b111111111;
assign micromatrizz[36][632] = 9'b111111111;
assign micromatrizz[36][633] = 9'b111111111;
assign micromatrizz[36][634] = 9'b111111111;
assign micromatrizz[36][635] = 9'b111111111;
assign micromatrizz[36][636] = 9'b111111111;
assign micromatrizz[36][637] = 9'b111111111;
assign micromatrizz[36][638] = 9'b111111111;
assign micromatrizz[36][639] = 9'b111111111;
assign micromatrizz[37][0] = 9'b111111111;
assign micromatrizz[37][1] = 9'b111111111;
assign micromatrizz[37][2] = 9'b111111111;
assign micromatrizz[37][3] = 9'b111111111;
assign micromatrizz[37][4] = 9'b111111111;
assign micromatrizz[37][5] = 9'b111111111;
assign micromatrizz[37][6] = 9'b111111111;
assign micromatrizz[37][7] = 9'b111111111;
assign micromatrizz[37][8] = 9'b111111111;
assign micromatrizz[37][9] = 9'b111111111;
assign micromatrizz[37][10] = 9'b111111111;
assign micromatrizz[37][11] = 9'b111111111;
assign micromatrizz[37][12] = 9'b111111111;
assign micromatrizz[37][13] = 9'b111111111;
assign micromatrizz[37][14] = 9'b111111111;
assign micromatrizz[37][15] = 9'b111111111;
assign micromatrizz[37][16] = 9'b111111111;
assign micromatrizz[37][17] = 9'b111111111;
assign micromatrizz[37][18] = 9'b111111111;
assign micromatrizz[37][19] = 9'b111111111;
assign micromatrizz[37][20] = 9'b111111111;
assign micromatrizz[37][21] = 9'b111111111;
assign micromatrizz[37][22] = 9'b111111111;
assign micromatrizz[37][23] = 9'b111111111;
assign micromatrizz[37][24] = 9'b111111111;
assign micromatrizz[37][25] = 9'b111111111;
assign micromatrizz[37][26] = 9'b111111111;
assign micromatrizz[37][27] = 9'b111111111;
assign micromatrizz[37][28] = 9'b111111111;
assign micromatrizz[37][29] = 9'b111111111;
assign micromatrizz[37][30] = 9'b111111111;
assign micromatrizz[37][31] = 9'b111111111;
assign micromatrizz[37][32] = 9'b111111111;
assign micromatrizz[37][33] = 9'b111111111;
assign micromatrizz[37][34] = 9'b111111111;
assign micromatrizz[37][35] = 9'b111111111;
assign micromatrizz[37][36] = 9'b111111111;
assign micromatrizz[37][37] = 9'b111111111;
assign micromatrizz[37][38] = 9'b111111111;
assign micromatrizz[37][39] = 9'b111111111;
assign micromatrizz[37][40] = 9'b111111111;
assign micromatrizz[37][41] = 9'b111111111;
assign micromatrizz[37][42] = 9'b111111111;
assign micromatrizz[37][43] = 9'b111111111;
assign micromatrizz[37][44] = 9'b111111111;
assign micromatrizz[37][45] = 9'b111111111;
assign micromatrizz[37][46] = 9'b111111111;
assign micromatrizz[37][47] = 9'b111111111;
assign micromatrizz[37][48] = 9'b111111111;
assign micromatrizz[37][49] = 9'b111111111;
assign micromatrizz[37][50] = 9'b111111111;
assign micromatrizz[37][51] = 9'b111111111;
assign micromatrizz[37][52] = 9'b111111111;
assign micromatrizz[37][53] = 9'b111111111;
assign micromatrizz[37][54] = 9'b111111111;
assign micromatrizz[37][55] = 9'b111111111;
assign micromatrizz[37][56] = 9'b111111111;
assign micromatrizz[37][57] = 9'b111111111;
assign micromatrizz[37][58] = 9'b111111111;
assign micromatrizz[37][59] = 9'b111111111;
assign micromatrizz[37][60] = 9'b111111111;
assign micromatrizz[37][61] = 9'b111111111;
assign micromatrizz[37][62] = 9'b111111111;
assign micromatrizz[37][63] = 9'b111111111;
assign micromatrizz[37][64] = 9'b111111111;
assign micromatrizz[37][65] = 9'b111111111;
assign micromatrizz[37][66] = 9'b111111111;
assign micromatrizz[37][67] = 9'b111111111;
assign micromatrizz[37][68] = 9'b111111111;
assign micromatrizz[37][69] = 9'b111111111;
assign micromatrizz[37][70] = 9'b111111111;
assign micromatrizz[37][71] = 9'b111111111;
assign micromatrizz[37][72] = 9'b111111111;
assign micromatrizz[37][73] = 9'b111111111;
assign micromatrizz[37][74] = 9'b111111111;
assign micromatrizz[37][75] = 9'b111111111;
assign micromatrizz[37][76] = 9'b111111111;
assign micromatrizz[37][77] = 9'b111111111;
assign micromatrizz[37][78] = 9'b111111111;
assign micromatrizz[37][79] = 9'b111111111;
assign micromatrizz[37][80] = 9'b111111111;
assign micromatrizz[37][81] = 9'b111111111;
assign micromatrizz[37][82] = 9'b111111111;
assign micromatrizz[37][83] = 9'b111111111;
assign micromatrizz[37][84] = 9'b111111111;
assign micromatrizz[37][85] = 9'b111111111;
assign micromatrizz[37][86] = 9'b111111111;
assign micromatrizz[37][87] = 9'b111111111;
assign micromatrizz[37][88] = 9'b111111111;
assign micromatrizz[37][89] = 9'b111111111;
assign micromatrizz[37][90] = 9'b111111111;
assign micromatrizz[37][91] = 9'b111111111;
assign micromatrizz[37][92] = 9'b111111111;
assign micromatrizz[37][93] = 9'b111111111;
assign micromatrizz[37][94] = 9'b111111111;
assign micromatrizz[37][95] = 9'b111111111;
assign micromatrizz[37][96] = 9'b111111111;
assign micromatrizz[37][97] = 9'b111111111;
assign micromatrizz[37][98] = 9'b111111111;
assign micromatrizz[37][99] = 9'b111111111;
assign micromatrizz[37][100] = 9'b111111111;
assign micromatrizz[37][101] = 9'b111111111;
assign micromatrizz[37][102] = 9'b111111111;
assign micromatrizz[37][103] = 9'b111111111;
assign micromatrizz[37][104] = 9'b111111111;
assign micromatrizz[37][105] = 9'b111111111;
assign micromatrizz[37][106] = 9'b111111111;
assign micromatrizz[37][107] = 9'b111111111;
assign micromatrizz[37][108] = 9'b111111111;
assign micromatrizz[37][109] = 9'b111111111;
assign micromatrizz[37][110] = 9'b111111111;
assign micromatrizz[37][111] = 9'b111111111;
assign micromatrizz[37][112] = 9'b111111111;
assign micromatrizz[37][113] = 9'b111111111;
assign micromatrizz[37][114] = 9'b111111111;
assign micromatrizz[37][115] = 9'b111111111;
assign micromatrizz[37][116] = 9'b111111111;
assign micromatrizz[37][117] = 9'b111111111;
assign micromatrizz[37][118] = 9'b111111111;
assign micromatrizz[37][119] = 9'b111111111;
assign micromatrizz[37][120] = 9'b111111111;
assign micromatrizz[37][121] = 9'b111111111;
assign micromatrizz[37][122] = 9'b111111111;
assign micromatrizz[37][123] = 9'b111111111;
assign micromatrizz[37][124] = 9'b111111111;
assign micromatrizz[37][125] = 9'b111111111;
assign micromatrizz[37][126] = 9'b111111111;
assign micromatrizz[37][127] = 9'b111111111;
assign micromatrizz[37][128] = 9'b111111111;
assign micromatrizz[37][129] = 9'b111111111;
assign micromatrizz[37][130] = 9'b111111111;
assign micromatrizz[37][131] = 9'b111111111;
assign micromatrizz[37][132] = 9'b111111111;
assign micromatrizz[37][133] = 9'b111111111;
assign micromatrizz[37][134] = 9'b111111111;
assign micromatrizz[37][135] = 9'b111111111;
assign micromatrizz[37][136] = 9'b111111111;
assign micromatrizz[37][137] = 9'b111111111;
assign micromatrizz[37][138] = 9'b111111111;
assign micromatrizz[37][139] = 9'b111111111;
assign micromatrizz[37][140] = 9'b111111111;
assign micromatrizz[37][141] = 9'b111111111;
assign micromatrizz[37][142] = 9'b111111111;
assign micromatrizz[37][143] = 9'b111111111;
assign micromatrizz[37][144] = 9'b111111111;
assign micromatrizz[37][145] = 9'b111111111;
assign micromatrizz[37][146] = 9'b111111111;
assign micromatrizz[37][147] = 9'b111111111;
assign micromatrizz[37][148] = 9'b111111111;
assign micromatrizz[37][149] = 9'b111111111;
assign micromatrizz[37][150] = 9'b111111111;
assign micromatrizz[37][151] = 9'b111111111;
assign micromatrizz[37][152] = 9'b111111111;
assign micromatrizz[37][153] = 9'b111111111;
assign micromatrizz[37][154] = 9'b111111111;
assign micromatrizz[37][155] = 9'b111111111;
assign micromatrizz[37][156] = 9'b111111111;
assign micromatrizz[37][157] = 9'b111111111;
assign micromatrizz[37][158] = 9'b111111111;
assign micromatrizz[37][159] = 9'b111111111;
assign micromatrizz[37][160] = 9'b111111111;
assign micromatrizz[37][161] = 9'b111111111;
assign micromatrizz[37][162] = 9'b111111111;
assign micromatrizz[37][163] = 9'b111111111;
assign micromatrizz[37][164] = 9'b111111111;
assign micromatrizz[37][165] = 9'b111111111;
assign micromatrizz[37][166] = 9'b111111111;
assign micromatrizz[37][167] = 9'b111111111;
assign micromatrizz[37][168] = 9'b111111111;
assign micromatrizz[37][169] = 9'b111111111;
assign micromatrizz[37][170] = 9'b111111111;
assign micromatrizz[37][171] = 9'b111111111;
assign micromatrizz[37][172] = 9'b111111111;
assign micromatrizz[37][173] = 9'b111111111;
assign micromatrizz[37][174] = 9'b111111111;
assign micromatrizz[37][175] = 9'b111111111;
assign micromatrizz[37][176] = 9'b111111111;
assign micromatrizz[37][177] = 9'b111111111;
assign micromatrizz[37][178] = 9'b111111111;
assign micromatrizz[37][179] = 9'b111111111;
assign micromatrizz[37][180] = 9'b111111111;
assign micromatrizz[37][181] = 9'b111111111;
assign micromatrizz[37][182] = 9'b111111111;
assign micromatrizz[37][183] = 9'b111111111;
assign micromatrizz[37][184] = 9'b111111111;
assign micromatrizz[37][185] = 9'b111111111;
assign micromatrizz[37][186] = 9'b111111111;
assign micromatrizz[37][187] = 9'b111111111;
assign micromatrizz[37][188] = 9'b111111111;
assign micromatrizz[37][189] = 9'b111111111;
assign micromatrizz[37][190] = 9'b111111111;
assign micromatrizz[37][191] = 9'b111111111;
assign micromatrizz[37][192] = 9'b111111111;
assign micromatrizz[37][193] = 9'b111111111;
assign micromatrizz[37][194] = 9'b111111111;
assign micromatrizz[37][195] = 9'b111111111;
assign micromatrizz[37][196] = 9'b111111111;
assign micromatrizz[37][197] = 9'b111111111;
assign micromatrizz[37][198] = 9'b111111111;
assign micromatrizz[37][199] = 9'b111111111;
assign micromatrizz[37][200] = 9'b111111111;
assign micromatrizz[37][201] = 9'b111111111;
assign micromatrizz[37][202] = 9'b111111111;
assign micromatrizz[37][203] = 9'b111111111;
assign micromatrizz[37][204] = 9'b111111111;
assign micromatrizz[37][205] = 9'b111111111;
assign micromatrizz[37][206] = 9'b111111111;
assign micromatrizz[37][207] = 9'b111111111;
assign micromatrizz[37][208] = 9'b111111111;
assign micromatrizz[37][209] = 9'b111111111;
assign micromatrizz[37][210] = 9'b111111111;
assign micromatrizz[37][211] = 9'b111111111;
assign micromatrizz[37][212] = 9'b111111111;
assign micromatrizz[37][213] = 9'b111111111;
assign micromatrizz[37][214] = 9'b111111111;
assign micromatrizz[37][215] = 9'b111111111;
assign micromatrizz[37][216] = 9'b111111111;
assign micromatrizz[37][217] = 9'b111111111;
assign micromatrizz[37][218] = 9'b111111111;
assign micromatrizz[37][219] = 9'b111111111;
assign micromatrizz[37][220] = 9'b111111111;
assign micromatrizz[37][221] = 9'b111111111;
assign micromatrizz[37][222] = 9'b111111111;
assign micromatrizz[37][223] = 9'b111111111;
assign micromatrizz[37][224] = 9'b111111111;
assign micromatrizz[37][225] = 9'b111111111;
assign micromatrizz[37][226] = 9'b111111111;
assign micromatrizz[37][227] = 9'b111111111;
assign micromatrizz[37][228] = 9'b111111111;
assign micromatrizz[37][229] = 9'b111111111;
assign micromatrizz[37][230] = 9'b111111111;
assign micromatrizz[37][231] = 9'b111111111;
assign micromatrizz[37][232] = 9'b111111111;
assign micromatrizz[37][233] = 9'b111111111;
assign micromatrizz[37][234] = 9'b111111111;
assign micromatrizz[37][235] = 9'b111111111;
assign micromatrizz[37][236] = 9'b111111111;
assign micromatrizz[37][237] = 9'b111111111;
assign micromatrizz[37][238] = 9'b111111111;
assign micromatrizz[37][239] = 9'b111111111;
assign micromatrizz[37][240] = 9'b111111111;
assign micromatrizz[37][241] = 9'b111111111;
assign micromatrizz[37][242] = 9'b111111111;
assign micromatrizz[37][243] = 9'b111111111;
assign micromatrizz[37][244] = 9'b111111111;
assign micromatrizz[37][245] = 9'b111111111;
assign micromatrizz[37][246] = 9'b111111111;
assign micromatrizz[37][247] = 9'b111111111;
assign micromatrizz[37][248] = 9'b111111111;
assign micromatrizz[37][249] = 9'b111111111;
assign micromatrizz[37][250] = 9'b111111111;
assign micromatrizz[37][251] = 9'b111111111;
assign micromatrizz[37][252] = 9'b111111111;
assign micromatrizz[37][253] = 9'b111111111;
assign micromatrizz[37][254] = 9'b111111111;
assign micromatrizz[37][255] = 9'b111111111;
assign micromatrizz[37][256] = 9'b111111111;
assign micromatrizz[37][257] = 9'b111111111;
assign micromatrizz[37][258] = 9'b111111111;
assign micromatrizz[37][259] = 9'b111111111;
assign micromatrizz[37][260] = 9'b111111111;
assign micromatrizz[37][261] = 9'b111111111;
assign micromatrizz[37][262] = 9'b111111111;
assign micromatrizz[37][263] = 9'b111111111;
assign micromatrizz[37][264] = 9'b111111111;
assign micromatrizz[37][265] = 9'b111111111;
assign micromatrizz[37][266] = 9'b111111111;
assign micromatrizz[37][267] = 9'b111111111;
assign micromatrizz[37][268] = 9'b111111111;
assign micromatrizz[37][269] = 9'b111111111;
assign micromatrizz[37][270] = 9'b111110111;
assign micromatrizz[37][271] = 9'b111110111;
assign micromatrizz[37][272] = 9'b111110111;
assign micromatrizz[37][273] = 9'b111110111;
assign micromatrizz[37][274] = 9'b111110111;
assign micromatrizz[37][275] = 9'b111110111;
assign micromatrizz[37][276] = 9'b111110111;
assign micromatrizz[37][277] = 9'b111110111;
assign micromatrizz[37][278] = 9'b111110111;
assign micromatrizz[37][279] = 9'b111110111;
assign micromatrizz[37][280] = 9'b111111111;
assign micromatrizz[37][281] = 9'b111111111;
assign micromatrizz[37][282] = 9'b111111111;
assign micromatrizz[37][283] = 9'b111111111;
assign micromatrizz[37][284] = 9'b111110111;
assign micromatrizz[37][285] = 9'b111110111;
assign micromatrizz[37][286] = 9'b111111111;
assign micromatrizz[37][287] = 9'b111111111;
assign micromatrizz[37][288] = 9'b111111111;
assign micromatrizz[37][289] = 9'b111111111;
assign micromatrizz[37][290] = 9'b111111111;
assign micromatrizz[37][291] = 9'b111111111;
assign micromatrizz[37][292] = 9'b111111111;
assign micromatrizz[37][293] = 9'b111111111;
assign micromatrizz[37][294] = 9'b111111111;
assign micromatrizz[37][295] = 9'b111111111;
assign micromatrizz[37][296] = 9'b111110111;
assign micromatrizz[37][297] = 9'b111110111;
assign micromatrizz[37][298] = 9'b111110111;
assign micromatrizz[37][299] = 9'b111110111;
assign micromatrizz[37][300] = 9'b111111111;
assign micromatrizz[37][301] = 9'b111111111;
assign micromatrizz[37][302] = 9'b111111111;
assign micromatrizz[37][303] = 9'b111111111;
assign micromatrizz[37][304] = 9'b111111111;
assign micromatrizz[37][305] = 9'b111111111;
assign micromatrizz[37][306] = 9'b111111111;
assign micromatrizz[37][307] = 9'b111111111;
assign micromatrizz[37][308] = 9'b111111111;
assign micromatrizz[37][309] = 9'b111111111;
assign micromatrizz[37][310] = 9'b111111111;
assign micromatrizz[37][311] = 9'b111111111;
assign micromatrizz[37][312] = 9'b111111111;
assign micromatrizz[37][313] = 9'b111110111;
assign micromatrizz[37][314] = 9'b111110111;
assign micromatrizz[37][315] = 9'b111110111;
assign micromatrizz[37][316] = 9'b111110111;
assign micromatrizz[37][317] = 9'b111111111;
assign micromatrizz[37][318] = 9'b111111111;
assign micromatrizz[37][319] = 9'b111111111;
assign micromatrizz[37][320] = 9'b111111111;
assign micromatrizz[37][321] = 9'b111111111;
assign micromatrizz[37][322] = 9'b111111111;
assign micromatrizz[37][323] = 9'b111111111;
assign micromatrizz[37][324] = 9'b111111111;
assign micromatrizz[37][325] = 9'b111111111;
assign micromatrizz[37][326] = 9'b111111111;
assign micromatrizz[37][327] = 9'b111111111;
assign micromatrizz[37][328] = 9'b111111111;
assign micromatrizz[37][329] = 9'b111111111;
assign micromatrizz[37][330] = 9'b111111111;
assign micromatrizz[37][331] = 9'b111111111;
assign micromatrizz[37][332] = 9'b111111111;
assign micromatrizz[37][333] = 9'b111111111;
assign micromatrizz[37][334] = 9'b111111111;
assign micromatrizz[37][335] = 9'b111111111;
assign micromatrizz[37][336] = 9'b111111111;
assign micromatrizz[37][337] = 9'b111111111;
assign micromatrizz[37][338] = 9'b111111111;
assign micromatrizz[37][339] = 9'b111111111;
assign micromatrizz[37][340] = 9'b111111111;
assign micromatrizz[37][341] = 9'b111111111;
assign micromatrizz[37][342] = 9'b111111111;
assign micromatrizz[37][343] = 9'b111111111;
assign micromatrizz[37][344] = 9'b111111111;
assign micromatrizz[37][345] = 9'b111111111;
assign micromatrizz[37][346] = 9'b111111111;
assign micromatrizz[37][347] = 9'b111111111;
assign micromatrizz[37][348] = 9'b111111111;
assign micromatrizz[37][349] = 9'b111111111;
assign micromatrizz[37][350] = 9'b111111111;
assign micromatrizz[37][351] = 9'b111111111;
assign micromatrizz[37][352] = 9'b111111111;
assign micromatrizz[37][353] = 9'b111111111;
assign micromatrizz[37][354] = 9'b111111111;
assign micromatrizz[37][355] = 9'b111111111;
assign micromatrizz[37][356] = 9'b111111111;
assign micromatrizz[37][357] = 9'b111111111;
assign micromatrizz[37][358] = 9'b111111111;
assign micromatrizz[37][359] = 9'b111111111;
assign micromatrizz[37][360] = 9'b111111111;
assign micromatrizz[37][361] = 9'b111111111;
assign micromatrizz[37][362] = 9'b111111111;
assign micromatrizz[37][363] = 9'b111111111;
assign micromatrizz[37][364] = 9'b111111111;
assign micromatrizz[37][365] = 9'b111111111;
assign micromatrizz[37][366] = 9'b111111111;
assign micromatrizz[37][367] = 9'b111111111;
assign micromatrizz[37][368] = 9'b111111111;
assign micromatrizz[37][369] = 9'b111111111;
assign micromatrizz[37][370] = 9'b111111111;
assign micromatrizz[37][371] = 9'b111111111;
assign micromatrizz[37][372] = 9'b111111111;
assign micromatrizz[37][373] = 9'b111111111;
assign micromatrizz[37][374] = 9'b111111111;
assign micromatrizz[37][375] = 9'b111111111;
assign micromatrizz[37][376] = 9'b111111111;
assign micromatrizz[37][377] = 9'b111111111;
assign micromatrizz[37][378] = 9'b111111111;
assign micromatrizz[37][379] = 9'b111111111;
assign micromatrizz[37][380] = 9'b111111111;
assign micromatrizz[37][381] = 9'b111111111;
assign micromatrizz[37][382] = 9'b111111111;
assign micromatrizz[37][383] = 9'b111111111;
assign micromatrizz[37][384] = 9'b111111111;
assign micromatrizz[37][385] = 9'b111111111;
assign micromatrizz[37][386] = 9'b111111111;
assign micromatrizz[37][387] = 9'b111111111;
assign micromatrizz[37][388] = 9'b111111111;
assign micromatrizz[37][389] = 9'b111111111;
assign micromatrizz[37][390] = 9'b111111111;
assign micromatrizz[37][391] = 9'b111111111;
assign micromatrizz[37][392] = 9'b111111111;
assign micromatrizz[37][393] = 9'b111111111;
assign micromatrizz[37][394] = 9'b111111111;
assign micromatrizz[37][395] = 9'b111111111;
assign micromatrizz[37][396] = 9'b111111111;
assign micromatrizz[37][397] = 9'b111111111;
assign micromatrizz[37][398] = 9'b111111111;
assign micromatrizz[37][399] = 9'b111111111;
assign micromatrizz[37][400] = 9'b111111111;
assign micromatrizz[37][401] = 9'b111111111;
assign micromatrizz[37][402] = 9'b111111111;
assign micromatrizz[37][403] = 9'b111111111;
assign micromatrizz[37][404] = 9'b111111111;
assign micromatrizz[37][405] = 9'b111111111;
assign micromatrizz[37][406] = 9'b111111111;
assign micromatrizz[37][407] = 9'b111111111;
assign micromatrizz[37][408] = 9'b111111111;
assign micromatrizz[37][409] = 9'b111111111;
assign micromatrizz[37][410] = 9'b111111111;
assign micromatrizz[37][411] = 9'b111111111;
assign micromatrizz[37][412] = 9'b111111111;
assign micromatrizz[37][413] = 9'b111111111;
assign micromatrizz[37][414] = 9'b111111111;
assign micromatrizz[37][415] = 9'b111111111;
assign micromatrizz[37][416] = 9'b111111111;
assign micromatrizz[37][417] = 9'b111111111;
assign micromatrizz[37][418] = 9'b111111111;
assign micromatrizz[37][419] = 9'b111111111;
assign micromatrizz[37][420] = 9'b111111111;
assign micromatrizz[37][421] = 9'b111111111;
assign micromatrizz[37][422] = 9'b111111111;
assign micromatrizz[37][423] = 9'b111111111;
assign micromatrizz[37][424] = 9'b111111111;
assign micromatrizz[37][425] = 9'b111111111;
assign micromatrizz[37][426] = 9'b111111111;
assign micromatrizz[37][427] = 9'b111111111;
assign micromatrizz[37][428] = 9'b111111111;
assign micromatrizz[37][429] = 9'b111111111;
assign micromatrizz[37][430] = 9'b111111111;
assign micromatrizz[37][431] = 9'b111111111;
assign micromatrizz[37][432] = 9'b111111111;
assign micromatrizz[37][433] = 9'b111111111;
assign micromatrizz[37][434] = 9'b111111111;
assign micromatrizz[37][435] = 9'b111111111;
assign micromatrizz[37][436] = 9'b111111111;
assign micromatrizz[37][437] = 9'b111111111;
assign micromatrizz[37][438] = 9'b111111111;
assign micromatrizz[37][439] = 9'b111111111;
assign micromatrizz[37][440] = 9'b111111111;
assign micromatrizz[37][441] = 9'b111111111;
assign micromatrizz[37][442] = 9'b111111111;
assign micromatrizz[37][443] = 9'b111111111;
assign micromatrizz[37][444] = 9'b111111111;
assign micromatrizz[37][445] = 9'b111111111;
assign micromatrizz[37][446] = 9'b111111111;
assign micromatrizz[37][447] = 9'b111111111;
assign micromatrizz[37][448] = 9'b111111111;
assign micromatrizz[37][449] = 9'b111111111;
assign micromatrizz[37][450] = 9'b111111111;
assign micromatrizz[37][451] = 9'b111111111;
assign micromatrizz[37][452] = 9'b111111111;
assign micromatrizz[37][453] = 9'b111111111;
assign micromatrizz[37][454] = 9'b111111111;
assign micromatrizz[37][455] = 9'b111111111;
assign micromatrizz[37][456] = 9'b111111111;
assign micromatrizz[37][457] = 9'b111111111;
assign micromatrizz[37][458] = 9'b111111111;
assign micromatrizz[37][459] = 9'b111111111;
assign micromatrizz[37][460] = 9'b111111111;
assign micromatrizz[37][461] = 9'b111111111;
assign micromatrizz[37][462] = 9'b111111111;
assign micromatrizz[37][463] = 9'b111111111;
assign micromatrizz[37][464] = 9'b111111111;
assign micromatrizz[37][465] = 9'b111111111;
assign micromatrizz[37][466] = 9'b111111111;
assign micromatrizz[37][467] = 9'b111111111;
assign micromatrizz[37][468] = 9'b111111111;
assign micromatrizz[37][469] = 9'b111111111;
assign micromatrizz[37][470] = 9'b111111111;
assign micromatrizz[37][471] = 9'b111111111;
assign micromatrizz[37][472] = 9'b111111111;
assign micromatrizz[37][473] = 9'b111111111;
assign micromatrizz[37][474] = 9'b111111111;
assign micromatrizz[37][475] = 9'b111111111;
assign micromatrizz[37][476] = 9'b111111111;
assign micromatrizz[37][477] = 9'b111111111;
assign micromatrizz[37][478] = 9'b111111111;
assign micromatrizz[37][479] = 9'b111111111;
assign micromatrizz[37][480] = 9'b111111111;
assign micromatrizz[37][481] = 9'b111111111;
assign micromatrizz[37][482] = 9'b111111111;
assign micromatrizz[37][483] = 9'b111111111;
assign micromatrizz[37][484] = 9'b111111111;
assign micromatrizz[37][485] = 9'b111111111;
assign micromatrizz[37][486] = 9'b111111111;
assign micromatrizz[37][487] = 9'b111111111;
assign micromatrizz[37][488] = 9'b111111111;
assign micromatrizz[37][489] = 9'b111111111;
assign micromatrizz[37][490] = 9'b111111111;
assign micromatrizz[37][491] = 9'b111111111;
assign micromatrizz[37][492] = 9'b111111111;
assign micromatrizz[37][493] = 9'b111111111;
assign micromatrizz[37][494] = 9'b111111111;
assign micromatrizz[37][495] = 9'b111111111;
assign micromatrizz[37][496] = 9'b111111111;
assign micromatrizz[37][497] = 9'b111111111;
assign micromatrizz[37][498] = 9'b111111111;
assign micromatrizz[37][499] = 9'b111111111;
assign micromatrizz[37][500] = 9'b111111111;
assign micromatrizz[37][501] = 9'b111111111;
assign micromatrizz[37][502] = 9'b111111111;
assign micromatrizz[37][503] = 9'b111111111;
assign micromatrizz[37][504] = 9'b111111111;
assign micromatrizz[37][505] = 9'b111111111;
assign micromatrizz[37][506] = 9'b111111111;
assign micromatrizz[37][507] = 9'b111111111;
assign micromatrizz[37][508] = 9'b111111111;
assign micromatrizz[37][509] = 9'b111111111;
assign micromatrizz[37][510] = 9'b111111111;
assign micromatrizz[37][511] = 9'b111111111;
assign micromatrizz[37][512] = 9'b111111111;
assign micromatrizz[37][513] = 9'b111111111;
assign micromatrizz[37][514] = 9'b111111111;
assign micromatrizz[37][515] = 9'b111111111;
assign micromatrizz[37][516] = 9'b111111111;
assign micromatrizz[37][517] = 9'b111111111;
assign micromatrizz[37][518] = 9'b111111111;
assign micromatrizz[37][519] = 9'b111111111;
assign micromatrizz[37][520] = 9'b111111111;
assign micromatrizz[37][521] = 9'b111111111;
assign micromatrizz[37][522] = 9'b111111111;
assign micromatrizz[37][523] = 9'b111111111;
assign micromatrizz[37][524] = 9'b111111111;
assign micromatrizz[37][525] = 9'b111111111;
assign micromatrizz[37][526] = 9'b111111111;
assign micromatrizz[37][527] = 9'b111111111;
assign micromatrizz[37][528] = 9'b111111111;
assign micromatrizz[37][529] = 9'b111111111;
assign micromatrizz[37][530] = 9'b111111111;
assign micromatrizz[37][531] = 9'b111111111;
assign micromatrizz[37][532] = 9'b111111111;
assign micromatrizz[37][533] = 9'b111111111;
assign micromatrizz[37][534] = 9'b111111111;
assign micromatrizz[37][535] = 9'b111111111;
assign micromatrizz[37][536] = 9'b111111111;
assign micromatrizz[37][537] = 9'b111111111;
assign micromatrizz[37][538] = 9'b111111111;
assign micromatrizz[37][539] = 9'b111111111;
assign micromatrizz[37][540] = 9'b111111111;
assign micromatrizz[37][541] = 9'b111111111;
assign micromatrizz[37][542] = 9'b111111111;
assign micromatrizz[37][543] = 9'b111111111;
assign micromatrizz[37][544] = 9'b111111111;
assign micromatrizz[37][545] = 9'b111111111;
assign micromatrizz[37][546] = 9'b111111111;
assign micromatrizz[37][547] = 9'b111111111;
assign micromatrizz[37][548] = 9'b111111111;
assign micromatrizz[37][549] = 9'b111111111;
assign micromatrizz[37][550] = 9'b111111111;
assign micromatrizz[37][551] = 9'b111111111;
assign micromatrizz[37][552] = 9'b111111111;
assign micromatrizz[37][553] = 9'b111111111;
assign micromatrizz[37][554] = 9'b111111111;
assign micromatrizz[37][555] = 9'b111111111;
assign micromatrizz[37][556] = 9'b111111111;
assign micromatrizz[37][557] = 9'b111111111;
assign micromatrizz[37][558] = 9'b111111111;
assign micromatrizz[37][559] = 9'b111111111;
assign micromatrizz[37][560] = 9'b111111111;
assign micromatrizz[37][561] = 9'b111111111;
assign micromatrizz[37][562] = 9'b111111111;
assign micromatrizz[37][563] = 9'b111111111;
assign micromatrizz[37][564] = 9'b111111111;
assign micromatrizz[37][565] = 9'b111111111;
assign micromatrizz[37][566] = 9'b111111111;
assign micromatrizz[37][567] = 9'b111111111;
assign micromatrizz[37][568] = 9'b111111111;
assign micromatrizz[37][569] = 9'b111111111;
assign micromatrizz[37][570] = 9'b111111111;
assign micromatrizz[37][571] = 9'b111111111;
assign micromatrizz[37][572] = 9'b111111111;
assign micromatrizz[37][573] = 9'b111111111;
assign micromatrizz[37][574] = 9'b111111111;
assign micromatrizz[37][575] = 9'b111111111;
assign micromatrizz[37][576] = 9'b111111111;
assign micromatrizz[37][577] = 9'b111111111;
assign micromatrizz[37][578] = 9'b111111111;
assign micromatrizz[37][579] = 9'b111111111;
assign micromatrizz[37][580] = 9'b111111111;
assign micromatrizz[37][581] = 9'b111111111;
assign micromatrizz[37][582] = 9'b111111111;
assign micromatrizz[37][583] = 9'b111111111;
assign micromatrizz[37][584] = 9'b111111111;
assign micromatrizz[37][585] = 9'b111111111;
assign micromatrizz[37][586] = 9'b111111111;
assign micromatrizz[37][587] = 9'b111111111;
assign micromatrizz[37][588] = 9'b111111111;
assign micromatrizz[37][589] = 9'b111111111;
assign micromatrizz[37][590] = 9'b111111111;
assign micromatrizz[37][591] = 9'b111111111;
assign micromatrizz[37][592] = 9'b111111111;
assign micromatrizz[37][593] = 9'b111111111;
assign micromatrizz[37][594] = 9'b111111111;
assign micromatrizz[37][595] = 9'b111111111;
assign micromatrizz[37][596] = 9'b111111111;
assign micromatrizz[37][597] = 9'b111111111;
assign micromatrizz[37][598] = 9'b111111111;
assign micromatrizz[37][599] = 9'b111111111;
assign micromatrizz[37][600] = 9'b111111111;
assign micromatrizz[37][601] = 9'b111111111;
assign micromatrizz[37][602] = 9'b111111111;
assign micromatrizz[37][603] = 9'b111111111;
assign micromatrizz[37][604] = 9'b111111111;
assign micromatrizz[37][605] = 9'b111111111;
assign micromatrizz[37][606] = 9'b111111111;
assign micromatrizz[37][607] = 9'b111111111;
assign micromatrizz[37][608] = 9'b111111111;
assign micromatrizz[37][609] = 9'b111111111;
assign micromatrizz[37][610] = 9'b111111111;
assign micromatrizz[37][611] = 9'b111111111;
assign micromatrizz[37][612] = 9'b111111111;
assign micromatrizz[37][613] = 9'b111111111;
assign micromatrizz[37][614] = 9'b111111111;
assign micromatrizz[37][615] = 9'b111111111;
assign micromatrizz[37][616] = 9'b111111111;
assign micromatrizz[37][617] = 9'b111111111;
assign micromatrizz[37][618] = 9'b111111111;
assign micromatrizz[37][619] = 9'b111111111;
assign micromatrizz[37][620] = 9'b111111111;
assign micromatrizz[37][621] = 9'b111111111;
assign micromatrizz[37][622] = 9'b111111111;
assign micromatrizz[37][623] = 9'b111111111;
assign micromatrizz[37][624] = 9'b111111111;
assign micromatrizz[37][625] = 9'b111111111;
assign micromatrizz[37][626] = 9'b111111111;
assign micromatrizz[37][627] = 9'b111111111;
assign micromatrizz[37][628] = 9'b111111111;
assign micromatrizz[37][629] = 9'b111111111;
assign micromatrizz[37][630] = 9'b111111111;
assign micromatrizz[37][631] = 9'b111111111;
assign micromatrizz[37][632] = 9'b111111111;
assign micromatrizz[37][633] = 9'b111111111;
assign micromatrizz[37][634] = 9'b111111111;
assign micromatrizz[37][635] = 9'b111111111;
assign micromatrizz[37][636] = 9'b111111111;
assign micromatrizz[37][637] = 9'b111111111;
assign micromatrizz[37][638] = 9'b111111111;
assign micromatrizz[37][639] = 9'b111111111;
assign micromatrizz[38][0] = 9'b111111111;
assign micromatrizz[38][1] = 9'b111111111;
assign micromatrizz[38][2] = 9'b111111111;
assign micromatrizz[38][3] = 9'b111111111;
assign micromatrizz[38][4] = 9'b111111111;
assign micromatrizz[38][5] = 9'b111111111;
assign micromatrizz[38][6] = 9'b111111111;
assign micromatrizz[38][7] = 9'b111111111;
assign micromatrizz[38][8] = 9'b111111111;
assign micromatrizz[38][9] = 9'b111111111;
assign micromatrizz[38][10] = 9'b111111111;
assign micromatrizz[38][11] = 9'b111111111;
assign micromatrizz[38][12] = 9'b111111111;
assign micromatrizz[38][13] = 9'b111111111;
assign micromatrizz[38][14] = 9'b111111111;
assign micromatrizz[38][15] = 9'b111111111;
assign micromatrizz[38][16] = 9'b111111111;
assign micromatrizz[38][17] = 9'b111111111;
assign micromatrizz[38][18] = 9'b111111111;
assign micromatrizz[38][19] = 9'b111111111;
assign micromatrizz[38][20] = 9'b111111111;
assign micromatrizz[38][21] = 9'b111111111;
assign micromatrizz[38][22] = 9'b111111111;
assign micromatrizz[38][23] = 9'b111111111;
assign micromatrizz[38][24] = 9'b111111111;
assign micromatrizz[38][25] = 9'b111111111;
assign micromatrizz[38][26] = 9'b111111111;
assign micromatrizz[38][27] = 9'b111111111;
assign micromatrizz[38][28] = 9'b111111111;
assign micromatrizz[38][29] = 9'b111111111;
assign micromatrizz[38][30] = 9'b111111111;
assign micromatrizz[38][31] = 9'b111111111;
assign micromatrizz[38][32] = 9'b111111111;
assign micromatrizz[38][33] = 9'b111111111;
assign micromatrizz[38][34] = 9'b111111111;
assign micromatrizz[38][35] = 9'b111111111;
assign micromatrizz[38][36] = 9'b111111111;
assign micromatrizz[38][37] = 9'b111111111;
assign micromatrizz[38][38] = 9'b111111111;
assign micromatrizz[38][39] = 9'b111111111;
assign micromatrizz[38][40] = 9'b111111111;
assign micromatrizz[38][41] = 9'b111111111;
assign micromatrizz[38][42] = 9'b111111111;
assign micromatrizz[38][43] = 9'b111111111;
assign micromatrizz[38][44] = 9'b111111111;
assign micromatrizz[38][45] = 9'b111111111;
assign micromatrizz[38][46] = 9'b111111111;
assign micromatrizz[38][47] = 9'b111111111;
assign micromatrizz[38][48] = 9'b111111111;
assign micromatrizz[38][49] = 9'b111111111;
assign micromatrizz[38][50] = 9'b111111111;
assign micromatrizz[38][51] = 9'b111111111;
assign micromatrizz[38][52] = 9'b111111111;
assign micromatrizz[38][53] = 9'b111111111;
assign micromatrizz[38][54] = 9'b111111111;
assign micromatrizz[38][55] = 9'b111111111;
assign micromatrizz[38][56] = 9'b111111111;
assign micromatrizz[38][57] = 9'b111111111;
assign micromatrizz[38][58] = 9'b111111111;
assign micromatrizz[38][59] = 9'b111111111;
assign micromatrizz[38][60] = 9'b111111111;
assign micromatrizz[38][61] = 9'b111111111;
assign micromatrizz[38][62] = 9'b111111111;
assign micromatrizz[38][63] = 9'b111111111;
assign micromatrizz[38][64] = 9'b111111111;
assign micromatrizz[38][65] = 9'b111111111;
assign micromatrizz[38][66] = 9'b111111111;
assign micromatrizz[38][67] = 9'b111111111;
assign micromatrizz[38][68] = 9'b111111111;
assign micromatrizz[38][69] = 9'b111111111;
assign micromatrizz[38][70] = 9'b111111111;
assign micromatrizz[38][71] = 9'b111111111;
assign micromatrizz[38][72] = 9'b111111111;
assign micromatrizz[38][73] = 9'b111111111;
assign micromatrizz[38][74] = 9'b111111111;
assign micromatrizz[38][75] = 9'b111111111;
assign micromatrizz[38][76] = 9'b111111111;
assign micromatrizz[38][77] = 9'b111111111;
assign micromatrizz[38][78] = 9'b111111111;
assign micromatrizz[38][79] = 9'b111111111;
assign micromatrizz[38][80] = 9'b111111111;
assign micromatrizz[38][81] = 9'b111111111;
assign micromatrizz[38][82] = 9'b111111111;
assign micromatrizz[38][83] = 9'b111111111;
assign micromatrizz[38][84] = 9'b111111111;
assign micromatrizz[38][85] = 9'b111111111;
assign micromatrizz[38][86] = 9'b111111111;
assign micromatrizz[38][87] = 9'b111111111;
assign micromatrizz[38][88] = 9'b111111111;
assign micromatrizz[38][89] = 9'b111111111;
assign micromatrizz[38][90] = 9'b111111111;
assign micromatrizz[38][91] = 9'b111111111;
assign micromatrizz[38][92] = 9'b111111111;
assign micromatrizz[38][93] = 9'b111111111;
assign micromatrizz[38][94] = 9'b111111111;
assign micromatrizz[38][95] = 9'b111111111;
assign micromatrizz[38][96] = 9'b111111111;
assign micromatrizz[38][97] = 9'b111111111;
assign micromatrizz[38][98] = 9'b111111111;
assign micromatrizz[38][99] = 9'b111111111;
assign micromatrizz[38][100] = 9'b111111111;
assign micromatrizz[38][101] = 9'b111111111;
assign micromatrizz[38][102] = 9'b111111111;
assign micromatrizz[38][103] = 9'b111111111;
assign micromatrizz[38][104] = 9'b111111111;
assign micromatrizz[38][105] = 9'b111111111;
assign micromatrizz[38][106] = 9'b111111111;
assign micromatrizz[38][107] = 9'b111111111;
assign micromatrizz[38][108] = 9'b111111111;
assign micromatrizz[38][109] = 9'b111111111;
assign micromatrizz[38][110] = 9'b111111111;
assign micromatrizz[38][111] = 9'b111111111;
assign micromatrizz[38][112] = 9'b111111111;
assign micromatrizz[38][113] = 9'b111111111;
assign micromatrizz[38][114] = 9'b111111111;
assign micromatrizz[38][115] = 9'b111111111;
assign micromatrizz[38][116] = 9'b111111111;
assign micromatrizz[38][117] = 9'b111111111;
assign micromatrizz[38][118] = 9'b111111111;
assign micromatrizz[38][119] = 9'b111111111;
assign micromatrizz[38][120] = 9'b111111111;
assign micromatrizz[38][121] = 9'b111111111;
assign micromatrizz[38][122] = 9'b111111111;
assign micromatrizz[38][123] = 9'b111111111;
assign micromatrizz[38][124] = 9'b111111111;
assign micromatrizz[38][125] = 9'b111111111;
assign micromatrizz[38][126] = 9'b111111111;
assign micromatrizz[38][127] = 9'b111111111;
assign micromatrizz[38][128] = 9'b111111111;
assign micromatrizz[38][129] = 9'b111111111;
assign micromatrizz[38][130] = 9'b111111111;
assign micromatrizz[38][131] = 9'b111111111;
assign micromatrizz[38][132] = 9'b111111111;
assign micromatrizz[38][133] = 9'b111111111;
assign micromatrizz[38][134] = 9'b111111111;
assign micromatrizz[38][135] = 9'b111111111;
assign micromatrizz[38][136] = 9'b111111111;
assign micromatrizz[38][137] = 9'b111111111;
assign micromatrizz[38][138] = 9'b111111111;
assign micromatrizz[38][139] = 9'b111111111;
assign micromatrizz[38][140] = 9'b111111111;
assign micromatrizz[38][141] = 9'b111111111;
assign micromatrizz[38][142] = 9'b111111111;
assign micromatrizz[38][143] = 9'b111111111;
assign micromatrizz[38][144] = 9'b111111111;
assign micromatrizz[38][145] = 9'b111111111;
assign micromatrizz[38][146] = 9'b111111111;
assign micromatrizz[38][147] = 9'b111111111;
assign micromatrizz[38][148] = 9'b111111111;
assign micromatrizz[38][149] = 9'b111111111;
assign micromatrizz[38][150] = 9'b111111111;
assign micromatrizz[38][151] = 9'b111111111;
assign micromatrizz[38][152] = 9'b111111111;
assign micromatrizz[38][153] = 9'b111111111;
assign micromatrizz[38][154] = 9'b111111111;
assign micromatrizz[38][155] = 9'b111111111;
assign micromatrizz[38][156] = 9'b111111111;
assign micromatrizz[38][157] = 9'b111111111;
assign micromatrizz[38][158] = 9'b111111111;
assign micromatrizz[38][159] = 9'b111111111;
assign micromatrizz[38][160] = 9'b111111111;
assign micromatrizz[38][161] = 9'b111111111;
assign micromatrizz[38][162] = 9'b111111111;
assign micromatrizz[38][163] = 9'b111111111;
assign micromatrizz[38][164] = 9'b111111111;
assign micromatrizz[38][165] = 9'b111111111;
assign micromatrizz[38][166] = 9'b111111111;
assign micromatrizz[38][167] = 9'b111111111;
assign micromatrizz[38][168] = 9'b111111111;
assign micromatrizz[38][169] = 9'b111111111;
assign micromatrizz[38][170] = 9'b111111111;
assign micromatrizz[38][171] = 9'b111111111;
assign micromatrizz[38][172] = 9'b111111111;
assign micromatrizz[38][173] = 9'b111111111;
assign micromatrizz[38][174] = 9'b111111111;
assign micromatrizz[38][175] = 9'b111111111;
assign micromatrizz[38][176] = 9'b111111111;
assign micromatrizz[38][177] = 9'b111111111;
assign micromatrizz[38][178] = 9'b111111111;
assign micromatrizz[38][179] = 9'b111111111;
assign micromatrizz[38][180] = 9'b111111111;
assign micromatrizz[38][181] = 9'b111111111;
assign micromatrizz[38][182] = 9'b111111111;
assign micromatrizz[38][183] = 9'b111111111;
assign micromatrizz[38][184] = 9'b111111111;
assign micromatrizz[38][185] = 9'b111111111;
assign micromatrizz[38][186] = 9'b111111111;
assign micromatrizz[38][187] = 9'b111111111;
assign micromatrizz[38][188] = 9'b111111111;
assign micromatrizz[38][189] = 9'b111111111;
assign micromatrizz[38][190] = 9'b111111111;
assign micromatrizz[38][191] = 9'b111111111;
assign micromatrizz[38][192] = 9'b111111111;
assign micromatrizz[38][193] = 9'b111111111;
assign micromatrizz[38][194] = 9'b111111111;
assign micromatrizz[38][195] = 9'b111111111;
assign micromatrizz[38][196] = 9'b111111111;
assign micromatrizz[38][197] = 9'b111111111;
assign micromatrizz[38][198] = 9'b111111111;
assign micromatrizz[38][199] = 9'b111111111;
assign micromatrizz[38][200] = 9'b111111111;
assign micromatrizz[38][201] = 9'b111111111;
assign micromatrizz[38][202] = 9'b111111111;
assign micromatrizz[38][203] = 9'b111111111;
assign micromatrizz[38][204] = 9'b111111111;
assign micromatrizz[38][205] = 9'b111111111;
assign micromatrizz[38][206] = 9'b111111111;
assign micromatrizz[38][207] = 9'b111111111;
assign micromatrizz[38][208] = 9'b111111111;
assign micromatrizz[38][209] = 9'b111111111;
assign micromatrizz[38][210] = 9'b111111111;
assign micromatrizz[38][211] = 9'b111111111;
assign micromatrizz[38][212] = 9'b111111111;
assign micromatrizz[38][213] = 9'b111111111;
assign micromatrizz[38][214] = 9'b111111111;
assign micromatrizz[38][215] = 9'b111111111;
assign micromatrizz[38][216] = 9'b111111111;
assign micromatrizz[38][217] = 9'b111111111;
assign micromatrizz[38][218] = 9'b111111111;
assign micromatrizz[38][219] = 9'b111111111;
assign micromatrizz[38][220] = 9'b111111111;
assign micromatrizz[38][221] = 9'b111111111;
assign micromatrizz[38][222] = 9'b111111111;
assign micromatrizz[38][223] = 9'b111111111;
assign micromatrizz[38][224] = 9'b111111111;
assign micromatrizz[38][225] = 9'b111111111;
assign micromatrizz[38][226] = 9'b111111111;
assign micromatrizz[38][227] = 9'b111111111;
assign micromatrizz[38][228] = 9'b111111111;
assign micromatrizz[38][229] = 9'b111111111;
assign micromatrizz[38][230] = 9'b111111111;
assign micromatrizz[38][231] = 9'b111111111;
assign micromatrizz[38][232] = 9'b111111111;
assign micromatrizz[38][233] = 9'b111111111;
assign micromatrizz[38][234] = 9'b111111111;
assign micromatrizz[38][235] = 9'b111111111;
assign micromatrizz[38][236] = 9'b111111111;
assign micromatrizz[38][237] = 9'b111111111;
assign micromatrizz[38][238] = 9'b111111111;
assign micromatrizz[38][239] = 9'b111111111;
assign micromatrizz[38][240] = 9'b111111111;
assign micromatrizz[38][241] = 9'b111111111;
assign micromatrizz[38][242] = 9'b111111111;
assign micromatrizz[38][243] = 9'b111111111;
assign micromatrizz[38][244] = 9'b111111111;
assign micromatrizz[38][245] = 9'b111111111;
assign micromatrizz[38][246] = 9'b111111111;
assign micromatrizz[38][247] = 9'b111111111;
assign micromatrizz[38][248] = 9'b111111111;
assign micromatrizz[38][249] = 9'b111111111;
assign micromatrizz[38][250] = 9'b111111111;
assign micromatrizz[38][251] = 9'b111111111;
assign micromatrizz[38][252] = 9'b111111111;
assign micromatrizz[38][253] = 9'b111111111;
assign micromatrizz[38][254] = 9'b111111111;
assign micromatrizz[38][255] = 9'b111111111;
assign micromatrizz[38][256] = 9'b111111111;
assign micromatrizz[38][257] = 9'b111111111;
assign micromatrizz[38][258] = 9'b111111111;
assign micromatrizz[38][259] = 9'b111111111;
assign micromatrizz[38][260] = 9'b111111111;
assign micromatrizz[38][261] = 9'b111111111;
assign micromatrizz[38][262] = 9'b111111111;
assign micromatrizz[38][263] = 9'b111111111;
assign micromatrizz[38][264] = 9'b111111111;
assign micromatrizz[38][265] = 9'b111111111;
assign micromatrizz[38][266] = 9'b111111111;
assign micromatrizz[38][267] = 9'b111111111;
assign micromatrizz[38][268] = 9'b111111111;
assign micromatrizz[38][269] = 9'b111111111;
assign micromatrizz[38][270] = 9'b111111111;
assign micromatrizz[38][271] = 9'b111111111;
assign micromatrizz[38][272] = 9'b111111111;
assign micromatrizz[38][273] = 9'b111111111;
assign micromatrizz[38][274] = 9'b111111111;
assign micromatrizz[38][275] = 9'b111111111;
assign micromatrizz[38][276] = 9'b111111111;
assign micromatrizz[38][277] = 9'b111111111;
assign micromatrizz[38][278] = 9'b111111111;
assign micromatrizz[38][279] = 9'b111111111;
assign micromatrizz[38][280] = 9'b111111111;
assign micromatrizz[38][281] = 9'b111111111;
assign micromatrizz[38][282] = 9'b111111111;
assign micromatrizz[38][283] = 9'b111111111;
assign micromatrizz[38][284] = 9'b111111111;
assign micromatrizz[38][285] = 9'b111111111;
assign micromatrizz[38][286] = 9'b111111111;
assign micromatrizz[38][287] = 9'b111111111;
assign micromatrizz[38][288] = 9'b111111111;
assign micromatrizz[38][289] = 9'b111111111;
assign micromatrizz[38][290] = 9'b111111111;
assign micromatrizz[38][291] = 9'b111111111;
assign micromatrizz[38][292] = 9'b111111111;
assign micromatrizz[38][293] = 9'b111111111;
assign micromatrizz[38][294] = 9'b111111111;
assign micromatrizz[38][295] = 9'b111111111;
assign micromatrizz[38][296] = 9'b111111111;
assign micromatrizz[38][297] = 9'b111111111;
assign micromatrizz[38][298] = 9'b111111111;
assign micromatrizz[38][299] = 9'b111111111;
assign micromatrizz[38][300] = 9'b111111111;
assign micromatrizz[38][301] = 9'b111111111;
assign micromatrizz[38][302] = 9'b111111111;
assign micromatrizz[38][303] = 9'b111111111;
assign micromatrizz[38][304] = 9'b111111111;
assign micromatrizz[38][305] = 9'b111111111;
assign micromatrizz[38][306] = 9'b111111111;
assign micromatrizz[38][307] = 9'b111111111;
assign micromatrizz[38][308] = 9'b111111111;
assign micromatrizz[38][309] = 9'b111111111;
assign micromatrizz[38][310] = 9'b111111111;
assign micromatrizz[38][311] = 9'b111111111;
assign micromatrizz[38][312] = 9'b111111111;
assign micromatrizz[38][313] = 9'b111111111;
assign micromatrizz[38][314] = 9'b111111111;
assign micromatrizz[38][315] = 9'b111111111;
assign micromatrizz[38][316] = 9'b111111111;
assign micromatrizz[38][317] = 9'b111111111;
assign micromatrizz[38][318] = 9'b111111111;
assign micromatrizz[38][319] = 9'b111111111;
assign micromatrizz[38][320] = 9'b111111111;
assign micromatrizz[38][321] = 9'b111111111;
assign micromatrizz[38][322] = 9'b111111111;
assign micromatrizz[38][323] = 9'b111111111;
assign micromatrizz[38][324] = 9'b111111111;
assign micromatrizz[38][325] = 9'b111111111;
assign micromatrizz[38][326] = 9'b111111111;
assign micromatrizz[38][327] = 9'b111111111;
assign micromatrizz[38][328] = 9'b111111111;
assign micromatrizz[38][329] = 9'b111111111;
assign micromatrizz[38][330] = 9'b111111111;
assign micromatrizz[38][331] = 9'b111111111;
assign micromatrizz[38][332] = 9'b111111111;
assign micromatrizz[38][333] = 9'b111111111;
assign micromatrizz[38][334] = 9'b111111111;
assign micromatrizz[38][335] = 9'b111111111;
assign micromatrizz[38][336] = 9'b111111111;
assign micromatrizz[38][337] = 9'b111111111;
assign micromatrizz[38][338] = 9'b111111111;
assign micromatrizz[38][339] = 9'b111111111;
assign micromatrizz[38][340] = 9'b111111111;
assign micromatrizz[38][341] = 9'b111111111;
assign micromatrizz[38][342] = 9'b111111111;
assign micromatrizz[38][343] = 9'b111111111;
assign micromatrizz[38][344] = 9'b111111111;
assign micromatrizz[38][345] = 9'b111111111;
assign micromatrizz[38][346] = 9'b111111111;
assign micromatrizz[38][347] = 9'b111111111;
assign micromatrizz[38][348] = 9'b111111111;
assign micromatrizz[38][349] = 9'b111111111;
assign micromatrizz[38][350] = 9'b111111111;
assign micromatrizz[38][351] = 9'b111111111;
assign micromatrizz[38][352] = 9'b111111111;
assign micromatrizz[38][353] = 9'b111111111;
assign micromatrizz[38][354] = 9'b111111111;
assign micromatrizz[38][355] = 9'b111111111;
assign micromatrizz[38][356] = 9'b111111111;
assign micromatrizz[38][357] = 9'b111111111;
assign micromatrizz[38][358] = 9'b111111111;
assign micromatrizz[38][359] = 9'b111111111;
assign micromatrizz[38][360] = 9'b111111111;
assign micromatrizz[38][361] = 9'b111111111;
assign micromatrizz[38][362] = 9'b111111111;
assign micromatrizz[38][363] = 9'b111111111;
assign micromatrizz[38][364] = 9'b111111111;
assign micromatrizz[38][365] = 9'b111111111;
assign micromatrizz[38][366] = 9'b111111111;
assign micromatrizz[38][367] = 9'b111111111;
assign micromatrizz[38][368] = 9'b111111111;
assign micromatrizz[38][369] = 9'b111111111;
assign micromatrizz[38][370] = 9'b111111111;
assign micromatrizz[38][371] = 9'b111111111;
assign micromatrizz[38][372] = 9'b111111111;
assign micromatrizz[38][373] = 9'b111111111;
assign micromatrizz[38][374] = 9'b111111111;
assign micromatrizz[38][375] = 9'b111111111;
assign micromatrizz[38][376] = 9'b111111111;
assign micromatrizz[38][377] = 9'b111111111;
assign micromatrizz[38][378] = 9'b111111111;
assign micromatrizz[38][379] = 9'b111111111;
assign micromatrizz[38][380] = 9'b111111111;
assign micromatrizz[38][381] = 9'b111111111;
assign micromatrizz[38][382] = 9'b111111111;
assign micromatrizz[38][383] = 9'b111111111;
assign micromatrizz[38][384] = 9'b111111111;
assign micromatrizz[38][385] = 9'b111111111;
assign micromatrizz[38][386] = 9'b111111111;
assign micromatrizz[38][387] = 9'b111111111;
assign micromatrizz[38][388] = 9'b111111111;
assign micromatrizz[38][389] = 9'b111111111;
assign micromatrizz[38][390] = 9'b111111111;
assign micromatrizz[38][391] = 9'b111111111;
assign micromatrizz[38][392] = 9'b111111111;
assign micromatrizz[38][393] = 9'b111111111;
assign micromatrizz[38][394] = 9'b111111111;
assign micromatrizz[38][395] = 9'b111111111;
assign micromatrizz[38][396] = 9'b111111111;
assign micromatrizz[38][397] = 9'b111111111;
assign micromatrizz[38][398] = 9'b111111111;
assign micromatrizz[38][399] = 9'b111111111;
assign micromatrizz[38][400] = 9'b111111111;
assign micromatrizz[38][401] = 9'b111111111;
assign micromatrizz[38][402] = 9'b111111111;
assign micromatrizz[38][403] = 9'b111111111;
assign micromatrizz[38][404] = 9'b111111111;
assign micromatrizz[38][405] = 9'b111111111;
assign micromatrizz[38][406] = 9'b111111111;
assign micromatrizz[38][407] = 9'b111111111;
assign micromatrizz[38][408] = 9'b111111111;
assign micromatrizz[38][409] = 9'b111111111;
assign micromatrizz[38][410] = 9'b111111111;
assign micromatrizz[38][411] = 9'b111111111;
assign micromatrizz[38][412] = 9'b111111111;
assign micromatrizz[38][413] = 9'b111111111;
assign micromatrizz[38][414] = 9'b111111111;
assign micromatrizz[38][415] = 9'b111111111;
assign micromatrizz[38][416] = 9'b111111111;
assign micromatrizz[38][417] = 9'b111111111;
assign micromatrizz[38][418] = 9'b111111111;
assign micromatrizz[38][419] = 9'b111111111;
assign micromatrizz[38][420] = 9'b111111111;
assign micromatrizz[38][421] = 9'b111111111;
assign micromatrizz[38][422] = 9'b111111111;
assign micromatrizz[38][423] = 9'b111111111;
assign micromatrizz[38][424] = 9'b111111111;
assign micromatrizz[38][425] = 9'b111111111;
assign micromatrizz[38][426] = 9'b111111111;
assign micromatrizz[38][427] = 9'b111111111;
assign micromatrizz[38][428] = 9'b111111111;
assign micromatrizz[38][429] = 9'b111111111;
assign micromatrizz[38][430] = 9'b111111111;
assign micromatrizz[38][431] = 9'b111111111;
assign micromatrizz[38][432] = 9'b111111111;
assign micromatrizz[38][433] = 9'b111111111;
assign micromatrizz[38][434] = 9'b111111111;
assign micromatrizz[38][435] = 9'b111111111;
assign micromatrizz[38][436] = 9'b111111111;
assign micromatrizz[38][437] = 9'b111111111;
assign micromatrizz[38][438] = 9'b111111111;
assign micromatrizz[38][439] = 9'b111111111;
assign micromatrizz[38][440] = 9'b111111111;
assign micromatrizz[38][441] = 9'b111111111;
assign micromatrizz[38][442] = 9'b111111111;
assign micromatrizz[38][443] = 9'b111111111;
assign micromatrizz[38][444] = 9'b111111111;
assign micromatrizz[38][445] = 9'b111111111;
assign micromatrizz[38][446] = 9'b111111111;
assign micromatrizz[38][447] = 9'b111111111;
assign micromatrizz[38][448] = 9'b111111111;
assign micromatrizz[38][449] = 9'b111111111;
assign micromatrizz[38][450] = 9'b111111111;
assign micromatrizz[38][451] = 9'b111111111;
assign micromatrizz[38][452] = 9'b111111111;
assign micromatrizz[38][453] = 9'b111111111;
assign micromatrizz[38][454] = 9'b111111111;
assign micromatrizz[38][455] = 9'b111111111;
assign micromatrizz[38][456] = 9'b111111111;
assign micromatrizz[38][457] = 9'b111111111;
assign micromatrizz[38][458] = 9'b111111111;
assign micromatrizz[38][459] = 9'b111111111;
assign micromatrizz[38][460] = 9'b111111111;
assign micromatrizz[38][461] = 9'b111111111;
assign micromatrizz[38][462] = 9'b111111111;
assign micromatrizz[38][463] = 9'b111111111;
assign micromatrizz[38][464] = 9'b111111111;
assign micromatrizz[38][465] = 9'b111111111;
assign micromatrizz[38][466] = 9'b111111111;
assign micromatrizz[38][467] = 9'b111111111;
assign micromatrizz[38][468] = 9'b111111111;
assign micromatrizz[38][469] = 9'b111111111;
assign micromatrizz[38][470] = 9'b111111111;
assign micromatrizz[38][471] = 9'b111111111;
assign micromatrizz[38][472] = 9'b111111111;
assign micromatrizz[38][473] = 9'b111111111;
assign micromatrizz[38][474] = 9'b111111111;
assign micromatrizz[38][475] = 9'b111111111;
assign micromatrizz[38][476] = 9'b111111111;
assign micromatrizz[38][477] = 9'b111111111;
assign micromatrizz[38][478] = 9'b111111111;
assign micromatrizz[38][479] = 9'b111111111;
assign micromatrizz[38][480] = 9'b111111111;
assign micromatrizz[38][481] = 9'b111111111;
assign micromatrizz[38][482] = 9'b111111111;
assign micromatrizz[38][483] = 9'b111111111;
assign micromatrizz[38][484] = 9'b111111111;
assign micromatrizz[38][485] = 9'b111111111;
assign micromatrizz[38][486] = 9'b111111111;
assign micromatrizz[38][487] = 9'b111111111;
assign micromatrizz[38][488] = 9'b111111111;
assign micromatrizz[38][489] = 9'b111111111;
assign micromatrizz[38][490] = 9'b111111111;
assign micromatrizz[38][491] = 9'b111111111;
assign micromatrizz[38][492] = 9'b111111111;
assign micromatrizz[38][493] = 9'b111111111;
assign micromatrizz[38][494] = 9'b111111111;
assign micromatrizz[38][495] = 9'b111111111;
assign micromatrizz[38][496] = 9'b111111111;
assign micromatrizz[38][497] = 9'b111111111;
assign micromatrizz[38][498] = 9'b111111111;
assign micromatrizz[38][499] = 9'b111111111;
assign micromatrizz[38][500] = 9'b111111111;
assign micromatrizz[38][501] = 9'b111111111;
assign micromatrizz[38][502] = 9'b111111111;
assign micromatrizz[38][503] = 9'b111111111;
assign micromatrizz[38][504] = 9'b111111111;
assign micromatrizz[38][505] = 9'b111111111;
assign micromatrizz[38][506] = 9'b111111111;
assign micromatrizz[38][507] = 9'b111111111;
assign micromatrizz[38][508] = 9'b111111111;
assign micromatrizz[38][509] = 9'b111111111;
assign micromatrizz[38][510] = 9'b111111111;
assign micromatrizz[38][511] = 9'b111111111;
assign micromatrizz[38][512] = 9'b111111111;
assign micromatrizz[38][513] = 9'b111111111;
assign micromatrizz[38][514] = 9'b111111111;
assign micromatrizz[38][515] = 9'b111111111;
assign micromatrizz[38][516] = 9'b111111111;
assign micromatrizz[38][517] = 9'b111111111;
assign micromatrizz[38][518] = 9'b111111111;
assign micromatrizz[38][519] = 9'b111111111;
assign micromatrizz[38][520] = 9'b111111111;
assign micromatrizz[38][521] = 9'b111111111;
assign micromatrizz[38][522] = 9'b111111111;
assign micromatrizz[38][523] = 9'b111111111;
assign micromatrizz[38][524] = 9'b111111111;
assign micromatrizz[38][525] = 9'b111111111;
assign micromatrizz[38][526] = 9'b111111111;
assign micromatrizz[38][527] = 9'b111111111;
assign micromatrizz[38][528] = 9'b111111111;
assign micromatrizz[38][529] = 9'b111111111;
assign micromatrizz[38][530] = 9'b111111111;
assign micromatrizz[38][531] = 9'b111111111;
assign micromatrizz[38][532] = 9'b111111111;
assign micromatrizz[38][533] = 9'b111111111;
assign micromatrizz[38][534] = 9'b111111111;
assign micromatrizz[38][535] = 9'b111111111;
assign micromatrizz[38][536] = 9'b111111111;
assign micromatrizz[38][537] = 9'b111111111;
assign micromatrizz[38][538] = 9'b111111111;
assign micromatrizz[38][539] = 9'b111111111;
assign micromatrizz[38][540] = 9'b111111111;
assign micromatrizz[38][541] = 9'b111111111;
assign micromatrizz[38][542] = 9'b111111111;
assign micromatrizz[38][543] = 9'b111111111;
assign micromatrizz[38][544] = 9'b111111111;
assign micromatrizz[38][545] = 9'b111111111;
assign micromatrizz[38][546] = 9'b111111111;
assign micromatrizz[38][547] = 9'b111111111;
assign micromatrizz[38][548] = 9'b111111111;
assign micromatrizz[38][549] = 9'b111111111;
assign micromatrizz[38][550] = 9'b111111111;
assign micromatrizz[38][551] = 9'b111111111;
assign micromatrizz[38][552] = 9'b111111111;
assign micromatrizz[38][553] = 9'b111111111;
assign micromatrizz[38][554] = 9'b111111111;
assign micromatrizz[38][555] = 9'b111111111;
assign micromatrizz[38][556] = 9'b111111111;
assign micromatrizz[38][557] = 9'b111111111;
assign micromatrizz[38][558] = 9'b111111111;
assign micromatrizz[38][559] = 9'b111111111;
assign micromatrizz[38][560] = 9'b111111111;
assign micromatrizz[38][561] = 9'b111111111;
assign micromatrizz[38][562] = 9'b111111111;
assign micromatrizz[38][563] = 9'b111111111;
assign micromatrizz[38][564] = 9'b111111111;
assign micromatrizz[38][565] = 9'b111111111;
assign micromatrizz[38][566] = 9'b111111111;
assign micromatrizz[38][567] = 9'b111111111;
assign micromatrizz[38][568] = 9'b111111111;
assign micromatrizz[38][569] = 9'b111111111;
assign micromatrizz[38][570] = 9'b111111111;
assign micromatrizz[38][571] = 9'b111111111;
assign micromatrizz[38][572] = 9'b111111111;
assign micromatrizz[38][573] = 9'b111111111;
assign micromatrizz[38][574] = 9'b111111111;
assign micromatrizz[38][575] = 9'b111111111;
assign micromatrizz[38][576] = 9'b111111111;
assign micromatrizz[38][577] = 9'b111111111;
assign micromatrizz[38][578] = 9'b111111111;
assign micromatrizz[38][579] = 9'b111111111;
assign micromatrizz[38][580] = 9'b111111111;
assign micromatrizz[38][581] = 9'b111111111;
assign micromatrizz[38][582] = 9'b111111111;
assign micromatrizz[38][583] = 9'b111111111;
assign micromatrizz[38][584] = 9'b111111111;
assign micromatrizz[38][585] = 9'b111111111;
assign micromatrizz[38][586] = 9'b111111111;
assign micromatrizz[38][587] = 9'b111111111;
assign micromatrizz[38][588] = 9'b111111111;
assign micromatrizz[38][589] = 9'b111111111;
assign micromatrizz[38][590] = 9'b111111111;
assign micromatrizz[38][591] = 9'b111111111;
assign micromatrizz[38][592] = 9'b111111111;
assign micromatrizz[38][593] = 9'b111111111;
assign micromatrizz[38][594] = 9'b111111111;
assign micromatrizz[38][595] = 9'b111111111;
assign micromatrizz[38][596] = 9'b111111111;
assign micromatrizz[38][597] = 9'b111111111;
assign micromatrizz[38][598] = 9'b111111111;
assign micromatrizz[38][599] = 9'b111111111;
assign micromatrizz[38][600] = 9'b111111111;
assign micromatrizz[38][601] = 9'b111111111;
assign micromatrizz[38][602] = 9'b111111111;
assign micromatrizz[38][603] = 9'b111111111;
assign micromatrizz[38][604] = 9'b111111111;
assign micromatrizz[38][605] = 9'b111111111;
assign micromatrizz[38][606] = 9'b111111111;
assign micromatrizz[38][607] = 9'b111111111;
assign micromatrizz[38][608] = 9'b111111111;
assign micromatrizz[38][609] = 9'b111111111;
assign micromatrizz[38][610] = 9'b111111111;
assign micromatrizz[38][611] = 9'b111111111;
assign micromatrizz[38][612] = 9'b111111111;
assign micromatrizz[38][613] = 9'b111111111;
assign micromatrizz[38][614] = 9'b111111111;
assign micromatrizz[38][615] = 9'b111111111;
assign micromatrizz[38][616] = 9'b111111111;
assign micromatrizz[38][617] = 9'b111111111;
assign micromatrizz[38][618] = 9'b111111111;
assign micromatrizz[38][619] = 9'b111111111;
assign micromatrizz[38][620] = 9'b111111111;
assign micromatrizz[38][621] = 9'b111111111;
assign micromatrizz[38][622] = 9'b111111111;
assign micromatrizz[38][623] = 9'b111111111;
assign micromatrizz[38][624] = 9'b111111111;
assign micromatrizz[38][625] = 9'b111111111;
assign micromatrizz[38][626] = 9'b111111111;
assign micromatrizz[38][627] = 9'b111111111;
assign micromatrizz[38][628] = 9'b111111111;
assign micromatrizz[38][629] = 9'b111111111;
assign micromatrizz[38][630] = 9'b111111111;
assign micromatrizz[38][631] = 9'b111111111;
assign micromatrizz[38][632] = 9'b111111111;
assign micromatrizz[38][633] = 9'b111111111;
assign micromatrizz[38][634] = 9'b111111111;
assign micromatrizz[38][635] = 9'b111111111;
assign micromatrizz[38][636] = 9'b111111111;
assign micromatrizz[38][637] = 9'b111111111;
assign micromatrizz[38][638] = 9'b111111111;
assign micromatrizz[38][639] = 9'b111111111;
assign micromatrizz[39][0] = 9'b111111111;
assign micromatrizz[39][1] = 9'b111111111;
assign micromatrizz[39][2] = 9'b111111111;
assign micromatrizz[39][3] = 9'b111111111;
assign micromatrizz[39][4] = 9'b111111111;
assign micromatrizz[39][5] = 9'b111111111;
assign micromatrizz[39][6] = 9'b111111111;
assign micromatrizz[39][7] = 9'b111111111;
assign micromatrizz[39][8] = 9'b111111111;
assign micromatrizz[39][9] = 9'b111111111;
assign micromatrizz[39][10] = 9'b111111111;
assign micromatrizz[39][11] = 9'b111111111;
assign micromatrizz[39][12] = 9'b111111111;
assign micromatrizz[39][13] = 9'b111111111;
assign micromatrizz[39][14] = 9'b111111111;
assign micromatrizz[39][15] = 9'b111111111;
assign micromatrizz[39][16] = 9'b111111111;
assign micromatrizz[39][17] = 9'b111111111;
assign micromatrizz[39][18] = 9'b111111111;
assign micromatrizz[39][19] = 9'b111111111;
assign micromatrizz[39][20] = 9'b111111111;
assign micromatrizz[39][21] = 9'b111111111;
assign micromatrizz[39][22] = 9'b111111111;
assign micromatrizz[39][23] = 9'b111111111;
assign micromatrizz[39][24] = 9'b111111111;
assign micromatrizz[39][25] = 9'b111111111;
assign micromatrizz[39][26] = 9'b111111111;
assign micromatrizz[39][27] = 9'b111111111;
assign micromatrizz[39][28] = 9'b111111111;
assign micromatrizz[39][29] = 9'b111111111;
assign micromatrizz[39][30] = 9'b111111111;
assign micromatrizz[39][31] = 9'b111111111;
assign micromatrizz[39][32] = 9'b111111111;
assign micromatrizz[39][33] = 9'b111111111;
assign micromatrizz[39][34] = 9'b111111111;
assign micromatrizz[39][35] = 9'b111111111;
assign micromatrizz[39][36] = 9'b111111111;
assign micromatrizz[39][37] = 9'b111111111;
assign micromatrizz[39][38] = 9'b111111111;
assign micromatrizz[39][39] = 9'b111111111;
assign micromatrizz[39][40] = 9'b111111111;
assign micromatrizz[39][41] = 9'b111111111;
assign micromatrizz[39][42] = 9'b111111111;
assign micromatrizz[39][43] = 9'b111111111;
assign micromatrizz[39][44] = 9'b111111111;
assign micromatrizz[39][45] = 9'b111111111;
assign micromatrizz[39][46] = 9'b111111111;
assign micromatrizz[39][47] = 9'b111111111;
assign micromatrizz[39][48] = 9'b111111111;
assign micromatrizz[39][49] = 9'b111111111;
assign micromatrizz[39][50] = 9'b111111111;
assign micromatrizz[39][51] = 9'b111111111;
assign micromatrizz[39][52] = 9'b111111111;
assign micromatrizz[39][53] = 9'b111111111;
assign micromatrizz[39][54] = 9'b111111111;
assign micromatrizz[39][55] = 9'b111111111;
assign micromatrizz[39][56] = 9'b111111111;
assign micromatrizz[39][57] = 9'b111111111;
assign micromatrizz[39][58] = 9'b111111111;
assign micromatrizz[39][59] = 9'b111111111;
assign micromatrizz[39][60] = 9'b111111111;
assign micromatrizz[39][61] = 9'b111111111;
assign micromatrizz[39][62] = 9'b111111111;
assign micromatrizz[39][63] = 9'b111111111;
assign micromatrizz[39][64] = 9'b111111111;
assign micromatrizz[39][65] = 9'b111111111;
assign micromatrizz[39][66] = 9'b111111111;
assign micromatrizz[39][67] = 9'b111111111;
assign micromatrizz[39][68] = 9'b111111111;
assign micromatrizz[39][69] = 9'b111111111;
assign micromatrizz[39][70] = 9'b111111111;
assign micromatrizz[39][71] = 9'b111111111;
assign micromatrizz[39][72] = 9'b111111111;
assign micromatrizz[39][73] = 9'b111111111;
assign micromatrizz[39][74] = 9'b111111111;
assign micromatrizz[39][75] = 9'b111111111;
assign micromatrizz[39][76] = 9'b111111111;
assign micromatrizz[39][77] = 9'b111111111;
assign micromatrizz[39][78] = 9'b111111111;
assign micromatrizz[39][79] = 9'b111111111;
assign micromatrizz[39][80] = 9'b111111111;
assign micromatrizz[39][81] = 9'b111111111;
assign micromatrizz[39][82] = 9'b111111111;
assign micromatrizz[39][83] = 9'b111111111;
assign micromatrizz[39][84] = 9'b111111111;
assign micromatrizz[39][85] = 9'b111111111;
assign micromatrizz[39][86] = 9'b111111111;
assign micromatrizz[39][87] = 9'b111111111;
assign micromatrizz[39][88] = 9'b111111111;
assign micromatrizz[39][89] = 9'b111111111;
assign micromatrizz[39][90] = 9'b111111111;
assign micromatrizz[39][91] = 9'b111111111;
assign micromatrizz[39][92] = 9'b111111111;
assign micromatrizz[39][93] = 9'b111111111;
assign micromatrizz[39][94] = 9'b111111111;
assign micromatrizz[39][95] = 9'b111111111;
assign micromatrizz[39][96] = 9'b111111111;
assign micromatrizz[39][97] = 9'b111111111;
assign micromatrizz[39][98] = 9'b111111111;
assign micromatrizz[39][99] = 9'b111111111;
assign micromatrizz[39][100] = 9'b111111111;
assign micromatrizz[39][101] = 9'b111111111;
assign micromatrizz[39][102] = 9'b111111111;
assign micromatrizz[39][103] = 9'b111111111;
assign micromatrizz[39][104] = 9'b111111111;
assign micromatrizz[39][105] = 9'b111111111;
assign micromatrizz[39][106] = 9'b111111111;
assign micromatrizz[39][107] = 9'b111111111;
assign micromatrizz[39][108] = 9'b111111111;
assign micromatrizz[39][109] = 9'b111111111;
assign micromatrizz[39][110] = 9'b111111111;
assign micromatrizz[39][111] = 9'b111111111;
assign micromatrizz[39][112] = 9'b111111111;
assign micromatrizz[39][113] = 9'b111111111;
assign micromatrizz[39][114] = 9'b111111111;
assign micromatrizz[39][115] = 9'b111111111;
assign micromatrizz[39][116] = 9'b111111111;
assign micromatrizz[39][117] = 9'b111111111;
assign micromatrizz[39][118] = 9'b111111111;
assign micromatrizz[39][119] = 9'b111111111;
assign micromatrizz[39][120] = 9'b111111111;
assign micromatrizz[39][121] = 9'b111111111;
assign micromatrizz[39][122] = 9'b111111111;
assign micromatrizz[39][123] = 9'b111111111;
assign micromatrizz[39][124] = 9'b111111111;
assign micromatrizz[39][125] = 9'b111111111;
assign micromatrizz[39][126] = 9'b111111111;
assign micromatrizz[39][127] = 9'b111111111;
assign micromatrizz[39][128] = 9'b111111111;
assign micromatrizz[39][129] = 9'b111111111;
assign micromatrizz[39][130] = 9'b111111111;
assign micromatrizz[39][131] = 9'b111111111;
assign micromatrizz[39][132] = 9'b111111111;
assign micromatrizz[39][133] = 9'b111111111;
assign micromatrizz[39][134] = 9'b111111111;
assign micromatrizz[39][135] = 9'b111111111;
assign micromatrizz[39][136] = 9'b111111111;
assign micromatrizz[39][137] = 9'b111111111;
assign micromatrizz[39][138] = 9'b111111111;
assign micromatrizz[39][139] = 9'b111111111;
assign micromatrizz[39][140] = 9'b111111111;
assign micromatrizz[39][141] = 9'b111111111;
assign micromatrizz[39][142] = 9'b111111111;
assign micromatrizz[39][143] = 9'b111111111;
assign micromatrizz[39][144] = 9'b111111111;
assign micromatrizz[39][145] = 9'b111111111;
assign micromatrizz[39][146] = 9'b111111111;
assign micromatrizz[39][147] = 9'b111111111;
assign micromatrizz[39][148] = 9'b111111111;
assign micromatrizz[39][149] = 9'b111111111;
assign micromatrizz[39][150] = 9'b111111111;
assign micromatrizz[39][151] = 9'b111111111;
assign micromatrizz[39][152] = 9'b111111111;
assign micromatrizz[39][153] = 9'b111111111;
assign micromatrizz[39][154] = 9'b111111111;
assign micromatrizz[39][155] = 9'b111111111;
assign micromatrizz[39][156] = 9'b111111111;
assign micromatrizz[39][157] = 9'b111111111;
assign micromatrizz[39][158] = 9'b111111111;
assign micromatrizz[39][159] = 9'b111111111;
assign micromatrizz[39][160] = 9'b111111111;
assign micromatrizz[39][161] = 9'b111111111;
assign micromatrizz[39][162] = 9'b111111111;
assign micromatrizz[39][163] = 9'b111111111;
assign micromatrizz[39][164] = 9'b111111111;
assign micromatrizz[39][165] = 9'b111111111;
assign micromatrizz[39][166] = 9'b111111111;
assign micromatrizz[39][167] = 9'b111111111;
assign micromatrizz[39][168] = 9'b111111111;
assign micromatrizz[39][169] = 9'b111111111;
assign micromatrizz[39][170] = 9'b111111111;
assign micromatrizz[39][171] = 9'b111111111;
assign micromatrizz[39][172] = 9'b111111111;
assign micromatrizz[39][173] = 9'b111111111;
assign micromatrizz[39][174] = 9'b111111111;
assign micromatrizz[39][175] = 9'b111111111;
assign micromatrizz[39][176] = 9'b111111111;
assign micromatrizz[39][177] = 9'b111111111;
assign micromatrizz[39][178] = 9'b111111111;
assign micromatrizz[39][179] = 9'b111111111;
assign micromatrizz[39][180] = 9'b111111111;
assign micromatrizz[39][181] = 9'b111111111;
assign micromatrizz[39][182] = 9'b111111111;
assign micromatrizz[39][183] = 9'b111111111;
assign micromatrizz[39][184] = 9'b111111111;
assign micromatrizz[39][185] = 9'b111111111;
assign micromatrizz[39][186] = 9'b111111111;
assign micromatrizz[39][187] = 9'b111111111;
assign micromatrizz[39][188] = 9'b111111111;
assign micromatrizz[39][189] = 9'b111111111;
assign micromatrizz[39][190] = 9'b111111111;
assign micromatrizz[39][191] = 9'b111111111;
assign micromatrizz[39][192] = 9'b111111111;
assign micromatrizz[39][193] = 9'b111111111;
assign micromatrizz[39][194] = 9'b111111111;
assign micromatrizz[39][195] = 9'b111111111;
assign micromatrizz[39][196] = 9'b111111111;
assign micromatrizz[39][197] = 9'b111111111;
assign micromatrizz[39][198] = 9'b111111111;
assign micromatrizz[39][199] = 9'b111111111;
assign micromatrizz[39][200] = 9'b111111111;
assign micromatrizz[39][201] = 9'b111111111;
assign micromatrizz[39][202] = 9'b111111111;
assign micromatrizz[39][203] = 9'b111111111;
assign micromatrizz[39][204] = 9'b111111111;
assign micromatrizz[39][205] = 9'b111111111;
assign micromatrizz[39][206] = 9'b111111111;
assign micromatrizz[39][207] = 9'b111111111;
assign micromatrizz[39][208] = 9'b111111111;
assign micromatrizz[39][209] = 9'b111111111;
assign micromatrizz[39][210] = 9'b111111111;
assign micromatrizz[39][211] = 9'b111111111;
assign micromatrizz[39][212] = 9'b111111111;
assign micromatrizz[39][213] = 9'b111111111;
assign micromatrizz[39][214] = 9'b111111111;
assign micromatrizz[39][215] = 9'b111111111;
assign micromatrizz[39][216] = 9'b111111111;
assign micromatrizz[39][217] = 9'b111111111;
assign micromatrizz[39][218] = 9'b111111111;
assign micromatrizz[39][219] = 9'b111111111;
assign micromatrizz[39][220] = 9'b111111111;
assign micromatrizz[39][221] = 9'b111111111;
assign micromatrizz[39][222] = 9'b111111111;
assign micromatrizz[39][223] = 9'b111111111;
assign micromatrizz[39][224] = 9'b111111111;
assign micromatrizz[39][225] = 9'b111111111;
assign micromatrizz[39][226] = 9'b111111111;
assign micromatrizz[39][227] = 9'b111111111;
assign micromatrizz[39][228] = 9'b111111111;
assign micromatrizz[39][229] = 9'b111111111;
assign micromatrizz[39][230] = 9'b111111111;
assign micromatrizz[39][231] = 9'b111111111;
assign micromatrizz[39][232] = 9'b111111111;
assign micromatrizz[39][233] = 9'b111111111;
assign micromatrizz[39][234] = 9'b111111111;
assign micromatrizz[39][235] = 9'b111111111;
assign micromatrizz[39][236] = 9'b111111111;
assign micromatrizz[39][237] = 9'b111111111;
assign micromatrizz[39][238] = 9'b111111111;
assign micromatrizz[39][239] = 9'b111111111;
assign micromatrizz[39][240] = 9'b111111111;
assign micromatrizz[39][241] = 9'b111111111;
assign micromatrizz[39][242] = 9'b111111111;
assign micromatrizz[39][243] = 9'b111111111;
assign micromatrizz[39][244] = 9'b111111111;
assign micromatrizz[39][245] = 9'b111111111;
assign micromatrizz[39][246] = 9'b111111111;
assign micromatrizz[39][247] = 9'b111111111;
assign micromatrizz[39][248] = 9'b111111111;
assign micromatrizz[39][249] = 9'b111111111;
assign micromatrizz[39][250] = 9'b111111111;
assign micromatrizz[39][251] = 9'b111111111;
assign micromatrizz[39][252] = 9'b111111111;
assign micromatrizz[39][253] = 9'b111111111;
assign micromatrizz[39][254] = 9'b111111111;
assign micromatrizz[39][255] = 9'b111111111;
assign micromatrizz[39][256] = 9'b111111111;
assign micromatrizz[39][257] = 9'b111111111;
assign micromatrizz[39][258] = 9'b111111111;
assign micromatrizz[39][259] = 9'b111111111;
assign micromatrizz[39][260] = 9'b111111111;
assign micromatrizz[39][261] = 9'b111111111;
assign micromatrizz[39][262] = 9'b111111111;
assign micromatrizz[39][263] = 9'b111111111;
assign micromatrizz[39][264] = 9'b111111111;
assign micromatrizz[39][265] = 9'b111111111;
assign micromatrizz[39][266] = 9'b111111111;
assign micromatrizz[39][267] = 9'b111111111;
assign micromatrizz[39][268] = 9'b111111111;
assign micromatrizz[39][269] = 9'b111111111;
assign micromatrizz[39][270] = 9'b111111111;
assign micromatrizz[39][271] = 9'b111111111;
assign micromatrizz[39][272] = 9'b111111111;
assign micromatrizz[39][273] = 9'b111111111;
assign micromatrizz[39][274] = 9'b111111111;
assign micromatrizz[39][275] = 9'b111111111;
assign micromatrizz[39][276] = 9'b111111111;
assign micromatrizz[39][277] = 9'b111111111;
assign micromatrizz[39][278] = 9'b111111111;
assign micromatrizz[39][279] = 9'b111111111;
assign micromatrizz[39][280] = 9'b111111111;
assign micromatrizz[39][281] = 9'b111111111;
assign micromatrizz[39][282] = 9'b111111111;
assign micromatrizz[39][283] = 9'b111111111;
assign micromatrizz[39][284] = 9'b111111111;
assign micromatrizz[39][285] = 9'b111111111;
assign micromatrizz[39][286] = 9'b111111111;
assign micromatrizz[39][287] = 9'b111111111;
assign micromatrizz[39][288] = 9'b111111111;
assign micromatrizz[39][289] = 9'b111111111;
assign micromatrizz[39][290] = 9'b111111111;
assign micromatrizz[39][291] = 9'b111111111;
assign micromatrizz[39][292] = 9'b111111111;
assign micromatrizz[39][293] = 9'b111111111;
assign micromatrizz[39][294] = 9'b111111111;
assign micromatrizz[39][295] = 9'b111111111;
assign micromatrizz[39][296] = 9'b111111111;
assign micromatrizz[39][297] = 9'b111111111;
assign micromatrizz[39][298] = 9'b111111111;
assign micromatrizz[39][299] = 9'b111111111;
assign micromatrizz[39][300] = 9'b111111111;
assign micromatrizz[39][301] = 9'b111111111;
assign micromatrizz[39][302] = 9'b111111111;
assign micromatrizz[39][303] = 9'b111111111;
assign micromatrizz[39][304] = 9'b111111111;
assign micromatrizz[39][305] = 9'b111111111;
assign micromatrizz[39][306] = 9'b111111111;
assign micromatrizz[39][307] = 9'b111111111;
assign micromatrizz[39][308] = 9'b111111111;
assign micromatrizz[39][309] = 9'b111111111;
assign micromatrizz[39][310] = 9'b111111111;
assign micromatrizz[39][311] = 9'b111111111;
assign micromatrizz[39][312] = 9'b111111111;
assign micromatrizz[39][313] = 9'b111111111;
assign micromatrizz[39][314] = 9'b111111111;
assign micromatrizz[39][315] = 9'b111111111;
assign micromatrizz[39][316] = 9'b111111111;
assign micromatrizz[39][317] = 9'b111111111;
assign micromatrizz[39][318] = 9'b111111111;
assign micromatrizz[39][319] = 9'b111111111;
assign micromatrizz[39][320] = 9'b111111111;
assign micromatrizz[39][321] = 9'b111111111;
assign micromatrizz[39][322] = 9'b111111111;
assign micromatrizz[39][323] = 9'b111111111;
assign micromatrizz[39][324] = 9'b111111111;
assign micromatrizz[39][325] = 9'b111111111;
assign micromatrizz[39][326] = 9'b111111111;
assign micromatrizz[39][327] = 9'b111111111;
assign micromatrizz[39][328] = 9'b111111111;
assign micromatrizz[39][329] = 9'b111111111;
assign micromatrizz[39][330] = 9'b111111111;
assign micromatrizz[39][331] = 9'b111111111;
assign micromatrizz[39][332] = 9'b111111111;
assign micromatrizz[39][333] = 9'b111111111;
assign micromatrizz[39][334] = 9'b111111111;
assign micromatrizz[39][335] = 9'b111111111;
assign micromatrizz[39][336] = 9'b111111111;
assign micromatrizz[39][337] = 9'b111111111;
assign micromatrizz[39][338] = 9'b111111111;
assign micromatrizz[39][339] = 9'b111111111;
assign micromatrizz[39][340] = 9'b111111111;
assign micromatrizz[39][341] = 9'b111111111;
assign micromatrizz[39][342] = 9'b111111111;
assign micromatrizz[39][343] = 9'b111111111;
assign micromatrizz[39][344] = 9'b111111111;
assign micromatrizz[39][345] = 9'b111111111;
assign micromatrizz[39][346] = 9'b111111111;
assign micromatrizz[39][347] = 9'b111111111;
assign micromatrizz[39][348] = 9'b111111111;
assign micromatrizz[39][349] = 9'b111111111;
assign micromatrizz[39][350] = 9'b111111111;
assign micromatrizz[39][351] = 9'b111111111;
assign micromatrizz[39][352] = 9'b111111111;
assign micromatrizz[39][353] = 9'b111111111;
assign micromatrizz[39][354] = 9'b111111111;
assign micromatrizz[39][355] = 9'b111111111;
assign micromatrizz[39][356] = 9'b111111111;
assign micromatrizz[39][357] = 9'b111111111;
assign micromatrizz[39][358] = 9'b111111111;
assign micromatrizz[39][359] = 9'b111111111;
assign micromatrizz[39][360] = 9'b111111111;
assign micromatrizz[39][361] = 9'b111111111;
assign micromatrizz[39][362] = 9'b111111111;
assign micromatrizz[39][363] = 9'b111111111;
assign micromatrizz[39][364] = 9'b111111111;
assign micromatrizz[39][365] = 9'b111111111;
assign micromatrizz[39][366] = 9'b111111111;
assign micromatrizz[39][367] = 9'b111111111;
assign micromatrizz[39][368] = 9'b111111111;
assign micromatrizz[39][369] = 9'b111111111;
assign micromatrizz[39][370] = 9'b111111111;
assign micromatrizz[39][371] = 9'b111111111;
assign micromatrizz[39][372] = 9'b111111111;
assign micromatrizz[39][373] = 9'b111111111;
assign micromatrizz[39][374] = 9'b111111111;
assign micromatrizz[39][375] = 9'b111111111;
assign micromatrizz[39][376] = 9'b111111111;
assign micromatrizz[39][377] = 9'b111111111;
assign micromatrizz[39][378] = 9'b111111111;
assign micromatrizz[39][379] = 9'b111111111;
assign micromatrizz[39][380] = 9'b111111111;
assign micromatrizz[39][381] = 9'b111111111;
assign micromatrizz[39][382] = 9'b111111111;
assign micromatrizz[39][383] = 9'b111111111;
assign micromatrizz[39][384] = 9'b111111111;
assign micromatrizz[39][385] = 9'b111111111;
assign micromatrizz[39][386] = 9'b111111111;
assign micromatrizz[39][387] = 9'b111111111;
assign micromatrizz[39][388] = 9'b111111111;
assign micromatrizz[39][389] = 9'b111111111;
assign micromatrizz[39][390] = 9'b111111111;
assign micromatrizz[39][391] = 9'b111111111;
assign micromatrizz[39][392] = 9'b111111111;
assign micromatrizz[39][393] = 9'b111111111;
assign micromatrizz[39][394] = 9'b111111111;
assign micromatrizz[39][395] = 9'b111111111;
assign micromatrizz[39][396] = 9'b111111111;
assign micromatrizz[39][397] = 9'b111111111;
assign micromatrizz[39][398] = 9'b111111111;
assign micromatrizz[39][399] = 9'b111111111;
assign micromatrizz[39][400] = 9'b111111111;
assign micromatrizz[39][401] = 9'b111111111;
assign micromatrizz[39][402] = 9'b111111111;
assign micromatrizz[39][403] = 9'b111111111;
assign micromatrizz[39][404] = 9'b111111111;
assign micromatrizz[39][405] = 9'b111111111;
assign micromatrizz[39][406] = 9'b111111111;
assign micromatrizz[39][407] = 9'b111111111;
assign micromatrizz[39][408] = 9'b111111111;
assign micromatrizz[39][409] = 9'b111111111;
assign micromatrizz[39][410] = 9'b111111111;
assign micromatrizz[39][411] = 9'b111111111;
assign micromatrizz[39][412] = 9'b111111111;
assign micromatrizz[39][413] = 9'b111111111;
assign micromatrizz[39][414] = 9'b111111111;
assign micromatrizz[39][415] = 9'b111111111;
assign micromatrizz[39][416] = 9'b111111111;
assign micromatrizz[39][417] = 9'b111111111;
assign micromatrizz[39][418] = 9'b111111111;
assign micromatrizz[39][419] = 9'b111111111;
assign micromatrizz[39][420] = 9'b111111111;
assign micromatrizz[39][421] = 9'b111111111;
assign micromatrizz[39][422] = 9'b111111111;
assign micromatrizz[39][423] = 9'b111111111;
assign micromatrizz[39][424] = 9'b111111111;
assign micromatrizz[39][425] = 9'b111111111;
assign micromatrizz[39][426] = 9'b111111111;
assign micromatrizz[39][427] = 9'b111111111;
assign micromatrizz[39][428] = 9'b111111111;
assign micromatrizz[39][429] = 9'b111111111;
assign micromatrizz[39][430] = 9'b111111111;
assign micromatrizz[39][431] = 9'b111111111;
assign micromatrizz[39][432] = 9'b111111111;
assign micromatrizz[39][433] = 9'b111111111;
assign micromatrizz[39][434] = 9'b111111111;
assign micromatrizz[39][435] = 9'b111111111;
assign micromatrizz[39][436] = 9'b111111111;
assign micromatrizz[39][437] = 9'b111111111;
assign micromatrizz[39][438] = 9'b111111111;
assign micromatrizz[39][439] = 9'b111111111;
assign micromatrizz[39][440] = 9'b111111111;
assign micromatrizz[39][441] = 9'b111111111;
assign micromatrizz[39][442] = 9'b111111111;
assign micromatrizz[39][443] = 9'b111111111;
assign micromatrizz[39][444] = 9'b111111111;
assign micromatrizz[39][445] = 9'b111111111;
assign micromatrizz[39][446] = 9'b111111111;
assign micromatrizz[39][447] = 9'b111111111;
assign micromatrizz[39][448] = 9'b111111111;
assign micromatrizz[39][449] = 9'b111111111;
assign micromatrizz[39][450] = 9'b111111111;
assign micromatrizz[39][451] = 9'b111111111;
assign micromatrizz[39][452] = 9'b111111111;
assign micromatrizz[39][453] = 9'b111111111;
assign micromatrizz[39][454] = 9'b111111111;
assign micromatrizz[39][455] = 9'b111111111;
assign micromatrizz[39][456] = 9'b111111111;
assign micromatrizz[39][457] = 9'b111111111;
assign micromatrizz[39][458] = 9'b111111111;
assign micromatrizz[39][459] = 9'b111111111;
assign micromatrizz[39][460] = 9'b111111111;
assign micromatrizz[39][461] = 9'b111111111;
assign micromatrizz[39][462] = 9'b111111111;
assign micromatrizz[39][463] = 9'b111111111;
assign micromatrizz[39][464] = 9'b111111111;
assign micromatrizz[39][465] = 9'b111111111;
assign micromatrizz[39][466] = 9'b111111111;
assign micromatrizz[39][467] = 9'b111111111;
assign micromatrizz[39][468] = 9'b111111111;
assign micromatrizz[39][469] = 9'b111111111;
assign micromatrizz[39][470] = 9'b111111111;
assign micromatrizz[39][471] = 9'b111111111;
assign micromatrizz[39][472] = 9'b111111111;
assign micromatrizz[39][473] = 9'b111111111;
assign micromatrizz[39][474] = 9'b111111111;
assign micromatrizz[39][475] = 9'b111111111;
assign micromatrizz[39][476] = 9'b111111111;
assign micromatrizz[39][477] = 9'b111111111;
assign micromatrizz[39][478] = 9'b111111111;
assign micromatrizz[39][479] = 9'b111111111;
assign micromatrizz[39][480] = 9'b111111111;
assign micromatrizz[39][481] = 9'b111111111;
assign micromatrizz[39][482] = 9'b111111111;
assign micromatrizz[39][483] = 9'b111111111;
assign micromatrizz[39][484] = 9'b111111111;
assign micromatrizz[39][485] = 9'b111111111;
assign micromatrizz[39][486] = 9'b111111111;
assign micromatrizz[39][487] = 9'b111111111;
assign micromatrizz[39][488] = 9'b111111111;
assign micromatrizz[39][489] = 9'b111111111;
assign micromatrizz[39][490] = 9'b111111111;
assign micromatrizz[39][491] = 9'b111111111;
assign micromatrizz[39][492] = 9'b111111111;
assign micromatrizz[39][493] = 9'b111111111;
assign micromatrizz[39][494] = 9'b111111111;
assign micromatrizz[39][495] = 9'b111111111;
assign micromatrizz[39][496] = 9'b111111111;
assign micromatrizz[39][497] = 9'b111111111;
assign micromatrizz[39][498] = 9'b111111111;
assign micromatrizz[39][499] = 9'b111111111;
assign micromatrizz[39][500] = 9'b111111111;
assign micromatrizz[39][501] = 9'b111111111;
assign micromatrizz[39][502] = 9'b111111111;
assign micromatrizz[39][503] = 9'b111111111;
assign micromatrizz[39][504] = 9'b111111111;
assign micromatrizz[39][505] = 9'b111111111;
assign micromatrizz[39][506] = 9'b111111111;
assign micromatrizz[39][507] = 9'b111111111;
assign micromatrizz[39][508] = 9'b111111111;
assign micromatrizz[39][509] = 9'b111111111;
assign micromatrizz[39][510] = 9'b111111111;
assign micromatrizz[39][511] = 9'b111111111;
assign micromatrizz[39][512] = 9'b111111111;
assign micromatrizz[39][513] = 9'b111111111;
assign micromatrizz[39][514] = 9'b111111111;
assign micromatrizz[39][515] = 9'b111111111;
assign micromatrizz[39][516] = 9'b111111111;
assign micromatrizz[39][517] = 9'b111111111;
assign micromatrizz[39][518] = 9'b111111111;
assign micromatrizz[39][519] = 9'b111111111;
assign micromatrizz[39][520] = 9'b111111111;
assign micromatrizz[39][521] = 9'b111111111;
assign micromatrizz[39][522] = 9'b111111111;
assign micromatrizz[39][523] = 9'b111111111;
assign micromatrizz[39][524] = 9'b111111111;
assign micromatrizz[39][525] = 9'b111111111;
assign micromatrizz[39][526] = 9'b111111111;
assign micromatrizz[39][527] = 9'b111111111;
assign micromatrizz[39][528] = 9'b111111111;
assign micromatrizz[39][529] = 9'b111111111;
assign micromatrizz[39][530] = 9'b111111111;
assign micromatrizz[39][531] = 9'b111111111;
assign micromatrizz[39][532] = 9'b111111111;
assign micromatrizz[39][533] = 9'b111111111;
assign micromatrizz[39][534] = 9'b111111111;
assign micromatrizz[39][535] = 9'b111111111;
assign micromatrizz[39][536] = 9'b111111111;
assign micromatrizz[39][537] = 9'b111111111;
assign micromatrizz[39][538] = 9'b111111111;
assign micromatrizz[39][539] = 9'b111111111;
assign micromatrizz[39][540] = 9'b111111111;
assign micromatrizz[39][541] = 9'b111111111;
assign micromatrizz[39][542] = 9'b111111111;
assign micromatrizz[39][543] = 9'b111111111;
assign micromatrizz[39][544] = 9'b111111111;
assign micromatrizz[39][545] = 9'b111111111;
assign micromatrizz[39][546] = 9'b111111111;
assign micromatrizz[39][547] = 9'b111111111;
assign micromatrizz[39][548] = 9'b111111111;
assign micromatrizz[39][549] = 9'b111111111;
assign micromatrizz[39][550] = 9'b111111111;
assign micromatrizz[39][551] = 9'b111111111;
assign micromatrizz[39][552] = 9'b111111111;
assign micromatrizz[39][553] = 9'b111111111;
assign micromatrizz[39][554] = 9'b111111111;
assign micromatrizz[39][555] = 9'b111111111;
assign micromatrizz[39][556] = 9'b111111111;
assign micromatrizz[39][557] = 9'b111111111;
assign micromatrizz[39][558] = 9'b111111111;
assign micromatrizz[39][559] = 9'b111111111;
assign micromatrizz[39][560] = 9'b111111111;
assign micromatrizz[39][561] = 9'b111111111;
assign micromatrizz[39][562] = 9'b111111111;
assign micromatrizz[39][563] = 9'b111111111;
assign micromatrizz[39][564] = 9'b111111111;
assign micromatrizz[39][565] = 9'b111111111;
assign micromatrizz[39][566] = 9'b111111111;
assign micromatrizz[39][567] = 9'b111111111;
assign micromatrizz[39][568] = 9'b111111111;
assign micromatrizz[39][569] = 9'b111111111;
assign micromatrizz[39][570] = 9'b111111111;
assign micromatrizz[39][571] = 9'b111111111;
assign micromatrizz[39][572] = 9'b111111111;
assign micromatrizz[39][573] = 9'b111111111;
assign micromatrizz[39][574] = 9'b111111111;
assign micromatrizz[39][575] = 9'b111111111;
assign micromatrizz[39][576] = 9'b111111111;
assign micromatrizz[39][577] = 9'b111111111;
assign micromatrizz[39][578] = 9'b111111111;
assign micromatrizz[39][579] = 9'b111111111;
assign micromatrizz[39][580] = 9'b111111111;
assign micromatrizz[39][581] = 9'b111111111;
assign micromatrizz[39][582] = 9'b111111111;
assign micromatrizz[39][583] = 9'b111111111;
assign micromatrizz[39][584] = 9'b111111111;
assign micromatrizz[39][585] = 9'b111111111;
assign micromatrizz[39][586] = 9'b111111111;
assign micromatrizz[39][587] = 9'b111111111;
assign micromatrizz[39][588] = 9'b111111111;
assign micromatrizz[39][589] = 9'b111111111;
assign micromatrizz[39][590] = 9'b111111111;
assign micromatrizz[39][591] = 9'b111111111;
assign micromatrizz[39][592] = 9'b111111111;
assign micromatrizz[39][593] = 9'b111111111;
assign micromatrizz[39][594] = 9'b111111111;
assign micromatrizz[39][595] = 9'b111111111;
assign micromatrizz[39][596] = 9'b111111111;
assign micromatrizz[39][597] = 9'b111111111;
assign micromatrizz[39][598] = 9'b111111111;
assign micromatrizz[39][599] = 9'b111111111;
assign micromatrizz[39][600] = 9'b111111111;
assign micromatrizz[39][601] = 9'b111111111;
assign micromatrizz[39][602] = 9'b111111111;
assign micromatrizz[39][603] = 9'b111111111;
assign micromatrizz[39][604] = 9'b111111111;
assign micromatrizz[39][605] = 9'b111111111;
assign micromatrizz[39][606] = 9'b111111111;
assign micromatrizz[39][607] = 9'b111111111;
assign micromatrizz[39][608] = 9'b111111111;
assign micromatrizz[39][609] = 9'b111111111;
assign micromatrizz[39][610] = 9'b111111111;
assign micromatrizz[39][611] = 9'b111111111;
assign micromatrizz[39][612] = 9'b111111111;
assign micromatrizz[39][613] = 9'b111111111;
assign micromatrizz[39][614] = 9'b111111111;
assign micromatrizz[39][615] = 9'b111111111;
assign micromatrizz[39][616] = 9'b111111111;
assign micromatrizz[39][617] = 9'b111111111;
assign micromatrizz[39][618] = 9'b111111111;
assign micromatrizz[39][619] = 9'b111111111;
assign micromatrizz[39][620] = 9'b111111111;
assign micromatrizz[39][621] = 9'b111111111;
assign micromatrizz[39][622] = 9'b111111111;
assign micromatrizz[39][623] = 9'b111111111;
assign micromatrizz[39][624] = 9'b111111111;
assign micromatrizz[39][625] = 9'b111111111;
assign micromatrizz[39][626] = 9'b111111111;
assign micromatrizz[39][627] = 9'b111111111;
assign micromatrizz[39][628] = 9'b111111111;
assign micromatrizz[39][629] = 9'b111111111;
assign micromatrizz[39][630] = 9'b111111111;
assign micromatrizz[39][631] = 9'b111111111;
assign micromatrizz[39][632] = 9'b111111111;
assign micromatrizz[39][633] = 9'b111111111;
assign micromatrizz[39][634] = 9'b111111111;
assign micromatrizz[39][635] = 9'b111111111;
assign micromatrizz[39][636] = 9'b111111111;
assign micromatrizz[39][637] = 9'b111111111;
assign micromatrizz[39][638] = 9'b111111111;
assign micromatrizz[39][639] = 9'b111111111;
assign micromatrizz[40][0] = 9'b111111111;
assign micromatrizz[40][1] = 9'b111111111;
assign micromatrizz[40][2] = 9'b111111111;
assign micromatrizz[40][3] = 9'b111111111;
assign micromatrizz[40][4] = 9'b111111111;
assign micromatrizz[40][5] = 9'b111111111;
assign micromatrizz[40][6] = 9'b111111111;
assign micromatrizz[40][7] = 9'b111111111;
assign micromatrizz[40][8] = 9'b111111111;
assign micromatrizz[40][9] = 9'b111111111;
assign micromatrizz[40][10] = 9'b111111111;
assign micromatrizz[40][11] = 9'b111111111;
assign micromatrizz[40][12] = 9'b111111111;
assign micromatrizz[40][13] = 9'b111111111;
assign micromatrizz[40][14] = 9'b111111111;
assign micromatrizz[40][15] = 9'b111111111;
assign micromatrizz[40][16] = 9'b111111111;
assign micromatrizz[40][17] = 9'b111111111;
assign micromatrizz[40][18] = 9'b111111111;
assign micromatrizz[40][19] = 9'b111111111;
assign micromatrizz[40][20] = 9'b111111111;
assign micromatrizz[40][21] = 9'b111111111;
assign micromatrizz[40][22] = 9'b111111111;
assign micromatrizz[40][23] = 9'b111111111;
assign micromatrizz[40][24] = 9'b111111111;
assign micromatrizz[40][25] = 9'b111111111;
assign micromatrizz[40][26] = 9'b111111111;
assign micromatrizz[40][27] = 9'b111111111;
assign micromatrizz[40][28] = 9'b111111111;
assign micromatrizz[40][29] = 9'b111111111;
assign micromatrizz[40][30] = 9'b111111111;
assign micromatrizz[40][31] = 9'b111111111;
assign micromatrizz[40][32] = 9'b111111111;
assign micromatrizz[40][33] = 9'b111111111;
assign micromatrizz[40][34] = 9'b111111111;
assign micromatrizz[40][35] = 9'b111111111;
assign micromatrizz[40][36] = 9'b111111111;
assign micromatrizz[40][37] = 9'b111111111;
assign micromatrizz[40][38] = 9'b111111111;
assign micromatrizz[40][39] = 9'b111111111;
assign micromatrizz[40][40] = 9'b111111111;
assign micromatrizz[40][41] = 9'b111111111;
assign micromatrizz[40][42] = 9'b111111111;
assign micromatrizz[40][43] = 9'b111111111;
assign micromatrizz[40][44] = 9'b111111111;
assign micromatrizz[40][45] = 9'b111111111;
assign micromatrizz[40][46] = 9'b111111111;
assign micromatrizz[40][47] = 9'b111111111;
assign micromatrizz[40][48] = 9'b111111111;
assign micromatrizz[40][49] = 9'b111111111;
assign micromatrizz[40][50] = 9'b111111111;
assign micromatrizz[40][51] = 9'b111111111;
assign micromatrizz[40][52] = 9'b111111111;
assign micromatrizz[40][53] = 9'b111111111;
assign micromatrizz[40][54] = 9'b111111111;
assign micromatrizz[40][55] = 9'b111111111;
assign micromatrizz[40][56] = 9'b111111111;
assign micromatrizz[40][57] = 9'b111111111;
assign micromatrizz[40][58] = 9'b111111111;
assign micromatrizz[40][59] = 9'b111111111;
assign micromatrizz[40][60] = 9'b111111111;
assign micromatrizz[40][61] = 9'b111111111;
assign micromatrizz[40][62] = 9'b111111111;
assign micromatrizz[40][63] = 9'b111111111;
assign micromatrizz[40][64] = 9'b111111111;
assign micromatrizz[40][65] = 9'b111111111;
assign micromatrizz[40][66] = 9'b111111111;
assign micromatrizz[40][67] = 9'b111111111;
assign micromatrizz[40][68] = 9'b111111111;
assign micromatrizz[40][69] = 9'b111111111;
assign micromatrizz[40][70] = 9'b111111111;
assign micromatrizz[40][71] = 9'b111111111;
assign micromatrizz[40][72] = 9'b111111111;
assign micromatrizz[40][73] = 9'b111111111;
assign micromatrizz[40][74] = 9'b111111111;
assign micromatrizz[40][75] = 9'b111111111;
assign micromatrizz[40][76] = 9'b111111111;
assign micromatrizz[40][77] = 9'b111111111;
assign micromatrizz[40][78] = 9'b111111111;
assign micromatrizz[40][79] = 9'b111111111;
assign micromatrizz[40][80] = 9'b111111111;
assign micromatrizz[40][81] = 9'b111111111;
assign micromatrizz[40][82] = 9'b111111111;
assign micromatrizz[40][83] = 9'b111111111;
assign micromatrizz[40][84] = 9'b111111111;
assign micromatrizz[40][85] = 9'b111111111;
assign micromatrizz[40][86] = 9'b111111111;
assign micromatrizz[40][87] = 9'b111111111;
assign micromatrizz[40][88] = 9'b111111111;
assign micromatrizz[40][89] = 9'b111111111;
assign micromatrizz[40][90] = 9'b111111111;
assign micromatrizz[40][91] = 9'b111111111;
assign micromatrizz[40][92] = 9'b111111111;
assign micromatrizz[40][93] = 9'b111111111;
assign micromatrizz[40][94] = 9'b111111111;
assign micromatrizz[40][95] = 9'b111111111;
assign micromatrizz[40][96] = 9'b111111111;
assign micromatrizz[40][97] = 9'b111111111;
assign micromatrizz[40][98] = 9'b111111111;
assign micromatrizz[40][99] = 9'b111111111;
assign micromatrizz[40][100] = 9'b111111111;
assign micromatrizz[40][101] = 9'b111111111;
assign micromatrizz[40][102] = 9'b111111111;
assign micromatrizz[40][103] = 9'b111111111;
assign micromatrizz[40][104] = 9'b111111111;
assign micromatrizz[40][105] = 9'b111111111;
assign micromatrizz[40][106] = 9'b111111111;
assign micromatrizz[40][107] = 9'b111111111;
assign micromatrizz[40][108] = 9'b111111111;
assign micromatrizz[40][109] = 9'b111111111;
assign micromatrizz[40][110] = 9'b111111111;
assign micromatrizz[40][111] = 9'b111111111;
assign micromatrizz[40][112] = 9'b111111111;
assign micromatrizz[40][113] = 9'b111111111;
assign micromatrizz[40][114] = 9'b111111111;
assign micromatrizz[40][115] = 9'b111111111;
assign micromatrizz[40][116] = 9'b111111111;
assign micromatrizz[40][117] = 9'b111111111;
assign micromatrizz[40][118] = 9'b111111111;
assign micromatrizz[40][119] = 9'b111111111;
assign micromatrizz[40][120] = 9'b111111111;
assign micromatrizz[40][121] = 9'b111111111;
assign micromatrizz[40][122] = 9'b111111111;
assign micromatrizz[40][123] = 9'b111111111;
assign micromatrizz[40][124] = 9'b111111111;
assign micromatrizz[40][125] = 9'b111111111;
assign micromatrizz[40][126] = 9'b111111111;
assign micromatrizz[40][127] = 9'b111111111;
assign micromatrizz[40][128] = 9'b111111111;
assign micromatrizz[40][129] = 9'b111111111;
assign micromatrizz[40][130] = 9'b111111111;
assign micromatrizz[40][131] = 9'b111111111;
assign micromatrizz[40][132] = 9'b111111111;
assign micromatrizz[40][133] = 9'b111111111;
assign micromatrizz[40][134] = 9'b111111111;
assign micromatrizz[40][135] = 9'b111111111;
assign micromatrizz[40][136] = 9'b111111111;
assign micromatrizz[40][137] = 9'b111111111;
assign micromatrizz[40][138] = 9'b111111111;
assign micromatrizz[40][139] = 9'b111111111;
assign micromatrizz[40][140] = 9'b111111111;
assign micromatrizz[40][141] = 9'b111111111;
assign micromatrizz[40][142] = 9'b111111111;
assign micromatrizz[40][143] = 9'b111111111;
assign micromatrizz[40][144] = 9'b111111111;
assign micromatrizz[40][145] = 9'b111111111;
assign micromatrizz[40][146] = 9'b111111111;
assign micromatrizz[40][147] = 9'b111111111;
assign micromatrizz[40][148] = 9'b111111111;
assign micromatrizz[40][149] = 9'b111111111;
assign micromatrizz[40][150] = 9'b111111111;
assign micromatrizz[40][151] = 9'b111111111;
assign micromatrizz[40][152] = 9'b111111111;
assign micromatrizz[40][153] = 9'b111111111;
assign micromatrizz[40][154] = 9'b111111111;
assign micromatrizz[40][155] = 9'b111111111;
assign micromatrizz[40][156] = 9'b111111111;
assign micromatrizz[40][157] = 9'b111111111;
assign micromatrizz[40][158] = 9'b111111111;
assign micromatrizz[40][159] = 9'b111111111;
assign micromatrizz[40][160] = 9'b111111111;
assign micromatrizz[40][161] = 9'b111111111;
assign micromatrizz[40][162] = 9'b111111111;
assign micromatrizz[40][163] = 9'b111111111;
assign micromatrizz[40][164] = 9'b111111111;
assign micromatrizz[40][165] = 9'b111111111;
assign micromatrizz[40][166] = 9'b111111111;
assign micromatrizz[40][167] = 9'b111111111;
assign micromatrizz[40][168] = 9'b111111111;
assign micromatrizz[40][169] = 9'b111111111;
assign micromatrizz[40][170] = 9'b111111111;
assign micromatrizz[40][171] = 9'b111111111;
assign micromatrizz[40][172] = 9'b111111111;
assign micromatrizz[40][173] = 9'b111111111;
assign micromatrizz[40][174] = 9'b111111111;
assign micromatrizz[40][175] = 9'b111111111;
assign micromatrizz[40][176] = 9'b111111111;
assign micromatrizz[40][177] = 9'b111111111;
assign micromatrizz[40][178] = 9'b111111111;
assign micromatrizz[40][179] = 9'b111111111;
assign micromatrizz[40][180] = 9'b111111111;
assign micromatrizz[40][181] = 9'b111111111;
assign micromatrizz[40][182] = 9'b111111111;
assign micromatrizz[40][183] = 9'b111111111;
assign micromatrizz[40][184] = 9'b111111111;
assign micromatrizz[40][185] = 9'b111111111;
assign micromatrizz[40][186] = 9'b111111111;
assign micromatrizz[40][187] = 9'b111111111;
assign micromatrizz[40][188] = 9'b111111111;
assign micromatrizz[40][189] = 9'b111111111;
assign micromatrizz[40][190] = 9'b111111111;
assign micromatrizz[40][191] = 9'b111111111;
assign micromatrizz[40][192] = 9'b111111111;
assign micromatrizz[40][193] = 9'b111111111;
assign micromatrizz[40][194] = 9'b111111111;
assign micromatrizz[40][195] = 9'b111111111;
assign micromatrizz[40][196] = 9'b111111111;
assign micromatrizz[40][197] = 9'b111111111;
assign micromatrizz[40][198] = 9'b111111111;
assign micromatrizz[40][199] = 9'b111111111;
assign micromatrizz[40][200] = 9'b111111111;
assign micromatrizz[40][201] = 9'b111111111;
assign micromatrizz[40][202] = 9'b111111111;
assign micromatrizz[40][203] = 9'b111111111;
assign micromatrizz[40][204] = 9'b111111111;
assign micromatrizz[40][205] = 9'b111111111;
assign micromatrizz[40][206] = 9'b111111111;
assign micromatrizz[40][207] = 9'b111111111;
assign micromatrizz[40][208] = 9'b111111111;
assign micromatrizz[40][209] = 9'b111111111;
assign micromatrizz[40][210] = 9'b111111111;
assign micromatrizz[40][211] = 9'b111111111;
assign micromatrizz[40][212] = 9'b111111111;
assign micromatrizz[40][213] = 9'b111111111;
assign micromatrizz[40][214] = 9'b111111111;
assign micromatrizz[40][215] = 9'b111111111;
assign micromatrizz[40][216] = 9'b111111111;
assign micromatrizz[40][217] = 9'b111111111;
assign micromatrizz[40][218] = 9'b111111111;
assign micromatrizz[40][219] = 9'b111111111;
assign micromatrizz[40][220] = 9'b111111111;
assign micromatrizz[40][221] = 9'b111111111;
assign micromatrizz[40][222] = 9'b111111111;
assign micromatrizz[40][223] = 9'b111111111;
assign micromatrizz[40][224] = 9'b111111111;
assign micromatrizz[40][225] = 9'b111111111;
assign micromatrizz[40][226] = 9'b111111111;
assign micromatrizz[40][227] = 9'b111111111;
assign micromatrizz[40][228] = 9'b111111111;
assign micromatrizz[40][229] = 9'b111111111;
assign micromatrizz[40][230] = 9'b111111111;
assign micromatrizz[40][231] = 9'b111111111;
assign micromatrizz[40][232] = 9'b111111111;
assign micromatrizz[40][233] = 9'b111111111;
assign micromatrizz[40][234] = 9'b111111111;
assign micromatrizz[40][235] = 9'b111111111;
assign micromatrizz[40][236] = 9'b111111111;
assign micromatrizz[40][237] = 9'b111111111;
assign micromatrizz[40][238] = 9'b111111111;
assign micromatrizz[40][239] = 9'b111111111;
assign micromatrizz[40][240] = 9'b111111111;
assign micromatrizz[40][241] = 9'b111111111;
assign micromatrizz[40][242] = 9'b111111111;
assign micromatrizz[40][243] = 9'b111111111;
assign micromatrizz[40][244] = 9'b111111111;
assign micromatrizz[40][245] = 9'b111111111;
assign micromatrizz[40][246] = 9'b111111111;
assign micromatrizz[40][247] = 9'b111111111;
assign micromatrizz[40][248] = 9'b111111111;
assign micromatrizz[40][249] = 9'b111111111;
assign micromatrizz[40][250] = 9'b111111111;
assign micromatrizz[40][251] = 9'b111111111;
assign micromatrizz[40][252] = 9'b111111111;
assign micromatrizz[40][253] = 9'b111111111;
assign micromatrizz[40][254] = 9'b111111111;
assign micromatrizz[40][255] = 9'b111111111;
assign micromatrizz[40][256] = 9'b111111111;
assign micromatrizz[40][257] = 9'b111111111;
assign micromatrizz[40][258] = 9'b111111111;
assign micromatrizz[40][259] = 9'b111111111;
assign micromatrizz[40][260] = 9'b111111111;
assign micromatrizz[40][261] = 9'b111111111;
assign micromatrizz[40][262] = 9'b111111111;
assign micromatrizz[40][263] = 9'b111111111;
assign micromatrizz[40][264] = 9'b111111111;
assign micromatrizz[40][265] = 9'b111111111;
assign micromatrizz[40][266] = 9'b111111111;
assign micromatrizz[40][267] = 9'b111111111;
assign micromatrizz[40][268] = 9'b111111111;
assign micromatrizz[40][269] = 9'b111111111;
assign micromatrizz[40][270] = 9'b111111111;
assign micromatrizz[40][271] = 9'b111111111;
assign micromatrizz[40][272] = 9'b111111111;
assign micromatrizz[40][273] = 9'b111111111;
assign micromatrizz[40][274] = 9'b111111111;
assign micromatrizz[40][275] = 9'b111111111;
assign micromatrizz[40][276] = 9'b111111111;
assign micromatrizz[40][277] = 9'b111111111;
assign micromatrizz[40][278] = 9'b111111111;
assign micromatrizz[40][279] = 9'b111111111;
assign micromatrizz[40][280] = 9'b111111111;
assign micromatrizz[40][281] = 9'b111111111;
assign micromatrizz[40][282] = 9'b111111111;
assign micromatrizz[40][283] = 9'b111111111;
assign micromatrizz[40][284] = 9'b111111111;
assign micromatrizz[40][285] = 9'b111111111;
assign micromatrizz[40][286] = 9'b111111111;
assign micromatrizz[40][287] = 9'b111111111;
assign micromatrizz[40][288] = 9'b111111111;
assign micromatrizz[40][289] = 9'b111111111;
assign micromatrizz[40][290] = 9'b111111111;
assign micromatrizz[40][291] = 9'b111111111;
assign micromatrizz[40][292] = 9'b111111111;
assign micromatrizz[40][293] = 9'b111111111;
assign micromatrizz[40][294] = 9'b111111111;
assign micromatrizz[40][295] = 9'b111111111;
assign micromatrizz[40][296] = 9'b111111111;
assign micromatrizz[40][297] = 9'b111111111;
assign micromatrizz[40][298] = 9'b111111111;
assign micromatrizz[40][299] = 9'b111111111;
assign micromatrizz[40][300] = 9'b111111111;
assign micromatrizz[40][301] = 9'b111111111;
assign micromatrizz[40][302] = 9'b111111111;
assign micromatrizz[40][303] = 9'b111111111;
assign micromatrizz[40][304] = 9'b111111111;
assign micromatrizz[40][305] = 9'b111111111;
assign micromatrizz[40][306] = 9'b111111111;
assign micromatrizz[40][307] = 9'b111111111;
assign micromatrizz[40][308] = 9'b111111111;
assign micromatrizz[40][309] = 9'b111111111;
assign micromatrizz[40][310] = 9'b111111111;
assign micromatrizz[40][311] = 9'b111111111;
assign micromatrizz[40][312] = 9'b111111111;
assign micromatrizz[40][313] = 9'b111111111;
assign micromatrizz[40][314] = 9'b111111111;
assign micromatrizz[40][315] = 9'b111111111;
assign micromatrizz[40][316] = 9'b111111111;
assign micromatrizz[40][317] = 9'b111111111;
assign micromatrizz[40][318] = 9'b111111111;
assign micromatrizz[40][319] = 9'b111111111;
assign micromatrizz[40][320] = 9'b111111111;
assign micromatrizz[40][321] = 9'b111111111;
assign micromatrizz[40][322] = 9'b111111111;
assign micromatrizz[40][323] = 9'b111111111;
assign micromatrizz[40][324] = 9'b111111111;
assign micromatrizz[40][325] = 9'b111111111;
assign micromatrizz[40][326] = 9'b111111111;
assign micromatrizz[40][327] = 9'b111111111;
assign micromatrizz[40][328] = 9'b111111111;
assign micromatrizz[40][329] = 9'b111111111;
assign micromatrizz[40][330] = 9'b111111111;
assign micromatrizz[40][331] = 9'b111111111;
assign micromatrizz[40][332] = 9'b111111111;
assign micromatrizz[40][333] = 9'b111111111;
assign micromatrizz[40][334] = 9'b111111111;
assign micromatrizz[40][335] = 9'b111111111;
assign micromatrizz[40][336] = 9'b111111111;
assign micromatrizz[40][337] = 9'b111111111;
assign micromatrizz[40][338] = 9'b111111111;
assign micromatrizz[40][339] = 9'b111111111;
assign micromatrizz[40][340] = 9'b111111111;
assign micromatrizz[40][341] = 9'b111111111;
assign micromatrizz[40][342] = 9'b111111111;
assign micromatrizz[40][343] = 9'b111111111;
assign micromatrizz[40][344] = 9'b111111111;
assign micromatrizz[40][345] = 9'b111111111;
assign micromatrizz[40][346] = 9'b111111111;
assign micromatrizz[40][347] = 9'b111111111;
assign micromatrizz[40][348] = 9'b111111111;
assign micromatrizz[40][349] = 9'b111111111;
assign micromatrizz[40][350] = 9'b111111111;
assign micromatrizz[40][351] = 9'b111111111;
assign micromatrizz[40][352] = 9'b111111111;
assign micromatrizz[40][353] = 9'b111111111;
assign micromatrizz[40][354] = 9'b111111111;
assign micromatrizz[40][355] = 9'b111111111;
assign micromatrizz[40][356] = 9'b111111111;
assign micromatrizz[40][357] = 9'b111111111;
assign micromatrizz[40][358] = 9'b111111111;
assign micromatrizz[40][359] = 9'b111111111;
assign micromatrizz[40][360] = 9'b111111111;
assign micromatrizz[40][361] = 9'b111111111;
assign micromatrizz[40][362] = 9'b111111111;
assign micromatrizz[40][363] = 9'b111111111;
assign micromatrizz[40][364] = 9'b111111111;
assign micromatrizz[40][365] = 9'b111111111;
assign micromatrizz[40][366] = 9'b111111111;
assign micromatrizz[40][367] = 9'b111111111;
assign micromatrizz[40][368] = 9'b111111111;
assign micromatrizz[40][369] = 9'b111111111;
assign micromatrizz[40][370] = 9'b111111111;
assign micromatrizz[40][371] = 9'b111111111;
assign micromatrizz[40][372] = 9'b111111111;
assign micromatrizz[40][373] = 9'b111111111;
assign micromatrizz[40][374] = 9'b111111111;
assign micromatrizz[40][375] = 9'b111111111;
assign micromatrizz[40][376] = 9'b111111111;
assign micromatrizz[40][377] = 9'b111111111;
assign micromatrizz[40][378] = 9'b111111111;
assign micromatrizz[40][379] = 9'b111111111;
assign micromatrizz[40][380] = 9'b111111111;
assign micromatrizz[40][381] = 9'b111111111;
assign micromatrizz[40][382] = 9'b111111111;
assign micromatrizz[40][383] = 9'b111111111;
assign micromatrizz[40][384] = 9'b111111111;
assign micromatrizz[40][385] = 9'b111111111;
assign micromatrizz[40][386] = 9'b111111111;
assign micromatrizz[40][387] = 9'b111111111;
assign micromatrizz[40][388] = 9'b111111111;
assign micromatrizz[40][389] = 9'b111111111;
assign micromatrizz[40][390] = 9'b111111111;
assign micromatrizz[40][391] = 9'b111111111;
assign micromatrizz[40][392] = 9'b111111111;
assign micromatrizz[40][393] = 9'b111111111;
assign micromatrizz[40][394] = 9'b111111111;
assign micromatrizz[40][395] = 9'b111111111;
assign micromatrizz[40][396] = 9'b111111111;
assign micromatrizz[40][397] = 9'b111111111;
assign micromatrizz[40][398] = 9'b111111111;
assign micromatrizz[40][399] = 9'b111111111;
assign micromatrizz[40][400] = 9'b111111111;
assign micromatrizz[40][401] = 9'b111111111;
assign micromatrizz[40][402] = 9'b111111111;
assign micromatrizz[40][403] = 9'b111111111;
assign micromatrizz[40][404] = 9'b111111111;
assign micromatrizz[40][405] = 9'b111111111;
assign micromatrizz[40][406] = 9'b111111111;
assign micromatrizz[40][407] = 9'b111111111;
assign micromatrizz[40][408] = 9'b111111111;
assign micromatrizz[40][409] = 9'b111111111;
assign micromatrizz[40][410] = 9'b111111111;
assign micromatrizz[40][411] = 9'b111111111;
assign micromatrizz[40][412] = 9'b111111111;
assign micromatrizz[40][413] = 9'b111111111;
assign micromatrizz[40][414] = 9'b111111111;
assign micromatrizz[40][415] = 9'b111111111;
assign micromatrizz[40][416] = 9'b111111111;
assign micromatrizz[40][417] = 9'b111111111;
assign micromatrizz[40][418] = 9'b111111111;
assign micromatrizz[40][419] = 9'b111111111;
assign micromatrizz[40][420] = 9'b111111111;
assign micromatrizz[40][421] = 9'b111111111;
assign micromatrizz[40][422] = 9'b111111111;
assign micromatrizz[40][423] = 9'b111111111;
assign micromatrizz[40][424] = 9'b111111111;
assign micromatrizz[40][425] = 9'b111111111;
assign micromatrizz[40][426] = 9'b111111111;
assign micromatrizz[40][427] = 9'b111111111;
assign micromatrizz[40][428] = 9'b111111111;
assign micromatrizz[40][429] = 9'b111111111;
assign micromatrizz[40][430] = 9'b111111111;
assign micromatrizz[40][431] = 9'b111111111;
assign micromatrizz[40][432] = 9'b111111111;
assign micromatrizz[40][433] = 9'b111111111;
assign micromatrizz[40][434] = 9'b111111111;
assign micromatrizz[40][435] = 9'b111111111;
assign micromatrizz[40][436] = 9'b111111111;
assign micromatrizz[40][437] = 9'b111111111;
assign micromatrizz[40][438] = 9'b111111111;
assign micromatrizz[40][439] = 9'b111111111;
assign micromatrizz[40][440] = 9'b111111111;
assign micromatrizz[40][441] = 9'b111111111;
assign micromatrizz[40][442] = 9'b111111111;
assign micromatrizz[40][443] = 9'b111111111;
assign micromatrizz[40][444] = 9'b111111111;
assign micromatrizz[40][445] = 9'b111111111;
assign micromatrizz[40][446] = 9'b111111111;
assign micromatrizz[40][447] = 9'b111111111;
assign micromatrizz[40][448] = 9'b111111111;
assign micromatrizz[40][449] = 9'b111111111;
assign micromatrizz[40][450] = 9'b111111111;
assign micromatrizz[40][451] = 9'b111111111;
assign micromatrizz[40][452] = 9'b111111111;
assign micromatrizz[40][453] = 9'b111111111;
assign micromatrizz[40][454] = 9'b111111111;
assign micromatrizz[40][455] = 9'b111111111;
assign micromatrizz[40][456] = 9'b111111111;
assign micromatrizz[40][457] = 9'b111111111;
assign micromatrizz[40][458] = 9'b111111111;
assign micromatrizz[40][459] = 9'b111111111;
assign micromatrizz[40][460] = 9'b111111111;
assign micromatrizz[40][461] = 9'b111111111;
assign micromatrizz[40][462] = 9'b111111111;
assign micromatrizz[40][463] = 9'b111111111;
assign micromatrizz[40][464] = 9'b111111111;
assign micromatrizz[40][465] = 9'b111111111;
assign micromatrizz[40][466] = 9'b111111111;
assign micromatrizz[40][467] = 9'b111111111;
assign micromatrizz[40][468] = 9'b111111111;
assign micromatrizz[40][469] = 9'b111111111;
assign micromatrizz[40][470] = 9'b111111111;
assign micromatrizz[40][471] = 9'b111111111;
assign micromatrizz[40][472] = 9'b111111111;
assign micromatrizz[40][473] = 9'b111111111;
assign micromatrizz[40][474] = 9'b111111111;
assign micromatrizz[40][475] = 9'b111111111;
assign micromatrizz[40][476] = 9'b111111111;
assign micromatrizz[40][477] = 9'b111111111;
assign micromatrizz[40][478] = 9'b111111111;
assign micromatrizz[40][479] = 9'b111111111;
assign micromatrizz[40][480] = 9'b111111111;
assign micromatrizz[40][481] = 9'b111111111;
assign micromatrizz[40][482] = 9'b111111111;
assign micromatrizz[40][483] = 9'b111111111;
assign micromatrizz[40][484] = 9'b111111111;
assign micromatrizz[40][485] = 9'b111111111;
assign micromatrizz[40][486] = 9'b111111111;
assign micromatrizz[40][487] = 9'b111111111;
assign micromatrizz[40][488] = 9'b111111111;
assign micromatrizz[40][489] = 9'b111111111;
assign micromatrizz[40][490] = 9'b111111111;
assign micromatrizz[40][491] = 9'b111111111;
assign micromatrizz[40][492] = 9'b111111111;
assign micromatrizz[40][493] = 9'b111111111;
assign micromatrizz[40][494] = 9'b111111111;
assign micromatrizz[40][495] = 9'b111111111;
assign micromatrizz[40][496] = 9'b111111111;
assign micromatrizz[40][497] = 9'b111111111;
assign micromatrizz[40][498] = 9'b111111111;
assign micromatrizz[40][499] = 9'b111111111;
assign micromatrizz[40][500] = 9'b111111111;
assign micromatrizz[40][501] = 9'b111111111;
assign micromatrizz[40][502] = 9'b111111111;
assign micromatrizz[40][503] = 9'b111111111;
assign micromatrizz[40][504] = 9'b111111111;
assign micromatrizz[40][505] = 9'b111111111;
assign micromatrizz[40][506] = 9'b111111111;
assign micromatrizz[40][507] = 9'b111111111;
assign micromatrizz[40][508] = 9'b111111111;
assign micromatrizz[40][509] = 9'b111111111;
assign micromatrizz[40][510] = 9'b111111111;
assign micromatrizz[40][511] = 9'b111111111;
assign micromatrizz[40][512] = 9'b111111111;
assign micromatrizz[40][513] = 9'b111111111;
assign micromatrizz[40][514] = 9'b111111111;
assign micromatrizz[40][515] = 9'b111111111;
assign micromatrizz[40][516] = 9'b111111111;
assign micromatrizz[40][517] = 9'b111111111;
assign micromatrizz[40][518] = 9'b111111111;
assign micromatrizz[40][519] = 9'b111111111;
assign micromatrizz[40][520] = 9'b111111111;
assign micromatrizz[40][521] = 9'b111111111;
assign micromatrizz[40][522] = 9'b111111111;
assign micromatrizz[40][523] = 9'b111111111;
assign micromatrizz[40][524] = 9'b111111111;
assign micromatrizz[40][525] = 9'b111111111;
assign micromatrizz[40][526] = 9'b111111111;
assign micromatrizz[40][527] = 9'b111111111;
assign micromatrizz[40][528] = 9'b111111111;
assign micromatrizz[40][529] = 9'b111111111;
assign micromatrizz[40][530] = 9'b111111111;
assign micromatrizz[40][531] = 9'b111111111;
assign micromatrizz[40][532] = 9'b111111111;
assign micromatrizz[40][533] = 9'b111111111;
assign micromatrizz[40][534] = 9'b111111111;
assign micromatrizz[40][535] = 9'b111111111;
assign micromatrizz[40][536] = 9'b111111111;
assign micromatrizz[40][537] = 9'b111111111;
assign micromatrizz[40][538] = 9'b111111111;
assign micromatrizz[40][539] = 9'b111111111;
assign micromatrizz[40][540] = 9'b111111111;
assign micromatrizz[40][541] = 9'b111111111;
assign micromatrizz[40][542] = 9'b111111111;
assign micromatrizz[40][543] = 9'b111111111;
assign micromatrizz[40][544] = 9'b111111111;
assign micromatrizz[40][545] = 9'b111111111;
assign micromatrizz[40][546] = 9'b111111111;
assign micromatrizz[40][547] = 9'b111111111;
assign micromatrizz[40][548] = 9'b111111111;
assign micromatrizz[40][549] = 9'b111111111;
assign micromatrizz[40][550] = 9'b111111111;
assign micromatrizz[40][551] = 9'b111111111;
assign micromatrizz[40][552] = 9'b111111111;
assign micromatrizz[40][553] = 9'b111111111;
assign micromatrizz[40][554] = 9'b111111111;
assign micromatrizz[40][555] = 9'b111111111;
assign micromatrizz[40][556] = 9'b111111111;
assign micromatrizz[40][557] = 9'b111111111;
assign micromatrizz[40][558] = 9'b111111111;
assign micromatrizz[40][559] = 9'b111111111;
assign micromatrizz[40][560] = 9'b111111111;
assign micromatrizz[40][561] = 9'b111111111;
assign micromatrizz[40][562] = 9'b111111111;
assign micromatrizz[40][563] = 9'b111111111;
assign micromatrizz[40][564] = 9'b111111111;
assign micromatrizz[40][565] = 9'b111111111;
assign micromatrizz[40][566] = 9'b111111111;
assign micromatrizz[40][567] = 9'b111111111;
assign micromatrizz[40][568] = 9'b111111111;
assign micromatrizz[40][569] = 9'b111111111;
assign micromatrizz[40][570] = 9'b111111111;
assign micromatrizz[40][571] = 9'b111111111;
assign micromatrizz[40][572] = 9'b111111111;
assign micromatrizz[40][573] = 9'b111111111;
assign micromatrizz[40][574] = 9'b111111111;
assign micromatrizz[40][575] = 9'b111111111;
assign micromatrizz[40][576] = 9'b111111111;
assign micromatrizz[40][577] = 9'b111111111;
assign micromatrizz[40][578] = 9'b111111111;
assign micromatrizz[40][579] = 9'b111111111;
assign micromatrizz[40][580] = 9'b111111111;
assign micromatrizz[40][581] = 9'b111111111;
assign micromatrizz[40][582] = 9'b111111111;
assign micromatrizz[40][583] = 9'b111111111;
assign micromatrizz[40][584] = 9'b111111111;
assign micromatrizz[40][585] = 9'b111111111;
assign micromatrizz[40][586] = 9'b111111111;
assign micromatrizz[40][587] = 9'b111111111;
assign micromatrizz[40][588] = 9'b111111111;
assign micromatrizz[40][589] = 9'b111111111;
assign micromatrizz[40][590] = 9'b111111111;
assign micromatrizz[40][591] = 9'b111111111;
assign micromatrizz[40][592] = 9'b111111111;
assign micromatrizz[40][593] = 9'b111111111;
assign micromatrizz[40][594] = 9'b111111111;
assign micromatrizz[40][595] = 9'b111111111;
assign micromatrizz[40][596] = 9'b111111111;
assign micromatrizz[40][597] = 9'b111111111;
assign micromatrizz[40][598] = 9'b111111111;
assign micromatrizz[40][599] = 9'b111111111;
assign micromatrizz[40][600] = 9'b111111111;
assign micromatrizz[40][601] = 9'b111111111;
assign micromatrizz[40][602] = 9'b111111111;
assign micromatrizz[40][603] = 9'b111111111;
assign micromatrizz[40][604] = 9'b111111111;
assign micromatrizz[40][605] = 9'b111111111;
assign micromatrizz[40][606] = 9'b111111111;
assign micromatrizz[40][607] = 9'b111111111;
assign micromatrizz[40][608] = 9'b111111111;
assign micromatrizz[40][609] = 9'b111111111;
assign micromatrizz[40][610] = 9'b111111111;
assign micromatrizz[40][611] = 9'b111111111;
assign micromatrizz[40][612] = 9'b111111111;
assign micromatrizz[40][613] = 9'b111111111;
assign micromatrizz[40][614] = 9'b111111111;
assign micromatrizz[40][615] = 9'b111111111;
assign micromatrizz[40][616] = 9'b111111111;
assign micromatrizz[40][617] = 9'b111111111;
assign micromatrizz[40][618] = 9'b111111111;
assign micromatrizz[40][619] = 9'b111111111;
assign micromatrizz[40][620] = 9'b111111111;
assign micromatrizz[40][621] = 9'b111111111;
assign micromatrizz[40][622] = 9'b111111111;
assign micromatrizz[40][623] = 9'b111111111;
assign micromatrizz[40][624] = 9'b111111111;
assign micromatrizz[40][625] = 9'b111111111;
assign micromatrizz[40][626] = 9'b111111111;
assign micromatrizz[40][627] = 9'b111111111;
assign micromatrizz[40][628] = 9'b111111111;
assign micromatrizz[40][629] = 9'b111111111;
assign micromatrizz[40][630] = 9'b111111111;
assign micromatrizz[40][631] = 9'b111111111;
assign micromatrizz[40][632] = 9'b111111111;
assign micromatrizz[40][633] = 9'b111111111;
assign micromatrizz[40][634] = 9'b111111111;
assign micromatrizz[40][635] = 9'b111111111;
assign micromatrizz[40][636] = 9'b111111111;
assign micromatrizz[40][637] = 9'b111111111;
assign micromatrizz[40][638] = 9'b111111111;
assign micromatrizz[40][639] = 9'b111111111;
assign micromatrizz[41][0] = 9'b111111111;
assign micromatrizz[41][1] = 9'b111111111;
assign micromatrizz[41][2] = 9'b111111111;
assign micromatrizz[41][3] = 9'b111111111;
assign micromatrizz[41][4] = 9'b111111111;
assign micromatrizz[41][5] = 9'b111111111;
assign micromatrizz[41][6] = 9'b111111111;
assign micromatrizz[41][7] = 9'b111111111;
assign micromatrizz[41][8] = 9'b111111111;
assign micromatrizz[41][9] = 9'b111111111;
assign micromatrizz[41][10] = 9'b111111111;
assign micromatrizz[41][11] = 9'b111111111;
assign micromatrizz[41][12] = 9'b111111111;
assign micromatrizz[41][13] = 9'b111111111;
assign micromatrizz[41][14] = 9'b111111111;
assign micromatrizz[41][15] = 9'b111111111;
assign micromatrizz[41][16] = 9'b111111111;
assign micromatrizz[41][17] = 9'b111111111;
assign micromatrizz[41][18] = 9'b111111111;
assign micromatrizz[41][19] = 9'b111111111;
assign micromatrizz[41][20] = 9'b111111111;
assign micromatrizz[41][21] = 9'b111111111;
assign micromatrizz[41][22] = 9'b111111111;
assign micromatrizz[41][23] = 9'b111111111;
assign micromatrizz[41][24] = 9'b111111111;
assign micromatrizz[41][25] = 9'b111111111;
assign micromatrizz[41][26] = 9'b111111111;
assign micromatrizz[41][27] = 9'b111111111;
assign micromatrizz[41][28] = 9'b111111111;
assign micromatrizz[41][29] = 9'b111111111;
assign micromatrizz[41][30] = 9'b111111111;
assign micromatrizz[41][31] = 9'b111111111;
assign micromatrizz[41][32] = 9'b111111111;
assign micromatrizz[41][33] = 9'b111111111;
assign micromatrizz[41][34] = 9'b111111111;
assign micromatrizz[41][35] = 9'b111111111;
assign micromatrizz[41][36] = 9'b111111111;
assign micromatrizz[41][37] = 9'b111111111;
assign micromatrizz[41][38] = 9'b111111111;
assign micromatrizz[41][39] = 9'b111111111;
assign micromatrizz[41][40] = 9'b111111111;
assign micromatrizz[41][41] = 9'b111111111;
assign micromatrizz[41][42] = 9'b111111111;
assign micromatrizz[41][43] = 9'b111111111;
assign micromatrizz[41][44] = 9'b111111111;
assign micromatrizz[41][45] = 9'b111111111;
assign micromatrizz[41][46] = 9'b111111111;
assign micromatrizz[41][47] = 9'b111111111;
assign micromatrizz[41][48] = 9'b111111111;
assign micromatrizz[41][49] = 9'b111111111;
assign micromatrizz[41][50] = 9'b111111111;
assign micromatrizz[41][51] = 9'b111111111;
assign micromatrizz[41][52] = 9'b111111111;
assign micromatrizz[41][53] = 9'b111111111;
assign micromatrizz[41][54] = 9'b111111111;
assign micromatrizz[41][55] = 9'b111111111;
assign micromatrizz[41][56] = 9'b111111111;
assign micromatrizz[41][57] = 9'b111111111;
assign micromatrizz[41][58] = 9'b111111111;
assign micromatrizz[41][59] = 9'b111111111;
assign micromatrizz[41][60] = 9'b111111111;
assign micromatrizz[41][61] = 9'b111111111;
assign micromatrizz[41][62] = 9'b111111111;
assign micromatrizz[41][63] = 9'b111111111;
assign micromatrizz[41][64] = 9'b111111111;
assign micromatrizz[41][65] = 9'b111111111;
assign micromatrizz[41][66] = 9'b111111111;
assign micromatrizz[41][67] = 9'b111111111;
assign micromatrizz[41][68] = 9'b111111111;
assign micromatrizz[41][69] = 9'b111111111;
assign micromatrizz[41][70] = 9'b111111111;
assign micromatrizz[41][71] = 9'b111111111;
assign micromatrizz[41][72] = 9'b111111111;
assign micromatrizz[41][73] = 9'b111111111;
assign micromatrizz[41][74] = 9'b111111111;
assign micromatrizz[41][75] = 9'b111111111;
assign micromatrizz[41][76] = 9'b111111111;
assign micromatrizz[41][77] = 9'b111111111;
assign micromatrizz[41][78] = 9'b111111111;
assign micromatrizz[41][79] = 9'b111111111;
assign micromatrizz[41][80] = 9'b111111111;
assign micromatrizz[41][81] = 9'b111111111;
assign micromatrizz[41][82] = 9'b111111111;
assign micromatrizz[41][83] = 9'b111111111;
assign micromatrizz[41][84] = 9'b111111111;
assign micromatrizz[41][85] = 9'b111111111;
assign micromatrizz[41][86] = 9'b111111111;
assign micromatrizz[41][87] = 9'b111111111;
assign micromatrizz[41][88] = 9'b111111111;
assign micromatrizz[41][89] = 9'b111111111;
assign micromatrizz[41][90] = 9'b111111111;
assign micromatrizz[41][91] = 9'b111111111;
assign micromatrizz[41][92] = 9'b111111111;
assign micromatrizz[41][93] = 9'b111111111;
assign micromatrizz[41][94] = 9'b111111111;
assign micromatrizz[41][95] = 9'b111111111;
assign micromatrizz[41][96] = 9'b111111111;
assign micromatrizz[41][97] = 9'b111111111;
assign micromatrizz[41][98] = 9'b111111111;
assign micromatrizz[41][99] = 9'b111111111;
assign micromatrizz[41][100] = 9'b111111111;
assign micromatrizz[41][101] = 9'b111111111;
assign micromatrizz[41][102] = 9'b111111111;
assign micromatrizz[41][103] = 9'b111111111;
assign micromatrizz[41][104] = 9'b111111111;
assign micromatrizz[41][105] = 9'b111111111;
assign micromatrizz[41][106] = 9'b111111111;
assign micromatrizz[41][107] = 9'b111111111;
assign micromatrizz[41][108] = 9'b111111111;
assign micromatrizz[41][109] = 9'b111111111;
assign micromatrizz[41][110] = 9'b111111111;
assign micromatrizz[41][111] = 9'b111111111;
assign micromatrizz[41][112] = 9'b111111111;
assign micromatrizz[41][113] = 9'b111111111;
assign micromatrizz[41][114] = 9'b111111111;
assign micromatrizz[41][115] = 9'b111111111;
assign micromatrizz[41][116] = 9'b111111111;
assign micromatrizz[41][117] = 9'b111111111;
assign micromatrizz[41][118] = 9'b111111111;
assign micromatrizz[41][119] = 9'b111111111;
assign micromatrizz[41][120] = 9'b111111111;
assign micromatrizz[41][121] = 9'b111111111;
assign micromatrizz[41][122] = 9'b111111111;
assign micromatrizz[41][123] = 9'b111111111;
assign micromatrizz[41][124] = 9'b111111111;
assign micromatrizz[41][125] = 9'b111111111;
assign micromatrizz[41][126] = 9'b111111111;
assign micromatrizz[41][127] = 9'b111111111;
assign micromatrizz[41][128] = 9'b111111111;
assign micromatrizz[41][129] = 9'b111111111;
assign micromatrizz[41][130] = 9'b111111111;
assign micromatrizz[41][131] = 9'b111111111;
assign micromatrizz[41][132] = 9'b111111111;
assign micromatrizz[41][133] = 9'b111111111;
assign micromatrizz[41][134] = 9'b111111111;
assign micromatrizz[41][135] = 9'b111111111;
assign micromatrizz[41][136] = 9'b111111111;
assign micromatrizz[41][137] = 9'b111111111;
assign micromatrizz[41][138] = 9'b111111111;
assign micromatrizz[41][139] = 9'b111111111;
assign micromatrizz[41][140] = 9'b111111111;
assign micromatrizz[41][141] = 9'b111111111;
assign micromatrizz[41][142] = 9'b111111111;
assign micromatrizz[41][143] = 9'b111111111;
assign micromatrizz[41][144] = 9'b111111111;
assign micromatrizz[41][145] = 9'b111111111;
assign micromatrizz[41][146] = 9'b111111111;
assign micromatrizz[41][147] = 9'b111111111;
assign micromatrizz[41][148] = 9'b111111111;
assign micromatrizz[41][149] = 9'b111111111;
assign micromatrizz[41][150] = 9'b111111111;
assign micromatrizz[41][151] = 9'b111111111;
assign micromatrizz[41][152] = 9'b111111111;
assign micromatrizz[41][153] = 9'b111111111;
assign micromatrizz[41][154] = 9'b111111111;
assign micromatrizz[41][155] = 9'b111111111;
assign micromatrizz[41][156] = 9'b111111111;
assign micromatrizz[41][157] = 9'b111111111;
assign micromatrizz[41][158] = 9'b111111111;
assign micromatrizz[41][159] = 9'b111111111;
assign micromatrizz[41][160] = 9'b111111111;
assign micromatrizz[41][161] = 9'b111111111;
assign micromatrizz[41][162] = 9'b111111111;
assign micromatrizz[41][163] = 9'b111111111;
assign micromatrizz[41][164] = 9'b111111111;
assign micromatrizz[41][165] = 9'b111111111;
assign micromatrizz[41][166] = 9'b111111111;
assign micromatrizz[41][167] = 9'b111111111;
assign micromatrizz[41][168] = 9'b111111111;
assign micromatrizz[41][169] = 9'b111111111;
assign micromatrizz[41][170] = 9'b111111111;
assign micromatrizz[41][171] = 9'b111111111;
assign micromatrizz[41][172] = 9'b111111111;
assign micromatrizz[41][173] = 9'b111111111;
assign micromatrizz[41][174] = 9'b111111111;
assign micromatrizz[41][175] = 9'b111111111;
assign micromatrizz[41][176] = 9'b111111111;
assign micromatrizz[41][177] = 9'b111111111;
assign micromatrizz[41][178] = 9'b111111111;
assign micromatrizz[41][179] = 9'b111111111;
assign micromatrizz[41][180] = 9'b111111111;
assign micromatrizz[41][181] = 9'b111111111;
assign micromatrizz[41][182] = 9'b111111111;
assign micromatrizz[41][183] = 9'b111111111;
assign micromatrizz[41][184] = 9'b111111111;
assign micromatrizz[41][185] = 9'b111111111;
assign micromatrizz[41][186] = 9'b111111111;
assign micromatrizz[41][187] = 9'b111111111;
assign micromatrizz[41][188] = 9'b111111111;
assign micromatrizz[41][189] = 9'b111111111;
assign micromatrizz[41][190] = 9'b111111111;
assign micromatrizz[41][191] = 9'b111111111;
assign micromatrizz[41][192] = 9'b111111111;
assign micromatrizz[41][193] = 9'b111111111;
assign micromatrizz[41][194] = 9'b111111111;
assign micromatrizz[41][195] = 9'b111111111;
assign micromatrizz[41][196] = 9'b111111111;
assign micromatrizz[41][197] = 9'b111111111;
assign micromatrizz[41][198] = 9'b111111111;
assign micromatrizz[41][199] = 9'b111111111;
assign micromatrizz[41][200] = 9'b111111111;
assign micromatrizz[41][201] = 9'b111111111;
assign micromatrizz[41][202] = 9'b111111111;
assign micromatrizz[41][203] = 9'b111111111;
assign micromatrizz[41][204] = 9'b111111111;
assign micromatrizz[41][205] = 9'b111111111;
assign micromatrizz[41][206] = 9'b111111111;
assign micromatrizz[41][207] = 9'b111111111;
assign micromatrizz[41][208] = 9'b111111111;
assign micromatrizz[41][209] = 9'b111111111;
assign micromatrizz[41][210] = 9'b111111111;
assign micromatrizz[41][211] = 9'b111111111;
assign micromatrizz[41][212] = 9'b111111111;
assign micromatrizz[41][213] = 9'b111111111;
assign micromatrizz[41][214] = 9'b111111111;
assign micromatrizz[41][215] = 9'b111111111;
assign micromatrizz[41][216] = 9'b111111111;
assign micromatrizz[41][217] = 9'b111111111;
assign micromatrizz[41][218] = 9'b111111111;
assign micromatrizz[41][219] = 9'b111111111;
assign micromatrizz[41][220] = 9'b111111111;
assign micromatrizz[41][221] = 9'b111111111;
assign micromatrizz[41][222] = 9'b111111111;
assign micromatrizz[41][223] = 9'b111111111;
assign micromatrizz[41][224] = 9'b111111111;
assign micromatrizz[41][225] = 9'b111111111;
assign micromatrizz[41][226] = 9'b111111111;
assign micromatrizz[41][227] = 9'b111111111;
assign micromatrizz[41][228] = 9'b111111111;
assign micromatrizz[41][229] = 9'b111111111;
assign micromatrizz[41][230] = 9'b111111111;
assign micromatrizz[41][231] = 9'b111111111;
assign micromatrizz[41][232] = 9'b111111111;
assign micromatrizz[41][233] = 9'b111111111;
assign micromatrizz[41][234] = 9'b111111111;
assign micromatrizz[41][235] = 9'b111111111;
assign micromatrizz[41][236] = 9'b111111111;
assign micromatrizz[41][237] = 9'b111111111;
assign micromatrizz[41][238] = 9'b111111111;
assign micromatrizz[41][239] = 9'b111111111;
assign micromatrizz[41][240] = 9'b111111111;
assign micromatrizz[41][241] = 9'b111111111;
assign micromatrizz[41][242] = 9'b111111111;
assign micromatrizz[41][243] = 9'b111111111;
assign micromatrizz[41][244] = 9'b111111111;
assign micromatrizz[41][245] = 9'b111111111;
assign micromatrizz[41][246] = 9'b111111111;
assign micromatrizz[41][247] = 9'b111111111;
assign micromatrizz[41][248] = 9'b111111111;
assign micromatrizz[41][249] = 9'b111111111;
assign micromatrizz[41][250] = 9'b111111111;
assign micromatrizz[41][251] = 9'b111111111;
assign micromatrizz[41][252] = 9'b111111111;
assign micromatrizz[41][253] = 9'b111111111;
assign micromatrizz[41][254] = 9'b111111111;
assign micromatrizz[41][255] = 9'b111111111;
assign micromatrizz[41][256] = 9'b111111111;
assign micromatrizz[41][257] = 9'b111111111;
assign micromatrizz[41][258] = 9'b111111111;
assign micromatrizz[41][259] = 9'b111111111;
assign micromatrizz[41][260] = 9'b111111111;
assign micromatrizz[41][261] = 9'b111111111;
assign micromatrizz[41][262] = 9'b111111111;
assign micromatrizz[41][263] = 9'b111111111;
assign micromatrizz[41][264] = 9'b111111111;
assign micromatrizz[41][265] = 9'b111111111;
assign micromatrizz[41][266] = 9'b111111111;
assign micromatrizz[41][267] = 9'b111111111;
assign micromatrizz[41][268] = 9'b111111111;
assign micromatrizz[41][269] = 9'b111111111;
assign micromatrizz[41][270] = 9'b111111111;
assign micromatrizz[41][271] = 9'b111111111;
assign micromatrizz[41][272] = 9'b111111111;
assign micromatrizz[41][273] = 9'b111111111;
assign micromatrizz[41][274] = 9'b111111111;
assign micromatrizz[41][275] = 9'b111111111;
assign micromatrizz[41][276] = 9'b111111111;
assign micromatrizz[41][277] = 9'b111111111;
assign micromatrizz[41][278] = 9'b111111111;
assign micromatrizz[41][279] = 9'b111111111;
assign micromatrizz[41][280] = 9'b111111111;
assign micromatrizz[41][281] = 9'b111111111;
assign micromatrizz[41][282] = 9'b111111111;
assign micromatrizz[41][283] = 9'b111111111;
assign micromatrizz[41][284] = 9'b111111111;
assign micromatrizz[41][285] = 9'b111111111;
assign micromatrizz[41][286] = 9'b111111111;
assign micromatrizz[41][287] = 9'b111111111;
assign micromatrizz[41][288] = 9'b111111111;
assign micromatrizz[41][289] = 9'b111111111;
assign micromatrizz[41][290] = 9'b111111111;
assign micromatrizz[41][291] = 9'b111111111;
assign micromatrizz[41][292] = 9'b111111111;
assign micromatrizz[41][293] = 9'b111111111;
assign micromatrizz[41][294] = 9'b111111111;
assign micromatrizz[41][295] = 9'b111111111;
assign micromatrizz[41][296] = 9'b111111111;
assign micromatrizz[41][297] = 9'b111111111;
assign micromatrizz[41][298] = 9'b111111111;
assign micromatrizz[41][299] = 9'b111111111;
assign micromatrizz[41][300] = 9'b111111111;
assign micromatrizz[41][301] = 9'b111111111;
assign micromatrizz[41][302] = 9'b111111111;
assign micromatrizz[41][303] = 9'b111111111;
assign micromatrizz[41][304] = 9'b111111111;
assign micromatrizz[41][305] = 9'b111111111;
assign micromatrizz[41][306] = 9'b111111111;
assign micromatrizz[41][307] = 9'b111111111;
assign micromatrizz[41][308] = 9'b111111111;
assign micromatrizz[41][309] = 9'b111111111;
assign micromatrizz[41][310] = 9'b111111111;
assign micromatrizz[41][311] = 9'b111111111;
assign micromatrizz[41][312] = 9'b111111111;
assign micromatrizz[41][313] = 9'b111111111;
assign micromatrizz[41][314] = 9'b111111111;
assign micromatrizz[41][315] = 9'b111111111;
assign micromatrizz[41][316] = 9'b111111111;
assign micromatrizz[41][317] = 9'b111111111;
assign micromatrizz[41][318] = 9'b111111111;
assign micromatrizz[41][319] = 9'b111111111;
assign micromatrizz[41][320] = 9'b111111111;
assign micromatrizz[41][321] = 9'b111111111;
assign micromatrizz[41][322] = 9'b111111111;
assign micromatrizz[41][323] = 9'b111111111;
assign micromatrizz[41][324] = 9'b111111111;
assign micromatrizz[41][325] = 9'b111111111;
assign micromatrizz[41][326] = 9'b111111111;
assign micromatrizz[41][327] = 9'b111111111;
assign micromatrizz[41][328] = 9'b111111111;
assign micromatrizz[41][329] = 9'b111111111;
assign micromatrizz[41][330] = 9'b111111111;
assign micromatrizz[41][331] = 9'b111111111;
assign micromatrizz[41][332] = 9'b111111111;
assign micromatrizz[41][333] = 9'b111111111;
assign micromatrizz[41][334] = 9'b111111111;
assign micromatrizz[41][335] = 9'b111111111;
assign micromatrizz[41][336] = 9'b111111111;
assign micromatrizz[41][337] = 9'b111111111;
assign micromatrizz[41][338] = 9'b111111111;
assign micromatrizz[41][339] = 9'b111111111;
assign micromatrizz[41][340] = 9'b111111111;
assign micromatrizz[41][341] = 9'b111111111;
assign micromatrizz[41][342] = 9'b111111111;
assign micromatrizz[41][343] = 9'b111111111;
assign micromatrizz[41][344] = 9'b111111111;
assign micromatrizz[41][345] = 9'b111111111;
assign micromatrizz[41][346] = 9'b111111111;
assign micromatrizz[41][347] = 9'b111111111;
assign micromatrizz[41][348] = 9'b111111111;
assign micromatrizz[41][349] = 9'b111111111;
assign micromatrizz[41][350] = 9'b111111111;
assign micromatrizz[41][351] = 9'b111111111;
assign micromatrizz[41][352] = 9'b111111111;
assign micromatrizz[41][353] = 9'b111111111;
assign micromatrizz[41][354] = 9'b111111111;
assign micromatrizz[41][355] = 9'b111111111;
assign micromatrizz[41][356] = 9'b111111111;
assign micromatrizz[41][357] = 9'b111111111;
assign micromatrizz[41][358] = 9'b111111111;
assign micromatrizz[41][359] = 9'b111111111;
assign micromatrizz[41][360] = 9'b111111111;
assign micromatrizz[41][361] = 9'b111111111;
assign micromatrizz[41][362] = 9'b111111111;
assign micromatrizz[41][363] = 9'b111111111;
assign micromatrizz[41][364] = 9'b111111111;
assign micromatrizz[41][365] = 9'b111111111;
assign micromatrizz[41][366] = 9'b111111111;
assign micromatrizz[41][367] = 9'b111111111;
assign micromatrizz[41][368] = 9'b111111111;
assign micromatrizz[41][369] = 9'b111111111;
assign micromatrizz[41][370] = 9'b111111111;
assign micromatrizz[41][371] = 9'b111111111;
assign micromatrizz[41][372] = 9'b111111111;
assign micromatrizz[41][373] = 9'b111111111;
assign micromatrizz[41][374] = 9'b111111111;
assign micromatrizz[41][375] = 9'b111111111;
assign micromatrizz[41][376] = 9'b111111111;
assign micromatrizz[41][377] = 9'b111111111;
assign micromatrizz[41][378] = 9'b111111111;
assign micromatrizz[41][379] = 9'b111111111;
assign micromatrizz[41][380] = 9'b111111111;
assign micromatrizz[41][381] = 9'b111111111;
assign micromatrizz[41][382] = 9'b111111111;
assign micromatrizz[41][383] = 9'b111111111;
assign micromatrizz[41][384] = 9'b111111111;
assign micromatrizz[41][385] = 9'b111111111;
assign micromatrizz[41][386] = 9'b111111111;
assign micromatrizz[41][387] = 9'b111111111;
assign micromatrizz[41][388] = 9'b111111111;
assign micromatrizz[41][389] = 9'b111111111;
assign micromatrizz[41][390] = 9'b111111111;
assign micromatrizz[41][391] = 9'b111111111;
assign micromatrizz[41][392] = 9'b111111111;
assign micromatrizz[41][393] = 9'b111111111;
assign micromatrizz[41][394] = 9'b111111111;
assign micromatrizz[41][395] = 9'b111111111;
assign micromatrizz[41][396] = 9'b111111111;
assign micromatrizz[41][397] = 9'b111111111;
assign micromatrizz[41][398] = 9'b111111111;
assign micromatrizz[41][399] = 9'b111111111;
assign micromatrizz[41][400] = 9'b111111111;
assign micromatrizz[41][401] = 9'b111111111;
assign micromatrizz[41][402] = 9'b111111111;
assign micromatrizz[41][403] = 9'b111111111;
assign micromatrizz[41][404] = 9'b111111111;
assign micromatrizz[41][405] = 9'b111111111;
assign micromatrizz[41][406] = 9'b111111111;
assign micromatrizz[41][407] = 9'b111111111;
assign micromatrizz[41][408] = 9'b111111111;
assign micromatrizz[41][409] = 9'b111111111;
assign micromatrizz[41][410] = 9'b111111111;
assign micromatrizz[41][411] = 9'b111111111;
assign micromatrizz[41][412] = 9'b111111111;
assign micromatrizz[41][413] = 9'b111111111;
assign micromatrizz[41][414] = 9'b111111111;
assign micromatrizz[41][415] = 9'b111111111;
assign micromatrizz[41][416] = 9'b111111111;
assign micromatrizz[41][417] = 9'b111111111;
assign micromatrizz[41][418] = 9'b111111111;
assign micromatrizz[41][419] = 9'b111111111;
assign micromatrizz[41][420] = 9'b111111111;
assign micromatrizz[41][421] = 9'b111111111;
assign micromatrizz[41][422] = 9'b111111111;
assign micromatrizz[41][423] = 9'b111111111;
assign micromatrizz[41][424] = 9'b111111111;
assign micromatrizz[41][425] = 9'b111111111;
assign micromatrizz[41][426] = 9'b111111111;
assign micromatrizz[41][427] = 9'b111111111;
assign micromatrizz[41][428] = 9'b111111111;
assign micromatrizz[41][429] = 9'b111111111;
assign micromatrizz[41][430] = 9'b111111111;
assign micromatrizz[41][431] = 9'b111111111;
assign micromatrizz[41][432] = 9'b111111111;
assign micromatrizz[41][433] = 9'b111111111;
assign micromatrizz[41][434] = 9'b111111111;
assign micromatrizz[41][435] = 9'b111111111;
assign micromatrizz[41][436] = 9'b111111111;
assign micromatrizz[41][437] = 9'b111111111;
assign micromatrizz[41][438] = 9'b111111111;
assign micromatrizz[41][439] = 9'b111111111;
assign micromatrizz[41][440] = 9'b111111111;
assign micromatrizz[41][441] = 9'b111111111;
assign micromatrizz[41][442] = 9'b111111111;
assign micromatrizz[41][443] = 9'b111111111;
assign micromatrizz[41][444] = 9'b111111111;
assign micromatrizz[41][445] = 9'b111111111;
assign micromatrizz[41][446] = 9'b111111111;
assign micromatrizz[41][447] = 9'b111111111;
assign micromatrizz[41][448] = 9'b111111111;
assign micromatrizz[41][449] = 9'b111111111;
assign micromatrizz[41][450] = 9'b111111111;
assign micromatrizz[41][451] = 9'b111111111;
assign micromatrizz[41][452] = 9'b111111111;
assign micromatrizz[41][453] = 9'b111111111;
assign micromatrizz[41][454] = 9'b111111111;
assign micromatrizz[41][455] = 9'b111111111;
assign micromatrizz[41][456] = 9'b111111111;
assign micromatrizz[41][457] = 9'b111111111;
assign micromatrizz[41][458] = 9'b111111111;
assign micromatrizz[41][459] = 9'b111111111;
assign micromatrizz[41][460] = 9'b111111111;
assign micromatrizz[41][461] = 9'b111111111;
assign micromatrizz[41][462] = 9'b111111111;
assign micromatrizz[41][463] = 9'b111111111;
assign micromatrizz[41][464] = 9'b111111111;
assign micromatrizz[41][465] = 9'b111111111;
assign micromatrizz[41][466] = 9'b111111111;
assign micromatrizz[41][467] = 9'b111111111;
assign micromatrizz[41][468] = 9'b111111111;
assign micromatrizz[41][469] = 9'b111111111;
assign micromatrizz[41][470] = 9'b111111111;
assign micromatrizz[41][471] = 9'b111111111;
assign micromatrizz[41][472] = 9'b111111111;
assign micromatrizz[41][473] = 9'b111111111;
assign micromatrizz[41][474] = 9'b111111111;
assign micromatrizz[41][475] = 9'b111111111;
assign micromatrizz[41][476] = 9'b111111111;
assign micromatrizz[41][477] = 9'b111111111;
assign micromatrizz[41][478] = 9'b111111111;
assign micromatrizz[41][479] = 9'b111111111;
assign micromatrizz[41][480] = 9'b111111111;
assign micromatrizz[41][481] = 9'b111111111;
assign micromatrizz[41][482] = 9'b111111111;
assign micromatrizz[41][483] = 9'b111111111;
assign micromatrizz[41][484] = 9'b111111111;
assign micromatrizz[41][485] = 9'b111111111;
assign micromatrizz[41][486] = 9'b111111111;
assign micromatrizz[41][487] = 9'b111111111;
assign micromatrizz[41][488] = 9'b111111111;
assign micromatrizz[41][489] = 9'b111111111;
assign micromatrizz[41][490] = 9'b111111111;
assign micromatrizz[41][491] = 9'b111111111;
assign micromatrizz[41][492] = 9'b111111111;
assign micromatrizz[41][493] = 9'b111111111;
assign micromatrizz[41][494] = 9'b111111111;
assign micromatrizz[41][495] = 9'b111111111;
assign micromatrizz[41][496] = 9'b111111111;
assign micromatrizz[41][497] = 9'b111111111;
assign micromatrizz[41][498] = 9'b111111111;
assign micromatrizz[41][499] = 9'b111111111;
assign micromatrizz[41][500] = 9'b111111111;
assign micromatrizz[41][501] = 9'b111111111;
assign micromatrizz[41][502] = 9'b111111111;
assign micromatrizz[41][503] = 9'b111111111;
assign micromatrizz[41][504] = 9'b111111111;
assign micromatrizz[41][505] = 9'b111111111;
assign micromatrizz[41][506] = 9'b111111111;
assign micromatrizz[41][507] = 9'b111111111;
assign micromatrizz[41][508] = 9'b111111111;
assign micromatrizz[41][509] = 9'b111111111;
assign micromatrizz[41][510] = 9'b111111111;
assign micromatrizz[41][511] = 9'b111111111;
assign micromatrizz[41][512] = 9'b111111111;
assign micromatrizz[41][513] = 9'b111111111;
assign micromatrizz[41][514] = 9'b111111111;
assign micromatrizz[41][515] = 9'b111111111;
assign micromatrizz[41][516] = 9'b111111111;
assign micromatrizz[41][517] = 9'b111111111;
assign micromatrizz[41][518] = 9'b111111111;
assign micromatrizz[41][519] = 9'b111111111;
assign micromatrizz[41][520] = 9'b111111111;
assign micromatrizz[41][521] = 9'b111111111;
assign micromatrizz[41][522] = 9'b111111111;
assign micromatrizz[41][523] = 9'b111111111;
assign micromatrizz[41][524] = 9'b111111111;
assign micromatrizz[41][525] = 9'b111111111;
assign micromatrizz[41][526] = 9'b111111111;
assign micromatrizz[41][527] = 9'b111111111;
assign micromatrizz[41][528] = 9'b111111111;
assign micromatrizz[41][529] = 9'b111111111;
assign micromatrizz[41][530] = 9'b111111111;
assign micromatrizz[41][531] = 9'b111111111;
assign micromatrizz[41][532] = 9'b111111111;
assign micromatrizz[41][533] = 9'b111111111;
assign micromatrizz[41][534] = 9'b111111111;
assign micromatrizz[41][535] = 9'b111111111;
assign micromatrizz[41][536] = 9'b111111111;
assign micromatrizz[41][537] = 9'b111111111;
assign micromatrizz[41][538] = 9'b111111111;
assign micromatrizz[41][539] = 9'b111111111;
assign micromatrizz[41][540] = 9'b111111111;
assign micromatrizz[41][541] = 9'b111111111;
assign micromatrizz[41][542] = 9'b111111111;
assign micromatrizz[41][543] = 9'b111111111;
assign micromatrizz[41][544] = 9'b111111111;
assign micromatrizz[41][545] = 9'b111111111;
assign micromatrizz[41][546] = 9'b111111111;
assign micromatrizz[41][547] = 9'b111111111;
assign micromatrizz[41][548] = 9'b111111111;
assign micromatrizz[41][549] = 9'b111111111;
assign micromatrizz[41][550] = 9'b111111111;
assign micromatrizz[41][551] = 9'b111111111;
assign micromatrizz[41][552] = 9'b111111111;
assign micromatrizz[41][553] = 9'b111111111;
assign micromatrizz[41][554] = 9'b111111111;
assign micromatrizz[41][555] = 9'b111111111;
assign micromatrizz[41][556] = 9'b111111111;
assign micromatrizz[41][557] = 9'b111111111;
assign micromatrizz[41][558] = 9'b111111111;
assign micromatrizz[41][559] = 9'b111111111;
assign micromatrizz[41][560] = 9'b111111111;
assign micromatrizz[41][561] = 9'b111111111;
assign micromatrizz[41][562] = 9'b111111111;
assign micromatrizz[41][563] = 9'b111111111;
assign micromatrizz[41][564] = 9'b111111111;
assign micromatrizz[41][565] = 9'b111111111;
assign micromatrizz[41][566] = 9'b111111111;
assign micromatrizz[41][567] = 9'b111111111;
assign micromatrizz[41][568] = 9'b111111111;
assign micromatrizz[41][569] = 9'b111111111;
assign micromatrizz[41][570] = 9'b111111111;
assign micromatrizz[41][571] = 9'b111111111;
assign micromatrizz[41][572] = 9'b111111111;
assign micromatrizz[41][573] = 9'b111111111;
assign micromatrizz[41][574] = 9'b111111111;
assign micromatrizz[41][575] = 9'b111111111;
assign micromatrizz[41][576] = 9'b111111111;
assign micromatrizz[41][577] = 9'b111111111;
assign micromatrizz[41][578] = 9'b111111111;
assign micromatrizz[41][579] = 9'b111111111;
assign micromatrizz[41][580] = 9'b111111111;
assign micromatrizz[41][581] = 9'b111111111;
assign micromatrizz[41][582] = 9'b111111111;
assign micromatrizz[41][583] = 9'b111111111;
assign micromatrizz[41][584] = 9'b111111111;
assign micromatrizz[41][585] = 9'b111111111;
assign micromatrizz[41][586] = 9'b111111111;
assign micromatrizz[41][587] = 9'b111111111;
assign micromatrizz[41][588] = 9'b111111111;
assign micromatrizz[41][589] = 9'b111111111;
assign micromatrizz[41][590] = 9'b111111111;
assign micromatrizz[41][591] = 9'b111111111;
assign micromatrizz[41][592] = 9'b111111111;
assign micromatrizz[41][593] = 9'b111111111;
assign micromatrizz[41][594] = 9'b111111111;
assign micromatrizz[41][595] = 9'b111111111;
assign micromatrizz[41][596] = 9'b111111111;
assign micromatrizz[41][597] = 9'b111111111;
assign micromatrizz[41][598] = 9'b111111111;
assign micromatrizz[41][599] = 9'b111111111;
assign micromatrizz[41][600] = 9'b111111111;
assign micromatrizz[41][601] = 9'b111111111;
assign micromatrizz[41][602] = 9'b111111111;
assign micromatrizz[41][603] = 9'b111111111;
assign micromatrizz[41][604] = 9'b111111111;
assign micromatrizz[41][605] = 9'b111111111;
assign micromatrizz[41][606] = 9'b111111111;
assign micromatrizz[41][607] = 9'b111111111;
assign micromatrizz[41][608] = 9'b111111111;
assign micromatrizz[41][609] = 9'b111111111;
assign micromatrizz[41][610] = 9'b111111111;
assign micromatrizz[41][611] = 9'b111111111;
assign micromatrizz[41][612] = 9'b111111111;
assign micromatrizz[41][613] = 9'b111111111;
assign micromatrizz[41][614] = 9'b111111111;
assign micromatrizz[41][615] = 9'b111111111;
assign micromatrizz[41][616] = 9'b111111111;
assign micromatrizz[41][617] = 9'b111111111;
assign micromatrizz[41][618] = 9'b111111111;
assign micromatrizz[41][619] = 9'b111111111;
assign micromatrizz[41][620] = 9'b111111111;
assign micromatrizz[41][621] = 9'b111111111;
assign micromatrizz[41][622] = 9'b111111111;
assign micromatrizz[41][623] = 9'b111111111;
assign micromatrizz[41][624] = 9'b111111111;
assign micromatrizz[41][625] = 9'b111111111;
assign micromatrizz[41][626] = 9'b111111111;
assign micromatrizz[41][627] = 9'b111111111;
assign micromatrizz[41][628] = 9'b111111111;
assign micromatrizz[41][629] = 9'b111111111;
assign micromatrizz[41][630] = 9'b111111111;
assign micromatrizz[41][631] = 9'b111111111;
assign micromatrizz[41][632] = 9'b111111111;
assign micromatrizz[41][633] = 9'b111111111;
assign micromatrizz[41][634] = 9'b111111111;
assign micromatrizz[41][635] = 9'b111111111;
assign micromatrizz[41][636] = 9'b111111111;
assign micromatrizz[41][637] = 9'b111111111;
assign micromatrizz[41][638] = 9'b111111111;
assign micromatrizz[41][639] = 9'b111111111;
assign micromatrizz[42][0] = 9'b111111111;
assign micromatrizz[42][1] = 9'b111111111;
assign micromatrizz[42][2] = 9'b111111111;
assign micromatrizz[42][3] = 9'b111111111;
assign micromatrizz[42][4] = 9'b111111111;
assign micromatrizz[42][5] = 9'b111111111;
assign micromatrizz[42][6] = 9'b111111111;
assign micromatrizz[42][7] = 9'b111111111;
assign micromatrizz[42][8] = 9'b111111111;
assign micromatrizz[42][9] = 9'b111111111;
assign micromatrizz[42][10] = 9'b111111111;
assign micromatrizz[42][11] = 9'b111111111;
assign micromatrizz[42][12] = 9'b111111111;
assign micromatrizz[42][13] = 9'b111111111;
assign micromatrizz[42][14] = 9'b111111111;
assign micromatrizz[42][15] = 9'b111111111;
assign micromatrizz[42][16] = 9'b111111111;
assign micromatrizz[42][17] = 9'b111111111;
assign micromatrizz[42][18] = 9'b111111111;
assign micromatrizz[42][19] = 9'b111111111;
assign micromatrizz[42][20] = 9'b111111111;
assign micromatrizz[42][21] = 9'b111111111;
assign micromatrizz[42][22] = 9'b111111111;
assign micromatrizz[42][23] = 9'b111111111;
assign micromatrizz[42][24] = 9'b111111111;
assign micromatrizz[42][25] = 9'b111111111;
assign micromatrizz[42][26] = 9'b111111111;
assign micromatrizz[42][27] = 9'b111111111;
assign micromatrizz[42][28] = 9'b111111111;
assign micromatrizz[42][29] = 9'b111111111;
assign micromatrizz[42][30] = 9'b111111111;
assign micromatrizz[42][31] = 9'b111111111;
assign micromatrizz[42][32] = 9'b111111111;
assign micromatrizz[42][33] = 9'b111111111;
assign micromatrizz[42][34] = 9'b111111111;
assign micromatrizz[42][35] = 9'b111111111;
assign micromatrizz[42][36] = 9'b111111111;
assign micromatrizz[42][37] = 9'b111111111;
assign micromatrizz[42][38] = 9'b111111111;
assign micromatrizz[42][39] = 9'b111111111;
assign micromatrizz[42][40] = 9'b111111111;
assign micromatrizz[42][41] = 9'b111111111;
assign micromatrizz[42][42] = 9'b111111111;
assign micromatrizz[42][43] = 9'b111111111;
assign micromatrizz[42][44] = 9'b111111111;
assign micromatrizz[42][45] = 9'b111111111;
assign micromatrizz[42][46] = 9'b111111111;
assign micromatrizz[42][47] = 9'b111111111;
assign micromatrizz[42][48] = 9'b111111111;
assign micromatrizz[42][49] = 9'b111111111;
assign micromatrizz[42][50] = 9'b111111111;
assign micromatrizz[42][51] = 9'b111111111;
assign micromatrizz[42][52] = 9'b111111111;
assign micromatrizz[42][53] = 9'b111111111;
assign micromatrizz[42][54] = 9'b111111111;
assign micromatrizz[42][55] = 9'b111111111;
assign micromatrizz[42][56] = 9'b111111111;
assign micromatrizz[42][57] = 9'b111111111;
assign micromatrizz[42][58] = 9'b111111111;
assign micromatrizz[42][59] = 9'b111111111;
assign micromatrizz[42][60] = 9'b111111111;
assign micromatrizz[42][61] = 9'b111111111;
assign micromatrizz[42][62] = 9'b111111111;
assign micromatrizz[42][63] = 9'b111111111;
assign micromatrizz[42][64] = 9'b111111111;
assign micromatrizz[42][65] = 9'b111111111;
assign micromatrizz[42][66] = 9'b111111111;
assign micromatrizz[42][67] = 9'b111111111;
assign micromatrizz[42][68] = 9'b111111111;
assign micromatrizz[42][69] = 9'b111111111;
assign micromatrizz[42][70] = 9'b111111111;
assign micromatrizz[42][71] = 9'b111111111;
assign micromatrizz[42][72] = 9'b111111111;
assign micromatrizz[42][73] = 9'b111111111;
assign micromatrizz[42][74] = 9'b111111111;
assign micromatrizz[42][75] = 9'b111111111;
assign micromatrizz[42][76] = 9'b111111111;
assign micromatrizz[42][77] = 9'b111111111;
assign micromatrizz[42][78] = 9'b111111111;
assign micromatrizz[42][79] = 9'b111111111;
assign micromatrizz[42][80] = 9'b111111111;
assign micromatrizz[42][81] = 9'b111111111;
assign micromatrizz[42][82] = 9'b111111111;
assign micromatrizz[42][83] = 9'b111111111;
assign micromatrizz[42][84] = 9'b111111111;
assign micromatrizz[42][85] = 9'b111111111;
assign micromatrizz[42][86] = 9'b111111111;
assign micromatrizz[42][87] = 9'b111111111;
assign micromatrizz[42][88] = 9'b111111111;
assign micromatrizz[42][89] = 9'b111111111;
assign micromatrizz[42][90] = 9'b111111111;
assign micromatrizz[42][91] = 9'b111111111;
assign micromatrizz[42][92] = 9'b111111111;
assign micromatrizz[42][93] = 9'b111111111;
assign micromatrizz[42][94] = 9'b111111111;
assign micromatrizz[42][95] = 9'b111111111;
assign micromatrizz[42][96] = 9'b111111111;
assign micromatrizz[42][97] = 9'b111111111;
assign micromatrizz[42][98] = 9'b111111111;
assign micromatrizz[42][99] = 9'b111111111;
assign micromatrizz[42][100] = 9'b111111111;
assign micromatrizz[42][101] = 9'b111111111;
assign micromatrizz[42][102] = 9'b111111111;
assign micromatrizz[42][103] = 9'b111111111;
assign micromatrizz[42][104] = 9'b111111111;
assign micromatrizz[42][105] = 9'b111111111;
assign micromatrizz[42][106] = 9'b111111111;
assign micromatrizz[42][107] = 9'b111111111;
assign micromatrizz[42][108] = 9'b111111111;
assign micromatrizz[42][109] = 9'b111111111;
assign micromatrizz[42][110] = 9'b111111111;
assign micromatrizz[42][111] = 9'b111111111;
assign micromatrizz[42][112] = 9'b111111111;
assign micromatrizz[42][113] = 9'b111111111;
assign micromatrizz[42][114] = 9'b111111111;
assign micromatrizz[42][115] = 9'b111111111;
assign micromatrizz[42][116] = 9'b111111111;
assign micromatrizz[42][117] = 9'b111111111;
assign micromatrizz[42][118] = 9'b111111111;
assign micromatrizz[42][119] = 9'b111111111;
assign micromatrizz[42][120] = 9'b111111111;
assign micromatrizz[42][121] = 9'b111111111;
assign micromatrizz[42][122] = 9'b111111111;
assign micromatrizz[42][123] = 9'b111111111;
assign micromatrizz[42][124] = 9'b111111111;
assign micromatrizz[42][125] = 9'b111111111;
assign micromatrizz[42][126] = 9'b111111111;
assign micromatrizz[42][127] = 9'b111111111;
assign micromatrizz[42][128] = 9'b111111111;
assign micromatrizz[42][129] = 9'b111111111;
assign micromatrizz[42][130] = 9'b111111111;
assign micromatrizz[42][131] = 9'b111111111;
assign micromatrizz[42][132] = 9'b111111111;
assign micromatrizz[42][133] = 9'b111111111;
assign micromatrizz[42][134] = 9'b111111111;
assign micromatrizz[42][135] = 9'b111111111;
assign micromatrizz[42][136] = 9'b111111111;
assign micromatrizz[42][137] = 9'b111111111;
assign micromatrizz[42][138] = 9'b111111111;
assign micromatrizz[42][139] = 9'b111111111;
assign micromatrizz[42][140] = 9'b111111111;
assign micromatrizz[42][141] = 9'b111111111;
assign micromatrizz[42][142] = 9'b111111111;
assign micromatrizz[42][143] = 9'b111111111;
assign micromatrizz[42][144] = 9'b111111111;
assign micromatrizz[42][145] = 9'b111111111;
assign micromatrizz[42][146] = 9'b111111111;
assign micromatrizz[42][147] = 9'b111111111;
assign micromatrizz[42][148] = 9'b111111111;
assign micromatrizz[42][149] = 9'b111111111;
assign micromatrizz[42][150] = 9'b111111111;
assign micromatrizz[42][151] = 9'b111111111;
assign micromatrizz[42][152] = 9'b111111111;
assign micromatrizz[42][153] = 9'b111111111;
assign micromatrizz[42][154] = 9'b111111111;
assign micromatrizz[42][155] = 9'b111111111;
assign micromatrizz[42][156] = 9'b111111111;
assign micromatrizz[42][157] = 9'b111111111;
assign micromatrizz[42][158] = 9'b111111111;
assign micromatrizz[42][159] = 9'b111111111;
assign micromatrizz[42][160] = 9'b111111111;
assign micromatrizz[42][161] = 9'b111111111;
assign micromatrizz[42][162] = 9'b111111111;
assign micromatrizz[42][163] = 9'b111111111;
assign micromatrizz[42][164] = 9'b111111111;
assign micromatrizz[42][165] = 9'b111111111;
assign micromatrizz[42][166] = 9'b111111111;
assign micromatrizz[42][167] = 9'b111111111;
assign micromatrizz[42][168] = 9'b111111111;
assign micromatrizz[42][169] = 9'b111111111;
assign micromatrizz[42][170] = 9'b111111111;
assign micromatrizz[42][171] = 9'b111111111;
assign micromatrizz[42][172] = 9'b111111111;
assign micromatrizz[42][173] = 9'b111111111;
assign micromatrizz[42][174] = 9'b111111111;
assign micromatrizz[42][175] = 9'b111111111;
assign micromatrizz[42][176] = 9'b111111111;
assign micromatrizz[42][177] = 9'b111111111;
assign micromatrizz[42][178] = 9'b111111111;
assign micromatrizz[42][179] = 9'b111111111;
assign micromatrizz[42][180] = 9'b111111111;
assign micromatrizz[42][181] = 9'b111111111;
assign micromatrizz[42][182] = 9'b111111111;
assign micromatrizz[42][183] = 9'b111111111;
assign micromatrizz[42][184] = 9'b111111111;
assign micromatrizz[42][185] = 9'b111111111;
assign micromatrizz[42][186] = 9'b111111111;
assign micromatrizz[42][187] = 9'b111111111;
assign micromatrizz[42][188] = 9'b111111111;
assign micromatrizz[42][189] = 9'b111111111;
assign micromatrizz[42][190] = 9'b111111111;
assign micromatrizz[42][191] = 9'b111111111;
assign micromatrizz[42][192] = 9'b111111111;
assign micromatrizz[42][193] = 9'b111111111;
assign micromatrizz[42][194] = 9'b111111111;
assign micromatrizz[42][195] = 9'b111111111;
assign micromatrizz[42][196] = 9'b111111111;
assign micromatrizz[42][197] = 9'b111111111;
assign micromatrizz[42][198] = 9'b111111111;
assign micromatrizz[42][199] = 9'b111111111;
assign micromatrizz[42][200] = 9'b111111111;
assign micromatrizz[42][201] = 9'b111111111;
assign micromatrizz[42][202] = 9'b111111111;
assign micromatrizz[42][203] = 9'b111111111;
assign micromatrizz[42][204] = 9'b111111111;
assign micromatrizz[42][205] = 9'b111111111;
assign micromatrizz[42][206] = 9'b111111111;
assign micromatrizz[42][207] = 9'b111111111;
assign micromatrizz[42][208] = 9'b111111111;
assign micromatrizz[42][209] = 9'b111111111;
assign micromatrizz[42][210] = 9'b111111111;
assign micromatrizz[42][211] = 9'b111111111;
assign micromatrizz[42][212] = 9'b111111111;
assign micromatrizz[42][213] = 9'b111111111;
assign micromatrizz[42][214] = 9'b111111111;
assign micromatrizz[42][215] = 9'b111111111;
assign micromatrizz[42][216] = 9'b111111111;
assign micromatrizz[42][217] = 9'b111111111;
assign micromatrizz[42][218] = 9'b111111111;
assign micromatrizz[42][219] = 9'b111111111;
assign micromatrizz[42][220] = 9'b111111111;
assign micromatrizz[42][221] = 9'b111111111;
assign micromatrizz[42][222] = 9'b111111111;
assign micromatrizz[42][223] = 9'b111111111;
assign micromatrizz[42][224] = 9'b111111111;
assign micromatrizz[42][225] = 9'b111111111;
assign micromatrizz[42][226] = 9'b111111111;
assign micromatrizz[42][227] = 9'b111111111;
assign micromatrizz[42][228] = 9'b111111111;
assign micromatrizz[42][229] = 9'b111111111;
assign micromatrizz[42][230] = 9'b111111111;
assign micromatrizz[42][231] = 9'b111111111;
assign micromatrizz[42][232] = 9'b111111111;
assign micromatrizz[42][233] = 9'b111111111;
assign micromatrizz[42][234] = 9'b111111111;
assign micromatrizz[42][235] = 9'b111111111;
assign micromatrizz[42][236] = 9'b111111111;
assign micromatrizz[42][237] = 9'b111111111;
assign micromatrizz[42][238] = 9'b111111111;
assign micromatrizz[42][239] = 9'b111111111;
assign micromatrizz[42][240] = 9'b111111111;
assign micromatrizz[42][241] = 9'b111111111;
assign micromatrizz[42][242] = 9'b111111111;
assign micromatrizz[42][243] = 9'b111111111;
assign micromatrizz[42][244] = 9'b111111111;
assign micromatrizz[42][245] = 9'b111111111;
assign micromatrizz[42][246] = 9'b111111111;
assign micromatrizz[42][247] = 9'b111111111;
assign micromatrizz[42][248] = 9'b111111111;
assign micromatrizz[42][249] = 9'b111111111;
assign micromatrizz[42][250] = 9'b111111111;
assign micromatrizz[42][251] = 9'b111111111;
assign micromatrizz[42][252] = 9'b111111111;
assign micromatrizz[42][253] = 9'b111111111;
assign micromatrizz[42][254] = 9'b111111111;
assign micromatrizz[42][255] = 9'b111111111;
assign micromatrizz[42][256] = 9'b111111111;
assign micromatrizz[42][257] = 9'b111111111;
assign micromatrizz[42][258] = 9'b111111111;
assign micromatrizz[42][259] = 9'b111111111;
assign micromatrizz[42][260] = 9'b111111111;
assign micromatrizz[42][261] = 9'b111111111;
assign micromatrizz[42][262] = 9'b111111111;
assign micromatrizz[42][263] = 9'b111111111;
assign micromatrizz[42][264] = 9'b111111111;
assign micromatrizz[42][265] = 9'b111111111;
assign micromatrizz[42][266] = 9'b111111111;
assign micromatrizz[42][267] = 9'b111111111;
assign micromatrizz[42][268] = 9'b111111111;
assign micromatrizz[42][269] = 9'b111111111;
assign micromatrizz[42][270] = 9'b111111111;
assign micromatrizz[42][271] = 9'b111111111;
assign micromatrizz[42][272] = 9'b111111111;
assign micromatrizz[42][273] = 9'b111111111;
assign micromatrizz[42][274] = 9'b111111111;
assign micromatrizz[42][275] = 9'b111111111;
assign micromatrizz[42][276] = 9'b111111111;
assign micromatrizz[42][277] = 9'b111111111;
assign micromatrizz[42][278] = 9'b111111111;
assign micromatrizz[42][279] = 9'b111111111;
assign micromatrizz[42][280] = 9'b111111111;
assign micromatrizz[42][281] = 9'b111111111;
assign micromatrizz[42][282] = 9'b111111111;
assign micromatrizz[42][283] = 9'b111111111;
assign micromatrizz[42][284] = 9'b111111111;
assign micromatrizz[42][285] = 9'b111111111;
assign micromatrizz[42][286] = 9'b111111111;
assign micromatrizz[42][287] = 9'b111111111;
assign micromatrizz[42][288] = 9'b111111111;
assign micromatrizz[42][289] = 9'b111111111;
assign micromatrizz[42][290] = 9'b111111111;
assign micromatrizz[42][291] = 9'b111111111;
assign micromatrizz[42][292] = 9'b111111111;
assign micromatrizz[42][293] = 9'b111111111;
assign micromatrizz[42][294] = 9'b111111111;
assign micromatrizz[42][295] = 9'b111111111;
assign micromatrizz[42][296] = 9'b111111111;
assign micromatrizz[42][297] = 9'b111111111;
assign micromatrizz[42][298] = 9'b111111111;
assign micromatrizz[42][299] = 9'b111111111;
assign micromatrizz[42][300] = 9'b111111111;
assign micromatrizz[42][301] = 9'b111111111;
assign micromatrizz[42][302] = 9'b111111111;
assign micromatrizz[42][303] = 9'b111111111;
assign micromatrizz[42][304] = 9'b111111111;
assign micromatrizz[42][305] = 9'b111111111;
assign micromatrizz[42][306] = 9'b111111111;
assign micromatrizz[42][307] = 9'b111111111;
assign micromatrizz[42][308] = 9'b111111111;
assign micromatrizz[42][309] = 9'b111111111;
assign micromatrizz[42][310] = 9'b111111111;
assign micromatrizz[42][311] = 9'b111111111;
assign micromatrizz[42][312] = 9'b111111111;
assign micromatrizz[42][313] = 9'b111111111;
assign micromatrizz[42][314] = 9'b111111111;
assign micromatrizz[42][315] = 9'b111111111;
assign micromatrizz[42][316] = 9'b111111111;
assign micromatrizz[42][317] = 9'b111111111;
assign micromatrizz[42][318] = 9'b111111111;
assign micromatrizz[42][319] = 9'b111111111;
assign micromatrizz[42][320] = 9'b111111111;
assign micromatrizz[42][321] = 9'b111111111;
assign micromatrizz[42][322] = 9'b111111111;
assign micromatrizz[42][323] = 9'b111111111;
assign micromatrizz[42][324] = 9'b111111111;
assign micromatrizz[42][325] = 9'b111111111;
assign micromatrizz[42][326] = 9'b111111111;
assign micromatrizz[42][327] = 9'b111111111;
assign micromatrizz[42][328] = 9'b111111111;
assign micromatrizz[42][329] = 9'b111111111;
assign micromatrizz[42][330] = 9'b111111111;
assign micromatrizz[42][331] = 9'b111111111;
assign micromatrizz[42][332] = 9'b111111111;
assign micromatrizz[42][333] = 9'b111111111;
assign micromatrizz[42][334] = 9'b111111111;
assign micromatrizz[42][335] = 9'b111111111;
assign micromatrizz[42][336] = 9'b111111111;
assign micromatrizz[42][337] = 9'b111111111;
assign micromatrizz[42][338] = 9'b111111111;
assign micromatrizz[42][339] = 9'b111111111;
assign micromatrizz[42][340] = 9'b111111111;
assign micromatrizz[42][341] = 9'b111111111;
assign micromatrizz[42][342] = 9'b111111111;
assign micromatrizz[42][343] = 9'b111111111;
assign micromatrizz[42][344] = 9'b111111111;
assign micromatrizz[42][345] = 9'b111111111;
assign micromatrizz[42][346] = 9'b111111111;
assign micromatrizz[42][347] = 9'b111111111;
assign micromatrizz[42][348] = 9'b111111111;
assign micromatrizz[42][349] = 9'b111111111;
assign micromatrizz[42][350] = 9'b111111111;
assign micromatrizz[42][351] = 9'b111111111;
assign micromatrizz[42][352] = 9'b111111111;
assign micromatrizz[42][353] = 9'b111111111;
assign micromatrizz[42][354] = 9'b111111111;
assign micromatrizz[42][355] = 9'b111111111;
assign micromatrizz[42][356] = 9'b111111111;
assign micromatrizz[42][357] = 9'b111111111;
assign micromatrizz[42][358] = 9'b111111111;
assign micromatrizz[42][359] = 9'b111111111;
assign micromatrizz[42][360] = 9'b111111111;
assign micromatrizz[42][361] = 9'b111111111;
assign micromatrizz[42][362] = 9'b111111111;
assign micromatrizz[42][363] = 9'b111111111;
assign micromatrizz[42][364] = 9'b111111111;
assign micromatrizz[42][365] = 9'b111111111;
assign micromatrizz[42][366] = 9'b111111111;
assign micromatrizz[42][367] = 9'b111111111;
assign micromatrizz[42][368] = 9'b111111111;
assign micromatrizz[42][369] = 9'b111111111;
assign micromatrizz[42][370] = 9'b111111111;
assign micromatrizz[42][371] = 9'b111111111;
assign micromatrizz[42][372] = 9'b111111111;
assign micromatrizz[42][373] = 9'b111111111;
assign micromatrizz[42][374] = 9'b111111111;
assign micromatrizz[42][375] = 9'b111111111;
assign micromatrizz[42][376] = 9'b111111111;
assign micromatrizz[42][377] = 9'b111111111;
assign micromatrizz[42][378] = 9'b111111111;
assign micromatrizz[42][379] = 9'b111111111;
assign micromatrizz[42][380] = 9'b111111111;
assign micromatrizz[42][381] = 9'b111111111;
assign micromatrizz[42][382] = 9'b111111111;
assign micromatrizz[42][383] = 9'b111111111;
assign micromatrizz[42][384] = 9'b111111111;
assign micromatrizz[42][385] = 9'b111111111;
assign micromatrizz[42][386] = 9'b111111111;
assign micromatrizz[42][387] = 9'b111111111;
assign micromatrizz[42][388] = 9'b111111111;
assign micromatrizz[42][389] = 9'b111111111;
assign micromatrizz[42][390] = 9'b111111111;
assign micromatrizz[42][391] = 9'b111111111;
assign micromatrizz[42][392] = 9'b111111111;
assign micromatrizz[42][393] = 9'b111111111;
assign micromatrizz[42][394] = 9'b111111111;
assign micromatrizz[42][395] = 9'b111111111;
assign micromatrizz[42][396] = 9'b111111111;
assign micromatrizz[42][397] = 9'b111111111;
assign micromatrizz[42][398] = 9'b111111111;
assign micromatrizz[42][399] = 9'b111111111;
assign micromatrizz[42][400] = 9'b111111111;
assign micromatrizz[42][401] = 9'b111111111;
assign micromatrizz[42][402] = 9'b111111111;
assign micromatrizz[42][403] = 9'b111111111;
assign micromatrizz[42][404] = 9'b111111111;
assign micromatrizz[42][405] = 9'b111111111;
assign micromatrizz[42][406] = 9'b111111111;
assign micromatrizz[42][407] = 9'b111111111;
assign micromatrizz[42][408] = 9'b111111111;
assign micromatrizz[42][409] = 9'b111111111;
assign micromatrizz[42][410] = 9'b111111111;
assign micromatrizz[42][411] = 9'b111111111;
assign micromatrizz[42][412] = 9'b111111111;
assign micromatrizz[42][413] = 9'b111111111;
assign micromatrizz[42][414] = 9'b111111111;
assign micromatrizz[42][415] = 9'b111111111;
assign micromatrizz[42][416] = 9'b111111111;
assign micromatrizz[42][417] = 9'b111111111;
assign micromatrizz[42][418] = 9'b111111111;
assign micromatrizz[42][419] = 9'b111111111;
assign micromatrizz[42][420] = 9'b111111111;
assign micromatrizz[42][421] = 9'b111111111;
assign micromatrizz[42][422] = 9'b111111111;
assign micromatrizz[42][423] = 9'b111111111;
assign micromatrizz[42][424] = 9'b111111111;
assign micromatrizz[42][425] = 9'b111111111;
assign micromatrizz[42][426] = 9'b111111111;
assign micromatrizz[42][427] = 9'b111111111;
assign micromatrizz[42][428] = 9'b111111111;
assign micromatrizz[42][429] = 9'b111111111;
assign micromatrizz[42][430] = 9'b111111111;
assign micromatrizz[42][431] = 9'b111111111;
assign micromatrizz[42][432] = 9'b111111111;
assign micromatrizz[42][433] = 9'b111111111;
assign micromatrizz[42][434] = 9'b111111111;
assign micromatrizz[42][435] = 9'b111111111;
assign micromatrizz[42][436] = 9'b111111111;
assign micromatrizz[42][437] = 9'b111111111;
assign micromatrizz[42][438] = 9'b111111111;
assign micromatrizz[42][439] = 9'b111111111;
assign micromatrizz[42][440] = 9'b111111111;
assign micromatrizz[42][441] = 9'b111111111;
assign micromatrizz[42][442] = 9'b111111111;
assign micromatrizz[42][443] = 9'b111111111;
assign micromatrizz[42][444] = 9'b111111111;
assign micromatrizz[42][445] = 9'b111111111;
assign micromatrizz[42][446] = 9'b111111111;
assign micromatrizz[42][447] = 9'b111111111;
assign micromatrizz[42][448] = 9'b111111111;
assign micromatrizz[42][449] = 9'b111111111;
assign micromatrizz[42][450] = 9'b111111111;
assign micromatrizz[42][451] = 9'b111111111;
assign micromatrizz[42][452] = 9'b111111111;
assign micromatrizz[42][453] = 9'b111111111;
assign micromatrizz[42][454] = 9'b111111111;
assign micromatrizz[42][455] = 9'b111111111;
assign micromatrizz[42][456] = 9'b111111111;
assign micromatrizz[42][457] = 9'b111111111;
assign micromatrizz[42][458] = 9'b111111111;
assign micromatrizz[42][459] = 9'b111111111;
assign micromatrizz[42][460] = 9'b111111111;
assign micromatrizz[42][461] = 9'b111111111;
assign micromatrizz[42][462] = 9'b111111111;
assign micromatrizz[42][463] = 9'b111111111;
assign micromatrizz[42][464] = 9'b111111111;
assign micromatrizz[42][465] = 9'b111111111;
assign micromatrizz[42][466] = 9'b111111111;
assign micromatrizz[42][467] = 9'b111111111;
assign micromatrizz[42][468] = 9'b111111111;
assign micromatrizz[42][469] = 9'b111111111;
assign micromatrizz[42][470] = 9'b111111111;
assign micromatrizz[42][471] = 9'b111111111;
assign micromatrizz[42][472] = 9'b111111111;
assign micromatrizz[42][473] = 9'b111111111;
assign micromatrizz[42][474] = 9'b111111111;
assign micromatrizz[42][475] = 9'b111111111;
assign micromatrizz[42][476] = 9'b111111111;
assign micromatrizz[42][477] = 9'b111111111;
assign micromatrizz[42][478] = 9'b111111111;
assign micromatrizz[42][479] = 9'b111111111;
assign micromatrizz[42][480] = 9'b111111111;
assign micromatrizz[42][481] = 9'b111111111;
assign micromatrizz[42][482] = 9'b111111111;
assign micromatrizz[42][483] = 9'b111111111;
assign micromatrizz[42][484] = 9'b111111111;
assign micromatrizz[42][485] = 9'b111111111;
assign micromatrizz[42][486] = 9'b111111111;
assign micromatrizz[42][487] = 9'b111111111;
assign micromatrizz[42][488] = 9'b111111111;
assign micromatrizz[42][489] = 9'b111111111;
assign micromatrizz[42][490] = 9'b111111111;
assign micromatrizz[42][491] = 9'b111111111;
assign micromatrizz[42][492] = 9'b111111111;
assign micromatrizz[42][493] = 9'b111111111;
assign micromatrizz[42][494] = 9'b111111111;
assign micromatrizz[42][495] = 9'b111111111;
assign micromatrizz[42][496] = 9'b111111111;
assign micromatrizz[42][497] = 9'b111111111;
assign micromatrizz[42][498] = 9'b111111111;
assign micromatrizz[42][499] = 9'b111111111;
assign micromatrizz[42][500] = 9'b111111111;
assign micromatrizz[42][501] = 9'b111111111;
assign micromatrizz[42][502] = 9'b111111111;
assign micromatrizz[42][503] = 9'b111111111;
assign micromatrizz[42][504] = 9'b111111111;
assign micromatrizz[42][505] = 9'b111111111;
assign micromatrizz[42][506] = 9'b111111111;
assign micromatrizz[42][507] = 9'b111111111;
assign micromatrizz[42][508] = 9'b111111111;
assign micromatrizz[42][509] = 9'b111111111;
assign micromatrizz[42][510] = 9'b111111111;
assign micromatrizz[42][511] = 9'b111111111;
assign micromatrizz[42][512] = 9'b111111111;
assign micromatrizz[42][513] = 9'b111111111;
assign micromatrizz[42][514] = 9'b111111111;
assign micromatrizz[42][515] = 9'b111111111;
assign micromatrizz[42][516] = 9'b111111111;
assign micromatrizz[42][517] = 9'b111111111;
assign micromatrizz[42][518] = 9'b111111111;
assign micromatrizz[42][519] = 9'b111111111;
assign micromatrizz[42][520] = 9'b111111111;
assign micromatrizz[42][521] = 9'b111111111;
assign micromatrizz[42][522] = 9'b111111111;
assign micromatrizz[42][523] = 9'b111111111;
assign micromatrizz[42][524] = 9'b111111111;
assign micromatrizz[42][525] = 9'b111111111;
assign micromatrizz[42][526] = 9'b111111111;
assign micromatrizz[42][527] = 9'b111111111;
assign micromatrizz[42][528] = 9'b111111111;
assign micromatrizz[42][529] = 9'b111111111;
assign micromatrizz[42][530] = 9'b111111111;
assign micromatrizz[42][531] = 9'b111111111;
assign micromatrizz[42][532] = 9'b111111111;
assign micromatrizz[42][533] = 9'b111111111;
assign micromatrizz[42][534] = 9'b111111111;
assign micromatrizz[42][535] = 9'b111111111;
assign micromatrizz[42][536] = 9'b111111111;
assign micromatrizz[42][537] = 9'b111111111;
assign micromatrizz[42][538] = 9'b111111111;
assign micromatrizz[42][539] = 9'b111111111;
assign micromatrizz[42][540] = 9'b111111111;
assign micromatrizz[42][541] = 9'b111111111;
assign micromatrizz[42][542] = 9'b111111111;
assign micromatrizz[42][543] = 9'b111111111;
assign micromatrizz[42][544] = 9'b111111111;
assign micromatrizz[42][545] = 9'b111111111;
assign micromatrizz[42][546] = 9'b111111111;
assign micromatrizz[42][547] = 9'b111111111;
assign micromatrizz[42][548] = 9'b111111111;
assign micromatrizz[42][549] = 9'b111111111;
assign micromatrizz[42][550] = 9'b111111111;
assign micromatrizz[42][551] = 9'b111111111;
assign micromatrizz[42][552] = 9'b111111111;
assign micromatrizz[42][553] = 9'b111111111;
assign micromatrizz[42][554] = 9'b111111111;
assign micromatrizz[42][555] = 9'b111111111;
assign micromatrizz[42][556] = 9'b111111111;
assign micromatrizz[42][557] = 9'b111111111;
assign micromatrizz[42][558] = 9'b111111111;
assign micromatrizz[42][559] = 9'b111111111;
assign micromatrizz[42][560] = 9'b111111111;
assign micromatrizz[42][561] = 9'b111111111;
assign micromatrizz[42][562] = 9'b111111111;
assign micromatrizz[42][563] = 9'b111111111;
assign micromatrizz[42][564] = 9'b111111111;
assign micromatrizz[42][565] = 9'b111111111;
assign micromatrizz[42][566] = 9'b111111111;
assign micromatrizz[42][567] = 9'b111111111;
assign micromatrizz[42][568] = 9'b111111111;
assign micromatrizz[42][569] = 9'b111111111;
assign micromatrizz[42][570] = 9'b111111111;
assign micromatrizz[42][571] = 9'b111111111;
assign micromatrizz[42][572] = 9'b111111111;
assign micromatrizz[42][573] = 9'b111111111;
assign micromatrizz[42][574] = 9'b111111111;
assign micromatrizz[42][575] = 9'b111111111;
assign micromatrizz[42][576] = 9'b111111111;
assign micromatrizz[42][577] = 9'b111111111;
assign micromatrizz[42][578] = 9'b111111111;
assign micromatrizz[42][579] = 9'b111111111;
assign micromatrizz[42][580] = 9'b111111111;
assign micromatrizz[42][581] = 9'b111111111;
assign micromatrizz[42][582] = 9'b111111111;
assign micromatrizz[42][583] = 9'b111111111;
assign micromatrizz[42][584] = 9'b111111111;
assign micromatrizz[42][585] = 9'b111111111;
assign micromatrizz[42][586] = 9'b111111111;
assign micromatrizz[42][587] = 9'b111111111;
assign micromatrizz[42][588] = 9'b111111111;
assign micromatrizz[42][589] = 9'b111111111;
assign micromatrizz[42][590] = 9'b111111111;
assign micromatrizz[42][591] = 9'b111111111;
assign micromatrizz[42][592] = 9'b111111111;
assign micromatrizz[42][593] = 9'b111111111;
assign micromatrizz[42][594] = 9'b111111111;
assign micromatrizz[42][595] = 9'b111111111;
assign micromatrizz[42][596] = 9'b111111111;
assign micromatrizz[42][597] = 9'b111111111;
assign micromatrizz[42][598] = 9'b111111111;
assign micromatrizz[42][599] = 9'b111111111;
assign micromatrizz[42][600] = 9'b111111111;
assign micromatrizz[42][601] = 9'b111111111;
assign micromatrizz[42][602] = 9'b111111111;
assign micromatrizz[42][603] = 9'b111111111;
assign micromatrizz[42][604] = 9'b111111111;
assign micromatrizz[42][605] = 9'b111111111;
assign micromatrizz[42][606] = 9'b111111111;
assign micromatrizz[42][607] = 9'b111111111;
assign micromatrizz[42][608] = 9'b111111111;
assign micromatrizz[42][609] = 9'b111111111;
assign micromatrizz[42][610] = 9'b111111111;
assign micromatrizz[42][611] = 9'b111111111;
assign micromatrizz[42][612] = 9'b111111111;
assign micromatrizz[42][613] = 9'b111111111;
assign micromatrizz[42][614] = 9'b111111111;
assign micromatrizz[42][615] = 9'b111111111;
assign micromatrizz[42][616] = 9'b111111111;
assign micromatrizz[42][617] = 9'b111111111;
assign micromatrizz[42][618] = 9'b111111111;
assign micromatrizz[42][619] = 9'b111111111;
assign micromatrizz[42][620] = 9'b111111111;
assign micromatrizz[42][621] = 9'b111111111;
assign micromatrizz[42][622] = 9'b111111111;
assign micromatrizz[42][623] = 9'b111111111;
assign micromatrizz[42][624] = 9'b111111111;
assign micromatrizz[42][625] = 9'b111111111;
assign micromatrizz[42][626] = 9'b111111111;
assign micromatrizz[42][627] = 9'b111111111;
assign micromatrizz[42][628] = 9'b111111111;
assign micromatrizz[42][629] = 9'b111111111;
assign micromatrizz[42][630] = 9'b111111111;
assign micromatrizz[42][631] = 9'b111111111;
assign micromatrizz[42][632] = 9'b111111111;
assign micromatrizz[42][633] = 9'b111111111;
assign micromatrizz[42][634] = 9'b111111111;
assign micromatrizz[42][635] = 9'b111111111;
assign micromatrizz[42][636] = 9'b111111111;
assign micromatrizz[42][637] = 9'b111111111;
assign micromatrizz[42][638] = 9'b111111111;
assign micromatrizz[42][639] = 9'b111111111;
assign micromatrizz[43][0] = 9'b111111111;
assign micromatrizz[43][1] = 9'b111111111;
assign micromatrizz[43][2] = 9'b111111111;
assign micromatrizz[43][3] = 9'b111111111;
assign micromatrizz[43][4] = 9'b111111111;
assign micromatrizz[43][5] = 9'b111111111;
assign micromatrizz[43][6] = 9'b111111111;
assign micromatrizz[43][7] = 9'b111111111;
assign micromatrizz[43][8] = 9'b111111111;
assign micromatrizz[43][9] = 9'b111111111;
assign micromatrizz[43][10] = 9'b111111111;
assign micromatrizz[43][11] = 9'b111111111;
assign micromatrizz[43][12] = 9'b111111111;
assign micromatrizz[43][13] = 9'b111111111;
assign micromatrizz[43][14] = 9'b111111111;
assign micromatrizz[43][15] = 9'b111111111;
assign micromatrizz[43][16] = 9'b111111111;
assign micromatrizz[43][17] = 9'b111111111;
assign micromatrizz[43][18] = 9'b111111111;
assign micromatrizz[43][19] = 9'b111111111;
assign micromatrizz[43][20] = 9'b111111111;
assign micromatrizz[43][21] = 9'b111111111;
assign micromatrizz[43][22] = 9'b111111111;
assign micromatrizz[43][23] = 9'b111111111;
assign micromatrizz[43][24] = 9'b111111111;
assign micromatrizz[43][25] = 9'b111111111;
assign micromatrizz[43][26] = 9'b111111111;
assign micromatrizz[43][27] = 9'b111111111;
assign micromatrizz[43][28] = 9'b111111111;
assign micromatrizz[43][29] = 9'b111111111;
assign micromatrizz[43][30] = 9'b111111111;
assign micromatrizz[43][31] = 9'b111111111;
assign micromatrizz[43][32] = 9'b111111111;
assign micromatrizz[43][33] = 9'b111111111;
assign micromatrizz[43][34] = 9'b111111111;
assign micromatrizz[43][35] = 9'b111111111;
assign micromatrizz[43][36] = 9'b111111111;
assign micromatrizz[43][37] = 9'b111111111;
assign micromatrizz[43][38] = 9'b111111111;
assign micromatrizz[43][39] = 9'b111111111;
assign micromatrizz[43][40] = 9'b111111111;
assign micromatrizz[43][41] = 9'b111111111;
assign micromatrizz[43][42] = 9'b111111111;
assign micromatrizz[43][43] = 9'b111111111;
assign micromatrizz[43][44] = 9'b111111111;
assign micromatrizz[43][45] = 9'b111111111;
assign micromatrizz[43][46] = 9'b111111111;
assign micromatrizz[43][47] = 9'b111111111;
assign micromatrizz[43][48] = 9'b111111111;
assign micromatrizz[43][49] = 9'b111111111;
assign micromatrizz[43][50] = 9'b111111111;
assign micromatrizz[43][51] = 9'b111111111;
assign micromatrizz[43][52] = 9'b111111111;
assign micromatrizz[43][53] = 9'b111111111;
assign micromatrizz[43][54] = 9'b111111111;
assign micromatrizz[43][55] = 9'b111111111;
assign micromatrizz[43][56] = 9'b111111111;
assign micromatrizz[43][57] = 9'b111111111;
assign micromatrizz[43][58] = 9'b111111111;
assign micromatrizz[43][59] = 9'b111111111;
assign micromatrizz[43][60] = 9'b111111111;
assign micromatrizz[43][61] = 9'b111111111;
assign micromatrizz[43][62] = 9'b111111111;
assign micromatrizz[43][63] = 9'b111111111;
assign micromatrizz[43][64] = 9'b111111111;
assign micromatrizz[43][65] = 9'b111111111;
assign micromatrizz[43][66] = 9'b111111111;
assign micromatrizz[43][67] = 9'b111111111;
assign micromatrizz[43][68] = 9'b111111111;
assign micromatrizz[43][69] = 9'b111111111;
assign micromatrizz[43][70] = 9'b111111111;
assign micromatrizz[43][71] = 9'b111111111;
assign micromatrizz[43][72] = 9'b111111111;
assign micromatrizz[43][73] = 9'b111111111;
assign micromatrizz[43][74] = 9'b111111111;
assign micromatrizz[43][75] = 9'b111111111;
assign micromatrizz[43][76] = 9'b111111111;
assign micromatrizz[43][77] = 9'b111111111;
assign micromatrizz[43][78] = 9'b111111111;
assign micromatrizz[43][79] = 9'b111111111;
assign micromatrizz[43][80] = 9'b111111111;
assign micromatrizz[43][81] = 9'b111111111;
assign micromatrizz[43][82] = 9'b111111111;
assign micromatrizz[43][83] = 9'b111111111;
assign micromatrizz[43][84] = 9'b111111111;
assign micromatrizz[43][85] = 9'b111111111;
assign micromatrizz[43][86] = 9'b111111111;
assign micromatrizz[43][87] = 9'b111111111;
assign micromatrizz[43][88] = 9'b111111111;
assign micromatrizz[43][89] = 9'b111111111;
assign micromatrizz[43][90] = 9'b111111111;
assign micromatrizz[43][91] = 9'b111111111;
assign micromatrizz[43][92] = 9'b111111111;
assign micromatrizz[43][93] = 9'b111111111;
assign micromatrizz[43][94] = 9'b111111111;
assign micromatrizz[43][95] = 9'b111111111;
assign micromatrizz[43][96] = 9'b111111111;
assign micromatrizz[43][97] = 9'b111111111;
assign micromatrizz[43][98] = 9'b111111111;
assign micromatrizz[43][99] = 9'b111111111;
assign micromatrizz[43][100] = 9'b111111111;
assign micromatrizz[43][101] = 9'b111111111;
assign micromatrizz[43][102] = 9'b111111111;
assign micromatrizz[43][103] = 9'b111111111;
assign micromatrizz[43][104] = 9'b111111111;
assign micromatrizz[43][105] = 9'b111111111;
assign micromatrizz[43][106] = 9'b111111111;
assign micromatrizz[43][107] = 9'b111111111;
assign micromatrizz[43][108] = 9'b111111111;
assign micromatrizz[43][109] = 9'b111111111;
assign micromatrizz[43][110] = 9'b111111111;
assign micromatrizz[43][111] = 9'b111111111;
assign micromatrizz[43][112] = 9'b111111111;
assign micromatrizz[43][113] = 9'b111111111;
assign micromatrizz[43][114] = 9'b111111111;
assign micromatrizz[43][115] = 9'b111111111;
assign micromatrizz[43][116] = 9'b111111111;
assign micromatrizz[43][117] = 9'b111111111;
assign micromatrizz[43][118] = 9'b111111111;
assign micromatrizz[43][119] = 9'b111111111;
assign micromatrizz[43][120] = 9'b111111111;
assign micromatrizz[43][121] = 9'b111111111;
assign micromatrizz[43][122] = 9'b111111111;
assign micromatrizz[43][123] = 9'b111111111;
assign micromatrizz[43][124] = 9'b111111111;
assign micromatrizz[43][125] = 9'b111111111;
assign micromatrizz[43][126] = 9'b111111111;
assign micromatrizz[43][127] = 9'b111111111;
assign micromatrizz[43][128] = 9'b111111111;
assign micromatrizz[43][129] = 9'b111111111;
assign micromatrizz[43][130] = 9'b111111111;
assign micromatrizz[43][131] = 9'b111111111;
assign micromatrizz[43][132] = 9'b111111111;
assign micromatrizz[43][133] = 9'b111111111;
assign micromatrizz[43][134] = 9'b111111111;
assign micromatrizz[43][135] = 9'b111111111;
assign micromatrizz[43][136] = 9'b111111111;
assign micromatrizz[43][137] = 9'b111111111;
assign micromatrizz[43][138] = 9'b111111111;
assign micromatrizz[43][139] = 9'b111111111;
assign micromatrizz[43][140] = 9'b111111111;
assign micromatrizz[43][141] = 9'b111111111;
assign micromatrizz[43][142] = 9'b111111111;
assign micromatrizz[43][143] = 9'b111111111;
assign micromatrizz[43][144] = 9'b111111111;
assign micromatrizz[43][145] = 9'b111111111;
assign micromatrizz[43][146] = 9'b111111111;
assign micromatrizz[43][147] = 9'b111111111;
assign micromatrizz[43][148] = 9'b111111111;
assign micromatrizz[43][149] = 9'b111111111;
assign micromatrizz[43][150] = 9'b111111111;
assign micromatrizz[43][151] = 9'b111111111;
assign micromatrizz[43][152] = 9'b111111111;
assign micromatrizz[43][153] = 9'b111111111;
assign micromatrizz[43][154] = 9'b111111111;
assign micromatrizz[43][155] = 9'b111111111;
assign micromatrizz[43][156] = 9'b111111111;
assign micromatrizz[43][157] = 9'b111111111;
assign micromatrizz[43][158] = 9'b111111111;
assign micromatrizz[43][159] = 9'b111111111;
assign micromatrizz[43][160] = 9'b111111111;
assign micromatrizz[43][161] = 9'b111111111;
assign micromatrizz[43][162] = 9'b111111111;
assign micromatrizz[43][163] = 9'b111111111;
assign micromatrizz[43][164] = 9'b111111111;
assign micromatrizz[43][165] = 9'b111111111;
assign micromatrizz[43][166] = 9'b111111111;
assign micromatrizz[43][167] = 9'b111111111;
assign micromatrizz[43][168] = 9'b111111111;
assign micromatrizz[43][169] = 9'b111111111;
assign micromatrizz[43][170] = 9'b111111111;
assign micromatrizz[43][171] = 9'b111111111;
assign micromatrizz[43][172] = 9'b111111111;
assign micromatrizz[43][173] = 9'b111111111;
assign micromatrizz[43][174] = 9'b111111111;
assign micromatrizz[43][175] = 9'b111111111;
assign micromatrizz[43][176] = 9'b111111111;
assign micromatrizz[43][177] = 9'b111111111;
assign micromatrizz[43][178] = 9'b111111111;
assign micromatrizz[43][179] = 9'b111111111;
assign micromatrizz[43][180] = 9'b111111111;
assign micromatrizz[43][181] = 9'b111111111;
assign micromatrizz[43][182] = 9'b111111111;
assign micromatrizz[43][183] = 9'b111111111;
assign micromatrizz[43][184] = 9'b111111111;
assign micromatrizz[43][185] = 9'b111111111;
assign micromatrizz[43][186] = 9'b111111111;
assign micromatrizz[43][187] = 9'b111111111;
assign micromatrizz[43][188] = 9'b111111111;
assign micromatrizz[43][189] = 9'b111111111;
assign micromatrizz[43][190] = 9'b111111111;
assign micromatrizz[43][191] = 9'b111111111;
assign micromatrizz[43][192] = 9'b111111111;
assign micromatrizz[43][193] = 9'b111111111;
assign micromatrizz[43][194] = 9'b111111111;
assign micromatrizz[43][195] = 9'b111111111;
assign micromatrizz[43][196] = 9'b111111111;
assign micromatrizz[43][197] = 9'b111111111;
assign micromatrizz[43][198] = 9'b111111111;
assign micromatrizz[43][199] = 9'b111111111;
assign micromatrizz[43][200] = 9'b111111111;
assign micromatrizz[43][201] = 9'b111111111;
assign micromatrizz[43][202] = 9'b111111111;
assign micromatrizz[43][203] = 9'b111111111;
assign micromatrizz[43][204] = 9'b111111111;
assign micromatrizz[43][205] = 9'b111111111;
assign micromatrizz[43][206] = 9'b111111111;
assign micromatrizz[43][207] = 9'b111111111;
assign micromatrizz[43][208] = 9'b111111111;
assign micromatrizz[43][209] = 9'b111111111;
assign micromatrizz[43][210] = 9'b111111111;
assign micromatrizz[43][211] = 9'b111111111;
assign micromatrizz[43][212] = 9'b111111111;
assign micromatrizz[43][213] = 9'b111111111;
assign micromatrizz[43][214] = 9'b111111111;
assign micromatrizz[43][215] = 9'b111111111;
assign micromatrizz[43][216] = 9'b111111111;
assign micromatrizz[43][217] = 9'b111111111;
assign micromatrizz[43][218] = 9'b111111111;
assign micromatrizz[43][219] = 9'b111111111;
assign micromatrizz[43][220] = 9'b111111111;
assign micromatrizz[43][221] = 9'b111111111;
assign micromatrizz[43][222] = 9'b111111111;
assign micromatrizz[43][223] = 9'b111111111;
assign micromatrizz[43][224] = 9'b111111111;
assign micromatrizz[43][225] = 9'b111111111;
assign micromatrizz[43][226] = 9'b111111111;
assign micromatrizz[43][227] = 9'b111111111;
assign micromatrizz[43][228] = 9'b111111111;
assign micromatrizz[43][229] = 9'b111111111;
assign micromatrizz[43][230] = 9'b111111111;
assign micromatrizz[43][231] = 9'b111111111;
assign micromatrizz[43][232] = 9'b111111111;
assign micromatrizz[43][233] = 9'b111111111;
assign micromatrizz[43][234] = 9'b111111111;
assign micromatrizz[43][235] = 9'b111111111;
assign micromatrizz[43][236] = 9'b111111111;
assign micromatrizz[43][237] = 9'b111111111;
assign micromatrizz[43][238] = 9'b111111111;
assign micromatrizz[43][239] = 9'b111111111;
assign micromatrizz[43][240] = 9'b111111111;
assign micromatrizz[43][241] = 9'b111111111;
assign micromatrizz[43][242] = 9'b111111111;
assign micromatrizz[43][243] = 9'b111111111;
assign micromatrizz[43][244] = 9'b111111111;
assign micromatrizz[43][245] = 9'b111111111;
assign micromatrizz[43][246] = 9'b111111111;
assign micromatrizz[43][247] = 9'b111111111;
assign micromatrizz[43][248] = 9'b111111111;
assign micromatrizz[43][249] = 9'b111111111;
assign micromatrizz[43][250] = 9'b111111111;
assign micromatrizz[43][251] = 9'b111111111;
assign micromatrizz[43][252] = 9'b111111111;
assign micromatrizz[43][253] = 9'b111111111;
assign micromatrizz[43][254] = 9'b111111111;
assign micromatrizz[43][255] = 9'b111111111;
assign micromatrizz[43][256] = 9'b111111111;
assign micromatrizz[43][257] = 9'b111111111;
assign micromatrizz[43][258] = 9'b111111111;
assign micromatrizz[43][259] = 9'b111111111;
assign micromatrizz[43][260] = 9'b111111111;
assign micromatrizz[43][261] = 9'b111111111;
assign micromatrizz[43][262] = 9'b111111111;
assign micromatrizz[43][263] = 9'b111111111;
assign micromatrizz[43][264] = 9'b111111111;
assign micromatrizz[43][265] = 9'b111111111;
assign micromatrizz[43][266] = 9'b111111111;
assign micromatrizz[43][267] = 9'b111111111;
assign micromatrizz[43][268] = 9'b111111111;
assign micromatrizz[43][269] = 9'b111111111;
assign micromatrizz[43][270] = 9'b111111111;
assign micromatrizz[43][271] = 9'b111111111;
assign micromatrizz[43][272] = 9'b111111111;
assign micromatrizz[43][273] = 9'b111111111;
assign micromatrizz[43][274] = 9'b111111111;
assign micromatrizz[43][275] = 9'b111111111;
assign micromatrizz[43][276] = 9'b111111111;
assign micromatrizz[43][277] = 9'b111111111;
assign micromatrizz[43][278] = 9'b111111111;
assign micromatrizz[43][279] = 9'b111111111;
assign micromatrizz[43][280] = 9'b111111111;
assign micromatrizz[43][281] = 9'b111111111;
assign micromatrizz[43][282] = 9'b111111111;
assign micromatrizz[43][283] = 9'b111111111;
assign micromatrizz[43][284] = 9'b111111111;
assign micromatrizz[43][285] = 9'b111111111;
assign micromatrizz[43][286] = 9'b111111111;
assign micromatrizz[43][287] = 9'b111111111;
assign micromatrizz[43][288] = 9'b111111111;
assign micromatrizz[43][289] = 9'b111111111;
assign micromatrizz[43][290] = 9'b111111111;
assign micromatrizz[43][291] = 9'b111111111;
assign micromatrizz[43][292] = 9'b111111111;
assign micromatrizz[43][293] = 9'b111111111;
assign micromatrizz[43][294] = 9'b111111111;
assign micromatrizz[43][295] = 9'b111111111;
assign micromatrizz[43][296] = 9'b111111111;
assign micromatrizz[43][297] = 9'b111111111;
assign micromatrizz[43][298] = 9'b111111111;
assign micromatrizz[43][299] = 9'b111111111;
assign micromatrizz[43][300] = 9'b111111111;
assign micromatrizz[43][301] = 9'b111111111;
assign micromatrizz[43][302] = 9'b111111111;
assign micromatrizz[43][303] = 9'b111111111;
assign micromatrizz[43][304] = 9'b111111111;
assign micromatrizz[43][305] = 9'b111111111;
assign micromatrizz[43][306] = 9'b111111111;
assign micromatrizz[43][307] = 9'b111111111;
assign micromatrizz[43][308] = 9'b111111111;
assign micromatrizz[43][309] = 9'b111111111;
assign micromatrizz[43][310] = 9'b111111111;
assign micromatrizz[43][311] = 9'b111111111;
assign micromatrizz[43][312] = 9'b111111111;
assign micromatrizz[43][313] = 9'b111111111;
assign micromatrizz[43][314] = 9'b111111111;
assign micromatrizz[43][315] = 9'b111111111;
assign micromatrizz[43][316] = 9'b111111111;
assign micromatrizz[43][317] = 9'b111111111;
assign micromatrizz[43][318] = 9'b111111111;
assign micromatrizz[43][319] = 9'b111111111;
assign micromatrizz[43][320] = 9'b111111111;
assign micromatrizz[43][321] = 9'b111111111;
assign micromatrizz[43][322] = 9'b111111111;
assign micromatrizz[43][323] = 9'b111111111;
assign micromatrizz[43][324] = 9'b111111111;
assign micromatrizz[43][325] = 9'b111111111;
assign micromatrizz[43][326] = 9'b111111111;
assign micromatrizz[43][327] = 9'b111111111;
assign micromatrizz[43][328] = 9'b111111111;
assign micromatrizz[43][329] = 9'b111111111;
assign micromatrizz[43][330] = 9'b111111111;
assign micromatrizz[43][331] = 9'b111111111;
assign micromatrizz[43][332] = 9'b111111111;
assign micromatrizz[43][333] = 9'b111111111;
assign micromatrizz[43][334] = 9'b111111111;
assign micromatrizz[43][335] = 9'b111111111;
assign micromatrizz[43][336] = 9'b111111111;
assign micromatrizz[43][337] = 9'b111111111;
assign micromatrizz[43][338] = 9'b111111111;
assign micromatrizz[43][339] = 9'b111111111;
assign micromatrizz[43][340] = 9'b111111111;
assign micromatrizz[43][341] = 9'b111111111;
assign micromatrizz[43][342] = 9'b111111111;
assign micromatrizz[43][343] = 9'b111111111;
assign micromatrizz[43][344] = 9'b111111111;
assign micromatrizz[43][345] = 9'b111111111;
assign micromatrizz[43][346] = 9'b111111111;
assign micromatrizz[43][347] = 9'b111111111;
assign micromatrizz[43][348] = 9'b111111111;
assign micromatrizz[43][349] = 9'b111111111;
assign micromatrizz[43][350] = 9'b111111111;
assign micromatrizz[43][351] = 9'b111111111;
assign micromatrizz[43][352] = 9'b111111111;
assign micromatrizz[43][353] = 9'b111111111;
assign micromatrizz[43][354] = 9'b111111111;
assign micromatrizz[43][355] = 9'b111111111;
assign micromatrizz[43][356] = 9'b111111111;
assign micromatrizz[43][357] = 9'b111111111;
assign micromatrizz[43][358] = 9'b111111111;
assign micromatrizz[43][359] = 9'b111111111;
assign micromatrizz[43][360] = 9'b111111111;
assign micromatrizz[43][361] = 9'b111111111;
assign micromatrizz[43][362] = 9'b111111111;
assign micromatrizz[43][363] = 9'b111111111;
assign micromatrizz[43][364] = 9'b111111111;
assign micromatrizz[43][365] = 9'b111111111;
assign micromatrizz[43][366] = 9'b111111111;
assign micromatrizz[43][367] = 9'b111111111;
assign micromatrizz[43][368] = 9'b111111111;
assign micromatrizz[43][369] = 9'b111111111;
assign micromatrizz[43][370] = 9'b111111111;
assign micromatrizz[43][371] = 9'b111111111;
assign micromatrizz[43][372] = 9'b111111111;
assign micromatrizz[43][373] = 9'b111111111;
assign micromatrizz[43][374] = 9'b111111111;
assign micromatrizz[43][375] = 9'b111111111;
assign micromatrizz[43][376] = 9'b111111111;
assign micromatrizz[43][377] = 9'b111111111;
assign micromatrizz[43][378] = 9'b111111111;
assign micromatrizz[43][379] = 9'b111111111;
assign micromatrizz[43][380] = 9'b111111111;
assign micromatrizz[43][381] = 9'b111111111;
assign micromatrizz[43][382] = 9'b111111111;
assign micromatrizz[43][383] = 9'b111111111;
assign micromatrizz[43][384] = 9'b111111111;
assign micromatrizz[43][385] = 9'b111111111;
assign micromatrizz[43][386] = 9'b111111111;
assign micromatrizz[43][387] = 9'b111111111;
assign micromatrizz[43][388] = 9'b111111111;
assign micromatrizz[43][389] = 9'b111111111;
assign micromatrizz[43][390] = 9'b111111111;
assign micromatrizz[43][391] = 9'b111111111;
assign micromatrizz[43][392] = 9'b111111111;
assign micromatrizz[43][393] = 9'b111111111;
assign micromatrizz[43][394] = 9'b111111111;
assign micromatrizz[43][395] = 9'b111111111;
assign micromatrizz[43][396] = 9'b111111111;
assign micromatrizz[43][397] = 9'b111111111;
assign micromatrizz[43][398] = 9'b111111111;
assign micromatrizz[43][399] = 9'b111111111;
assign micromatrizz[43][400] = 9'b111111111;
assign micromatrizz[43][401] = 9'b111111111;
assign micromatrizz[43][402] = 9'b111111111;
assign micromatrizz[43][403] = 9'b111111111;
assign micromatrizz[43][404] = 9'b111111111;
assign micromatrizz[43][405] = 9'b111111111;
assign micromatrizz[43][406] = 9'b111111111;
assign micromatrizz[43][407] = 9'b111111111;
assign micromatrizz[43][408] = 9'b111111111;
assign micromatrizz[43][409] = 9'b111111111;
assign micromatrizz[43][410] = 9'b111111111;
assign micromatrizz[43][411] = 9'b111111111;
assign micromatrizz[43][412] = 9'b111111111;
assign micromatrizz[43][413] = 9'b111111111;
assign micromatrizz[43][414] = 9'b111111111;
assign micromatrizz[43][415] = 9'b111111111;
assign micromatrizz[43][416] = 9'b111111111;
assign micromatrizz[43][417] = 9'b111111111;
assign micromatrizz[43][418] = 9'b111111111;
assign micromatrizz[43][419] = 9'b111111111;
assign micromatrizz[43][420] = 9'b111111111;
assign micromatrizz[43][421] = 9'b111111111;
assign micromatrizz[43][422] = 9'b111111111;
assign micromatrizz[43][423] = 9'b111111111;
assign micromatrizz[43][424] = 9'b111111111;
assign micromatrizz[43][425] = 9'b111111111;
assign micromatrizz[43][426] = 9'b111111111;
assign micromatrizz[43][427] = 9'b111111111;
assign micromatrizz[43][428] = 9'b111111111;
assign micromatrizz[43][429] = 9'b111111111;
assign micromatrizz[43][430] = 9'b111111111;
assign micromatrizz[43][431] = 9'b111111111;
assign micromatrizz[43][432] = 9'b111111111;
assign micromatrizz[43][433] = 9'b111111111;
assign micromatrizz[43][434] = 9'b111111111;
assign micromatrizz[43][435] = 9'b111111111;
assign micromatrizz[43][436] = 9'b111111111;
assign micromatrizz[43][437] = 9'b111111111;
assign micromatrizz[43][438] = 9'b111111111;
assign micromatrizz[43][439] = 9'b111111111;
assign micromatrizz[43][440] = 9'b111111111;
assign micromatrizz[43][441] = 9'b111111111;
assign micromatrizz[43][442] = 9'b111111111;
assign micromatrizz[43][443] = 9'b111111111;
assign micromatrizz[43][444] = 9'b111111111;
assign micromatrizz[43][445] = 9'b111111111;
assign micromatrizz[43][446] = 9'b111111111;
assign micromatrizz[43][447] = 9'b111111111;
assign micromatrizz[43][448] = 9'b111111111;
assign micromatrizz[43][449] = 9'b111111111;
assign micromatrizz[43][450] = 9'b111111111;
assign micromatrizz[43][451] = 9'b111111111;
assign micromatrizz[43][452] = 9'b111111111;
assign micromatrizz[43][453] = 9'b111111111;
assign micromatrizz[43][454] = 9'b111111111;
assign micromatrizz[43][455] = 9'b111111111;
assign micromatrizz[43][456] = 9'b111111111;
assign micromatrizz[43][457] = 9'b111111111;
assign micromatrizz[43][458] = 9'b111111111;
assign micromatrizz[43][459] = 9'b111111111;
assign micromatrizz[43][460] = 9'b111111111;
assign micromatrizz[43][461] = 9'b111111111;
assign micromatrizz[43][462] = 9'b111111111;
assign micromatrizz[43][463] = 9'b111111111;
assign micromatrizz[43][464] = 9'b111111111;
assign micromatrizz[43][465] = 9'b111111111;
assign micromatrizz[43][466] = 9'b111111111;
assign micromatrizz[43][467] = 9'b111111111;
assign micromatrizz[43][468] = 9'b111111111;
assign micromatrizz[43][469] = 9'b111111111;
assign micromatrizz[43][470] = 9'b111111111;
assign micromatrizz[43][471] = 9'b111111111;
assign micromatrizz[43][472] = 9'b111111111;
assign micromatrizz[43][473] = 9'b111111111;
assign micromatrizz[43][474] = 9'b111111111;
assign micromatrizz[43][475] = 9'b111111111;
assign micromatrizz[43][476] = 9'b111111111;
assign micromatrizz[43][477] = 9'b111111111;
assign micromatrizz[43][478] = 9'b111111111;
assign micromatrizz[43][479] = 9'b111111111;
assign micromatrizz[43][480] = 9'b111111111;
assign micromatrizz[43][481] = 9'b111111111;
assign micromatrizz[43][482] = 9'b111111111;
assign micromatrizz[43][483] = 9'b111111111;
assign micromatrizz[43][484] = 9'b111111111;
assign micromatrizz[43][485] = 9'b111111111;
assign micromatrizz[43][486] = 9'b111111111;
assign micromatrizz[43][487] = 9'b111111111;
assign micromatrizz[43][488] = 9'b111111111;
assign micromatrizz[43][489] = 9'b111111111;
assign micromatrizz[43][490] = 9'b111111111;
assign micromatrizz[43][491] = 9'b111111111;
assign micromatrizz[43][492] = 9'b111111111;
assign micromatrizz[43][493] = 9'b111111111;
assign micromatrizz[43][494] = 9'b111111111;
assign micromatrizz[43][495] = 9'b111111111;
assign micromatrizz[43][496] = 9'b111111111;
assign micromatrizz[43][497] = 9'b111111111;
assign micromatrizz[43][498] = 9'b111111111;
assign micromatrizz[43][499] = 9'b111111111;
assign micromatrizz[43][500] = 9'b111111111;
assign micromatrizz[43][501] = 9'b111111111;
assign micromatrizz[43][502] = 9'b111111111;
assign micromatrizz[43][503] = 9'b111111111;
assign micromatrizz[43][504] = 9'b111111111;
assign micromatrizz[43][505] = 9'b111111111;
assign micromatrizz[43][506] = 9'b111111111;
assign micromatrizz[43][507] = 9'b111111111;
assign micromatrizz[43][508] = 9'b111111111;
assign micromatrizz[43][509] = 9'b111111111;
assign micromatrizz[43][510] = 9'b111111111;
assign micromatrizz[43][511] = 9'b111111111;
assign micromatrizz[43][512] = 9'b111111111;
assign micromatrizz[43][513] = 9'b111111111;
assign micromatrizz[43][514] = 9'b111111111;
assign micromatrizz[43][515] = 9'b111111111;
assign micromatrizz[43][516] = 9'b111111111;
assign micromatrizz[43][517] = 9'b111111111;
assign micromatrizz[43][518] = 9'b111111111;
assign micromatrizz[43][519] = 9'b111111111;
assign micromatrizz[43][520] = 9'b111111111;
assign micromatrizz[43][521] = 9'b111111111;
assign micromatrizz[43][522] = 9'b111111111;
assign micromatrizz[43][523] = 9'b111111111;
assign micromatrizz[43][524] = 9'b111111111;
assign micromatrizz[43][525] = 9'b111111111;
assign micromatrizz[43][526] = 9'b111111111;
assign micromatrizz[43][527] = 9'b111111111;
assign micromatrizz[43][528] = 9'b111111111;
assign micromatrizz[43][529] = 9'b111111111;
assign micromatrizz[43][530] = 9'b111111111;
assign micromatrizz[43][531] = 9'b111111111;
assign micromatrizz[43][532] = 9'b111111111;
assign micromatrizz[43][533] = 9'b111111111;
assign micromatrizz[43][534] = 9'b111111111;
assign micromatrizz[43][535] = 9'b111111111;
assign micromatrizz[43][536] = 9'b111111111;
assign micromatrizz[43][537] = 9'b111111111;
assign micromatrizz[43][538] = 9'b111111111;
assign micromatrizz[43][539] = 9'b111111111;
assign micromatrizz[43][540] = 9'b111111111;
assign micromatrizz[43][541] = 9'b111111111;
assign micromatrizz[43][542] = 9'b111111111;
assign micromatrizz[43][543] = 9'b111111111;
assign micromatrizz[43][544] = 9'b111111111;
assign micromatrizz[43][545] = 9'b111111111;
assign micromatrizz[43][546] = 9'b111111111;
assign micromatrizz[43][547] = 9'b111111111;
assign micromatrizz[43][548] = 9'b111111111;
assign micromatrizz[43][549] = 9'b111111111;
assign micromatrizz[43][550] = 9'b111111111;
assign micromatrizz[43][551] = 9'b111111111;
assign micromatrizz[43][552] = 9'b111111111;
assign micromatrizz[43][553] = 9'b111111111;
assign micromatrizz[43][554] = 9'b111111111;
assign micromatrizz[43][555] = 9'b111111111;
assign micromatrizz[43][556] = 9'b111111111;
assign micromatrizz[43][557] = 9'b111111111;
assign micromatrizz[43][558] = 9'b111111111;
assign micromatrizz[43][559] = 9'b111111111;
assign micromatrizz[43][560] = 9'b111111111;
assign micromatrizz[43][561] = 9'b111111111;
assign micromatrizz[43][562] = 9'b111111111;
assign micromatrizz[43][563] = 9'b111111111;
assign micromatrizz[43][564] = 9'b111111111;
assign micromatrizz[43][565] = 9'b111111111;
assign micromatrizz[43][566] = 9'b111111111;
assign micromatrizz[43][567] = 9'b111111111;
assign micromatrizz[43][568] = 9'b111111111;
assign micromatrizz[43][569] = 9'b111111111;
assign micromatrizz[43][570] = 9'b111111111;
assign micromatrizz[43][571] = 9'b111111111;
assign micromatrizz[43][572] = 9'b111111111;
assign micromatrizz[43][573] = 9'b111111111;
assign micromatrizz[43][574] = 9'b111111111;
assign micromatrizz[43][575] = 9'b111111111;
assign micromatrizz[43][576] = 9'b111111111;
assign micromatrizz[43][577] = 9'b111111111;
assign micromatrizz[43][578] = 9'b111111111;
assign micromatrizz[43][579] = 9'b111111111;
assign micromatrizz[43][580] = 9'b111111111;
assign micromatrizz[43][581] = 9'b111111111;
assign micromatrizz[43][582] = 9'b111111111;
assign micromatrizz[43][583] = 9'b111111111;
assign micromatrizz[43][584] = 9'b111111111;
assign micromatrizz[43][585] = 9'b111111111;
assign micromatrizz[43][586] = 9'b111111111;
assign micromatrizz[43][587] = 9'b111111111;
assign micromatrizz[43][588] = 9'b111111111;
assign micromatrizz[43][589] = 9'b111111111;
assign micromatrizz[43][590] = 9'b111111111;
assign micromatrizz[43][591] = 9'b111111111;
assign micromatrizz[43][592] = 9'b111111111;
assign micromatrizz[43][593] = 9'b111111111;
assign micromatrizz[43][594] = 9'b111111111;
assign micromatrizz[43][595] = 9'b111111111;
assign micromatrizz[43][596] = 9'b111111111;
assign micromatrizz[43][597] = 9'b111111111;
assign micromatrizz[43][598] = 9'b111111111;
assign micromatrizz[43][599] = 9'b111111111;
assign micromatrizz[43][600] = 9'b111111111;
assign micromatrizz[43][601] = 9'b111111111;
assign micromatrizz[43][602] = 9'b111111111;
assign micromatrizz[43][603] = 9'b111111111;
assign micromatrizz[43][604] = 9'b111111111;
assign micromatrizz[43][605] = 9'b111111111;
assign micromatrizz[43][606] = 9'b111111111;
assign micromatrizz[43][607] = 9'b111111111;
assign micromatrizz[43][608] = 9'b111111111;
assign micromatrizz[43][609] = 9'b111111111;
assign micromatrizz[43][610] = 9'b111111111;
assign micromatrizz[43][611] = 9'b111111111;
assign micromatrizz[43][612] = 9'b111111111;
assign micromatrizz[43][613] = 9'b111111111;
assign micromatrizz[43][614] = 9'b111111111;
assign micromatrizz[43][615] = 9'b111111111;
assign micromatrizz[43][616] = 9'b111111111;
assign micromatrizz[43][617] = 9'b111111111;
assign micromatrizz[43][618] = 9'b111111111;
assign micromatrizz[43][619] = 9'b111111111;
assign micromatrizz[43][620] = 9'b111111111;
assign micromatrizz[43][621] = 9'b111111111;
assign micromatrizz[43][622] = 9'b111111111;
assign micromatrizz[43][623] = 9'b111111111;
assign micromatrizz[43][624] = 9'b111111111;
assign micromatrizz[43][625] = 9'b111111111;
assign micromatrizz[43][626] = 9'b111111111;
assign micromatrizz[43][627] = 9'b111111111;
assign micromatrizz[43][628] = 9'b111111111;
assign micromatrizz[43][629] = 9'b111111111;
assign micromatrizz[43][630] = 9'b111111111;
assign micromatrizz[43][631] = 9'b111111111;
assign micromatrizz[43][632] = 9'b111111111;
assign micromatrizz[43][633] = 9'b111111111;
assign micromatrizz[43][634] = 9'b111111111;
assign micromatrizz[43][635] = 9'b111111111;
assign micromatrizz[43][636] = 9'b111111111;
assign micromatrizz[43][637] = 9'b111111111;
assign micromatrizz[43][638] = 9'b111111111;
assign micromatrizz[43][639] = 9'b111111111;
assign micromatrizz[44][0] = 9'b111111111;
assign micromatrizz[44][1] = 9'b111111111;
assign micromatrizz[44][2] = 9'b111111111;
assign micromatrizz[44][3] = 9'b111111111;
assign micromatrizz[44][4] = 9'b111111111;
assign micromatrizz[44][5] = 9'b111111111;
assign micromatrizz[44][6] = 9'b111111111;
assign micromatrizz[44][7] = 9'b111111111;
assign micromatrizz[44][8] = 9'b111111111;
assign micromatrizz[44][9] = 9'b111111111;
assign micromatrizz[44][10] = 9'b111111111;
assign micromatrizz[44][11] = 9'b111111111;
assign micromatrizz[44][12] = 9'b111111111;
assign micromatrizz[44][13] = 9'b111111111;
assign micromatrizz[44][14] = 9'b111111111;
assign micromatrizz[44][15] = 9'b111111111;
assign micromatrizz[44][16] = 9'b111111111;
assign micromatrizz[44][17] = 9'b111111111;
assign micromatrizz[44][18] = 9'b111111111;
assign micromatrizz[44][19] = 9'b111111111;
assign micromatrizz[44][20] = 9'b111111111;
assign micromatrizz[44][21] = 9'b111111111;
assign micromatrizz[44][22] = 9'b111111111;
assign micromatrizz[44][23] = 9'b111111111;
assign micromatrizz[44][24] = 9'b111111111;
assign micromatrizz[44][25] = 9'b111111111;
assign micromatrizz[44][26] = 9'b111111111;
assign micromatrizz[44][27] = 9'b111111111;
assign micromatrizz[44][28] = 9'b111111111;
assign micromatrizz[44][29] = 9'b111111111;
assign micromatrizz[44][30] = 9'b111111111;
assign micromatrizz[44][31] = 9'b111111111;
assign micromatrizz[44][32] = 9'b111111111;
assign micromatrizz[44][33] = 9'b111111111;
assign micromatrizz[44][34] = 9'b111111111;
assign micromatrizz[44][35] = 9'b111111111;
assign micromatrizz[44][36] = 9'b111111111;
assign micromatrizz[44][37] = 9'b111111111;
assign micromatrizz[44][38] = 9'b111111111;
assign micromatrizz[44][39] = 9'b111111111;
assign micromatrizz[44][40] = 9'b111111111;
assign micromatrizz[44][41] = 9'b111111111;
assign micromatrizz[44][42] = 9'b111111111;
assign micromatrizz[44][43] = 9'b111111111;
assign micromatrizz[44][44] = 9'b111111111;
assign micromatrizz[44][45] = 9'b111111111;
assign micromatrizz[44][46] = 9'b111111111;
assign micromatrizz[44][47] = 9'b111111111;
assign micromatrizz[44][48] = 9'b111111111;
assign micromatrizz[44][49] = 9'b111111111;
assign micromatrizz[44][50] = 9'b111111111;
assign micromatrizz[44][51] = 9'b111111111;
assign micromatrizz[44][52] = 9'b111111111;
assign micromatrizz[44][53] = 9'b111111111;
assign micromatrizz[44][54] = 9'b111111111;
assign micromatrizz[44][55] = 9'b111111111;
assign micromatrizz[44][56] = 9'b111111111;
assign micromatrizz[44][57] = 9'b111111111;
assign micromatrizz[44][58] = 9'b111111111;
assign micromatrizz[44][59] = 9'b111111111;
assign micromatrizz[44][60] = 9'b111111111;
assign micromatrizz[44][61] = 9'b111111111;
assign micromatrizz[44][62] = 9'b111111111;
assign micromatrizz[44][63] = 9'b111111111;
assign micromatrizz[44][64] = 9'b111111111;
assign micromatrizz[44][65] = 9'b111111111;
assign micromatrizz[44][66] = 9'b111111111;
assign micromatrizz[44][67] = 9'b111111111;
assign micromatrizz[44][68] = 9'b111111111;
assign micromatrizz[44][69] = 9'b111111111;
assign micromatrizz[44][70] = 9'b111111111;
assign micromatrizz[44][71] = 9'b111111111;
assign micromatrizz[44][72] = 9'b111111111;
assign micromatrizz[44][73] = 9'b111111111;
assign micromatrizz[44][74] = 9'b111111111;
assign micromatrizz[44][75] = 9'b111111111;
assign micromatrizz[44][76] = 9'b111111111;
assign micromatrizz[44][77] = 9'b111111111;
assign micromatrizz[44][78] = 9'b111111111;
assign micromatrizz[44][79] = 9'b111111111;
assign micromatrizz[44][80] = 9'b111111111;
assign micromatrizz[44][81] = 9'b111111111;
assign micromatrizz[44][82] = 9'b111111111;
assign micromatrizz[44][83] = 9'b111111111;
assign micromatrizz[44][84] = 9'b111111111;
assign micromatrizz[44][85] = 9'b111111111;
assign micromatrizz[44][86] = 9'b111111111;
assign micromatrizz[44][87] = 9'b111111111;
assign micromatrizz[44][88] = 9'b111111111;
assign micromatrizz[44][89] = 9'b111111111;
assign micromatrizz[44][90] = 9'b111111111;
assign micromatrizz[44][91] = 9'b111111111;
assign micromatrizz[44][92] = 9'b111111111;
assign micromatrizz[44][93] = 9'b111111111;
assign micromatrizz[44][94] = 9'b111111111;
assign micromatrizz[44][95] = 9'b111111111;
assign micromatrizz[44][96] = 9'b111111111;
assign micromatrizz[44][97] = 9'b111111111;
assign micromatrizz[44][98] = 9'b111111111;
assign micromatrizz[44][99] = 9'b111111111;
assign micromatrizz[44][100] = 9'b111111111;
assign micromatrizz[44][101] = 9'b111111111;
assign micromatrizz[44][102] = 9'b111111111;
assign micromatrizz[44][103] = 9'b111111111;
assign micromatrizz[44][104] = 9'b111111111;
assign micromatrizz[44][105] = 9'b111111111;
assign micromatrizz[44][106] = 9'b111111111;
assign micromatrizz[44][107] = 9'b111111111;
assign micromatrizz[44][108] = 9'b111111111;
assign micromatrizz[44][109] = 9'b111111111;
assign micromatrizz[44][110] = 9'b111111111;
assign micromatrizz[44][111] = 9'b111111111;
assign micromatrizz[44][112] = 9'b111111111;
assign micromatrizz[44][113] = 9'b111111111;
assign micromatrizz[44][114] = 9'b111111111;
assign micromatrizz[44][115] = 9'b111111111;
assign micromatrizz[44][116] = 9'b111111111;
assign micromatrizz[44][117] = 9'b111111111;
assign micromatrizz[44][118] = 9'b111111111;
assign micromatrizz[44][119] = 9'b111111111;
assign micromatrizz[44][120] = 9'b111111111;
assign micromatrizz[44][121] = 9'b111111111;
assign micromatrizz[44][122] = 9'b111111111;
assign micromatrizz[44][123] = 9'b111111111;
assign micromatrizz[44][124] = 9'b111111111;
assign micromatrizz[44][125] = 9'b111111111;
assign micromatrizz[44][126] = 9'b111111111;
assign micromatrizz[44][127] = 9'b111111111;
assign micromatrizz[44][128] = 9'b111111111;
assign micromatrizz[44][129] = 9'b111111111;
assign micromatrizz[44][130] = 9'b111111111;
assign micromatrizz[44][131] = 9'b111111111;
assign micromatrizz[44][132] = 9'b111111111;
assign micromatrizz[44][133] = 9'b111111111;
assign micromatrizz[44][134] = 9'b111111111;
assign micromatrizz[44][135] = 9'b111111111;
assign micromatrizz[44][136] = 9'b111111111;
assign micromatrizz[44][137] = 9'b111111111;
assign micromatrizz[44][138] = 9'b111111111;
assign micromatrizz[44][139] = 9'b111111111;
assign micromatrizz[44][140] = 9'b111111111;
assign micromatrizz[44][141] = 9'b111111111;
assign micromatrizz[44][142] = 9'b111111111;
assign micromatrizz[44][143] = 9'b111111111;
assign micromatrizz[44][144] = 9'b111111111;
assign micromatrizz[44][145] = 9'b111111111;
assign micromatrizz[44][146] = 9'b111111111;
assign micromatrizz[44][147] = 9'b111111111;
assign micromatrizz[44][148] = 9'b111111111;
assign micromatrizz[44][149] = 9'b111111111;
assign micromatrizz[44][150] = 9'b111111111;
assign micromatrizz[44][151] = 9'b111111111;
assign micromatrizz[44][152] = 9'b111111111;
assign micromatrizz[44][153] = 9'b111111111;
assign micromatrizz[44][154] = 9'b111111111;
assign micromatrizz[44][155] = 9'b111111111;
assign micromatrizz[44][156] = 9'b111111111;
assign micromatrizz[44][157] = 9'b111111111;
assign micromatrizz[44][158] = 9'b111111111;
assign micromatrizz[44][159] = 9'b111111111;
assign micromatrizz[44][160] = 9'b111111111;
assign micromatrizz[44][161] = 9'b111111111;
assign micromatrizz[44][162] = 9'b111111111;
assign micromatrizz[44][163] = 9'b111111111;
assign micromatrizz[44][164] = 9'b111111111;
assign micromatrizz[44][165] = 9'b111111111;
assign micromatrizz[44][166] = 9'b111111111;
assign micromatrizz[44][167] = 9'b111111111;
assign micromatrizz[44][168] = 9'b111111111;
assign micromatrizz[44][169] = 9'b111111111;
assign micromatrizz[44][170] = 9'b111111111;
assign micromatrizz[44][171] = 9'b111111111;
assign micromatrizz[44][172] = 9'b111111111;
assign micromatrizz[44][173] = 9'b111111111;
assign micromatrizz[44][174] = 9'b111111111;
assign micromatrizz[44][175] = 9'b111111111;
assign micromatrizz[44][176] = 9'b111111111;
assign micromatrizz[44][177] = 9'b111111111;
assign micromatrizz[44][178] = 9'b111111111;
assign micromatrizz[44][179] = 9'b111111111;
assign micromatrizz[44][180] = 9'b111111111;
assign micromatrizz[44][181] = 9'b111111111;
assign micromatrizz[44][182] = 9'b111111111;
assign micromatrizz[44][183] = 9'b111111111;
assign micromatrizz[44][184] = 9'b111111111;
assign micromatrizz[44][185] = 9'b111111111;
assign micromatrizz[44][186] = 9'b111111111;
assign micromatrizz[44][187] = 9'b111111111;
assign micromatrizz[44][188] = 9'b111111111;
assign micromatrizz[44][189] = 9'b111111111;
assign micromatrizz[44][190] = 9'b111111111;
assign micromatrizz[44][191] = 9'b111111111;
assign micromatrizz[44][192] = 9'b111111111;
assign micromatrizz[44][193] = 9'b111111111;
assign micromatrizz[44][194] = 9'b111111111;
assign micromatrizz[44][195] = 9'b111111111;
assign micromatrizz[44][196] = 9'b111111111;
assign micromatrizz[44][197] = 9'b111111111;
assign micromatrizz[44][198] = 9'b111111111;
assign micromatrizz[44][199] = 9'b111111111;
assign micromatrizz[44][200] = 9'b111111111;
assign micromatrizz[44][201] = 9'b111111111;
assign micromatrizz[44][202] = 9'b111111111;
assign micromatrizz[44][203] = 9'b111111111;
assign micromatrizz[44][204] = 9'b111111111;
assign micromatrizz[44][205] = 9'b111111111;
assign micromatrizz[44][206] = 9'b111111111;
assign micromatrizz[44][207] = 9'b111111111;
assign micromatrizz[44][208] = 9'b111111111;
assign micromatrizz[44][209] = 9'b111111111;
assign micromatrizz[44][210] = 9'b111111111;
assign micromatrizz[44][211] = 9'b111111111;
assign micromatrizz[44][212] = 9'b111111111;
assign micromatrizz[44][213] = 9'b111111111;
assign micromatrizz[44][214] = 9'b111111111;
assign micromatrizz[44][215] = 9'b111111111;
assign micromatrizz[44][216] = 9'b111111111;
assign micromatrizz[44][217] = 9'b111111111;
assign micromatrizz[44][218] = 9'b111111111;
assign micromatrizz[44][219] = 9'b111111111;
assign micromatrizz[44][220] = 9'b111111111;
assign micromatrizz[44][221] = 9'b111111111;
assign micromatrizz[44][222] = 9'b111111111;
assign micromatrizz[44][223] = 9'b111111111;
assign micromatrizz[44][224] = 9'b111111111;
assign micromatrizz[44][225] = 9'b111111111;
assign micromatrizz[44][226] = 9'b111111111;
assign micromatrizz[44][227] = 9'b111111111;
assign micromatrizz[44][228] = 9'b111111111;
assign micromatrizz[44][229] = 9'b111111111;
assign micromatrizz[44][230] = 9'b111111111;
assign micromatrizz[44][231] = 9'b111111111;
assign micromatrizz[44][232] = 9'b111111111;
assign micromatrizz[44][233] = 9'b111111111;
assign micromatrizz[44][234] = 9'b111111111;
assign micromatrizz[44][235] = 9'b111111111;
assign micromatrizz[44][236] = 9'b111111111;
assign micromatrizz[44][237] = 9'b111111111;
assign micromatrizz[44][238] = 9'b111111111;
assign micromatrizz[44][239] = 9'b111111111;
assign micromatrizz[44][240] = 9'b111111111;
assign micromatrizz[44][241] = 9'b111111111;
assign micromatrizz[44][242] = 9'b111111111;
assign micromatrizz[44][243] = 9'b111111111;
assign micromatrizz[44][244] = 9'b111111111;
assign micromatrizz[44][245] = 9'b111111111;
assign micromatrizz[44][246] = 9'b111111111;
assign micromatrizz[44][247] = 9'b111111111;
assign micromatrizz[44][248] = 9'b111111111;
assign micromatrizz[44][249] = 9'b111111111;
assign micromatrizz[44][250] = 9'b111111111;
assign micromatrizz[44][251] = 9'b111111111;
assign micromatrizz[44][252] = 9'b111111111;
assign micromatrizz[44][253] = 9'b111111111;
assign micromatrizz[44][254] = 9'b111111111;
assign micromatrizz[44][255] = 9'b111111111;
assign micromatrizz[44][256] = 9'b111111111;
assign micromatrizz[44][257] = 9'b111111111;
assign micromatrizz[44][258] = 9'b111111111;
assign micromatrizz[44][259] = 9'b111111111;
assign micromatrizz[44][260] = 9'b111111111;
assign micromatrizz[44][261] = 9'b111111111;
assign micromatrizz[44][262] = 9'b111111111;
assign micromatrizz[44][263] = 9'b111111111;
assign micromatrizz[44][264] = 9'b111111111;
assign micromatrizz[44][265] = 9'b111111111;
assign micromatrizz[44][266] = 9'b111111111;
assign micromatrizz[44][267] = 9'b111111111;
assign micromatrizz[44][268] = 9'b111111111;
assign micromatrizz[44][269] = 9'b111111111;
assign micromatrizz[44][270] = 9'b111111111;
assign micromatrizz[44][271] = 9'b111111111;
assign micromatrizz[44][272] = 9'b111111111;
assign micromatrizz[44][273] = 9'b111111111;
assign micromatrizz[44][274] = 9'b111111111;
assign micromatrizz[44][275] = 9'b111111111;
assign micromatrizz[44][276] = 9'b111111111;
assign micromatrizz[44][277] = 9'b111111111;
assign micromatrizz[44][278] = 9'b111111111;
assign micromatrizz[44][279] = 9'b111111111;
assign micromatrizz[44][280] = 9'b111111111;
assign micromatrizz[44][281] = 9'b111111111;
assign micromatrizz[44][282] = 9'b111111111;
assign micromatrizz[44][283] = 9'b111111111;
assign micromatrizz[44][284] = 9'b111111111;
assign micromatrizz[44][285] = 9'b111111111;
assign micromatrizz[44][286] = 9'b111111111;
assign micromatrizz[44][287] = 9'b111111111;
assign micromatrizz[44][288] = 9'b111111111;
assign micromatrizz[44][289] = 9'b111111111;
assign micromatrizz[44][290] = 9'b111111111;
assign micromatrizz[44][291] = 9'b111111111;
assign micromatrizz[44][292] = 9'b111111111;
assign micromatrizz[44][293] = 9'b111111111;
assign micromatrizz[44][294] = 9'b111111111;
assign micromatrizz[44][295] = 9'b111111111;
assign micromatrizz[44][296] = 9'b111111111;
assign micromatrizz[44][297] = 9'b111111111;
assign micromatrizz[44][298] = 9'b111111111;
assign micromatrizz[44][299] = 9'b111111111;
assign micromatrizz[44][300] = 9'b111111111;
assign micromatrizz[44][301] = 9'b111111111;
assign micromatrizz[44][302] = 9'b111111111;
assign micromatrizz[44][303] = 9'b111111111;
assign micromatrizz[44][304] = 9'b111111111;
assign micromatrizz[44][305] = 9'b111111111;
assign micromatrizz[44][306] = 9'b111111111;
assign micromatrizz[44][307] = 9'b111111111;
assign micromatrizz[44][308] = 9'b111111111;
assign micromatrizz[44][309] = 9'b111111111;
assign micromatrizz[44][310] = 9'b111111111;
assign micromatrizz[44][311] = 9'b111111111;
assign micromatrizz[44][312] = 9'b111111111;
assign micromatrizz[44][313] = 9'b111111111;
assign micromatrizz[44][314] = 9'b111111111;
assign micromatrizz[44][315] = 9'b111111111;
assign micromatrizz[44][316] = 9'b111111111;
assign micromatrizz[44][317] = 9'b111111111;
assign micromatrizz[44][318] = 9'b111111111;
assign micromatrizz[44][319] = 9'b111111111;
assign micromatrizz[44][320] = 9'b111111111;
assign micromatrizz[44][321] = 9'b111111111;
assign micromatrizz[44][322] = 9'b111111111;
assign micromatrizz[44][323] = 9'b111111111;
assign micromatrizz[44][324] = 9'b111111111;
assign micromatrizz[44][325] = 9'b111111111;
assign micromatrizz[44][326] = 9'b111111111;
assign micromatrizz[44][327] = 9'b111111111;
assign micromatrizz[44][328] = 9'b111111111;
assign micromatrizz[44][329] = 9'b111111111;
assign micromatrizz[44][330] = 9'b111111111;
assign micromatrizz[44][331] = 9'b111111111;
assign micromatrizz[44][332] = 9'b111111111;
assign micromatrizz[44][333] = 9'b111111111;
assign micromatrizz[44][334] = 9'b111111111;
assign micromatrizz[44][335] = 9'b111111111;
assign micromatrizz[44][336] = 9'b111111111;
assign micromatrizz[44][337] = 9'b111111111;
assign micromatrizz[44][338] = 9'b111111111;
assign micromatrizz[44][339] = 9'b111111111;
assign micromatrizz[44][340] = 9'b111111111;
assign micromatrizz[44][341] = 9'b111111111;
assign micromatrizz[44][342] = 9'b111111111;
assign micromatrizz[44][343] = 9'b111111111;
assign micromatrizz[44][344] = 9'b111111111;
assign micromatrizz[44][345] = 9'b111111111;
assign micromatrizz[44][346] = 9'b111111111;
assign micromatrizz[44][347] = 9'b111111111;
assign micromatrizz[44][348] = 9'b111111111;
assign micromatrizz[44][349] = 9'b111111111;
assign micromatrizz[44][350] = 9'b111111111;
assign micromatrizz[44][351] = 9'b111111111;
assign micromatrizz[44][352] = 9'b111111111;
assign micromatrizz[44][353] = 9'b111111111;
assign micromatrizz[44][354] = 9'b111111111;
assign micromatrizz[44][355] = 9'b111111111;
assign micromatrizz[44][356] = 9'b111111111;
assign micromatrizz[44][357] = 9'b111111111;
assign micromatrizz[44][358] = 9'b111111111;
assign micromatrizz[44][359] = 9'b111111111;
assign micromatrizz[44][360] = 9'b111111111;
assign micromatrizz[44][361] = 9'b111111111;
assign micromatrizz[44][362] = 9'b111111111;
assign micromatrizz[44][363] = 9'b111111111;
assign micromatrizz[44][364] = 9'b111111111;
assign micromatrizz[44][365] = 9'b111111111;
assign micromatrizz[44][366] = 9'b111111111;
assign micromatrizz[44][367] = 9'b111111111;
assign micromatrizz[44][368] = 9'b111111111;
assign micromatrizz[44][369] = 9'b111111111;
assign micromatrizz[44][370] = 9'b111111111;
assign micromatrizz[44][371] = 9'b111111111;
assign micromatrizz[44][372] = 9'b111111111;
assign micromatrizz[44][373] = 9'b111111111;
assign micromatrizz[44][374] = 9'b111111111;
assign micromatrizz[44][375] = 9'b111111111;
assign micromatrizz[44][376] = 9'b111111111;
assign micromatrizz[44][377] = 9'b111111111;
assign micromatrizz[44][378] = 9'b111111111;
assign micromatrizz[44][379] = 9'b111111111;
assign micromatrizz[44][380] = 9'b111111111;
assign micromatrizz[44][381] = 9'b111111111;
assign micromatrizz[44][382] = 9'b111111111;
assign micromatrizz[44][383] = 9'b111111111;
assign micromatrizz[44][384] = 9'b111111111;
assign micromatrizz[44][385] = 9'b111111111;
assign micromatrizz[44][386] = 9'b111111111;
assign micromatrizz[44][387] = 9'b111111111;
assign micromatrizz[44][388] = 9'b111111111;
assign micromatrizz[44][389] = 9'b111111111;
assign micromatrizz[44][390] = 9'b111111111;
assign micromatrizz[44][391] = 9'b111111111;
assign micromatrizz[44][392] = 9'b111111111;
assign micromatrizz[44][393] = 9'b111111111;
assign micromatrizz[44][394] = 9'b111111111;
assign micromatrizz[44][395] = 9'b111111111;
assign micromatrizz[44][396] = 9'b111111111;
assign micromatrizz[44][397] = 9'b111111111;
assign micromatrizz[44][398] = 9'b111111111;
assign micromatrizz[44][399] = 9'b111111111;
assign micromatrizz[44][400] = 9'b111111111;
assign micromatrizz[44][401] = 9'b111111111;
assign micromatrizz[44][402] = 9'b111111111;
assign micromatrizz[44][403] = 9'b111111111;
assign micromatrizz[44][404] = 9'b111111111;
assign micromatrizz[44][405] = 9'b111111111;
assign micromatrizz[44][406] = 9'b111111111;
assign micromatrizz[44][407] = 9'b111111111;
assign micromatrizz[44][408] = 9'b111111111;
assign micromatrizz[44][409] = 9'b111111111;
assign micromatrizz[44][410] = 9'b111111111;
assign micromatrizz[44][411] = 9'b111111111;
assign micromatrizz[44][412] = 9'b111111111;
assign micromatrizz[44][413] = 9'b111111111;
assign micromatrizz[44][414] = 9'b111111111;
assign micromatrizz[44][415] = 9'b111111111;
assign micromatrizz[44][416] = 9'b111111111;
assign micromatrizz[44][417] = 9'b111111111;
assign micromatrizz[44][418] = 9'b111111111;
assign micromatrizz[44][419] = 9'b111111111;
assign micromatrizz[44][420] = 9'b111111111;
assign micromatrizz[44][421] = 9'b111111111;
assign micromatrizz[44][422] = 9'b111111111;
assign micromatrizz[44][423] = 9'b111111111;
assign micromatrizz[44][424] = 9'b111111111;
assign micromatrizz[44][425] = 9'b111111111;
assign micromatrizz[44][426] = 9'b111111111;
assign micromatrizz[44][427] = 9'b111111111;
assign micromatrizz[44][428] = 9'b111111111;
assign micromatrizz[44][429] = 9'b111111111;
assign micromatrizz[44][430] = 9'b111111111;
assign micromatrizz[44][431] = 9'b111111111;
assign micromatrizz[44][432] = 9'b111111111;
assign micromatrizz[44][433] = 9'b111111111;
assign micromatrizz[44][434] = 9'b111111111;
assign micromatrizz[44][435] = 9'b111111111;
assign micromatrizz[44][436] = 9'b111111111;
assign micromatrizz[44][437] = 9'b111111111;
assign micromatrizz[44][438] = 9'b111111111;
assign micromatrizz[44][439] = 9'b111111111;
assign micromatrizz[44][440] = 9'b111111111;
assign micromatrizz[44][441] = 9'b111111111;
assign micromatrizz[44][442] = 9'b111111111;
assign micromatrizz[44][443] = 9'b111111111;
assign micromatrizz[44][444] = 9'b111111111;
assign micromatrizz[44][445] = 9'b111111111;
assign micromatrizz[44][446] = 9'b111111111;
assign micromatrizz[44][447] = 9'b111111111;
assign micromatrizz[44][448] = 9'b111111111;
assign micromatrizz[44][449] = 9'b111111111;
assign micromatrizz[44][450] = 9'b111111111;
assign micromatrizz[44][451] = 9'b111111111;
assign micromatrizz[44][452] = 9'b111111111;
assign micromatrizz[44][453] = 9'b111111111;
assign micromatrizz[44][454] = 9'b111111111;
assign micromatrizz[44][455] = 9'b111111111;
assign micromatrizz[44][456] = 9'b111111111;
assign micromatrizz[44][457] = 9'b111111111;
assign micromatrizz[44][458] = 9'b111111111;
assign micromatrizz[44][459] = 9'b111111111;
assign micromatrizz[44][460] = 9'b111111111;
assign micromatrizz[44][461] = 9'b111111111;
assign micromatrizz[44][462] = 9'b111111111;
assign micromatrizz[44][463] = 9'b111111111;
assign micromatrizz[44][464] = 9'b111111111;
assign micromatrizz[44][465] = 9'b111111111;
assign micromatrizz[44][466] = 9'b111111111;
assign micromatrizz[44][467] = 9'b111111111;
assign micromatrizz[44][468] = 9'b111111111;
assign micromatrizz[44][469] = 9'b111111111;
assign micromatrizz[44][470] = 9'b111111111;
assign micromatrizz[44][471] = 9'b111111111;
assign micromatrizz[44][472] = 9'b111111111;
assign micromatrizz[44][473] = 9'b111111111;
assign micromatrizz[44][474] = 9'b111111111;
assign micromatrizz[44][475] = 9'b111111111;
assign micromatrizz[44][476] = 9'b111111111;
assign micromatrizz[44][477] = 9'b111111111;
assign micromatrizz[44][478] = 9'b111111111;
assign micromatrizz[44][479] = 9'b111111111;
assign micromatrizz[44][480] = 9'b111111111;
assign micromatrizz[44][481] = 9'b111111111;
assign micromatrizz[44][482] = 9'b111111111;
assign micromatrizz[44][483] = 9'b111111111;
assign micromatrizz[44][484] = 9'b111111111;
assign micromatrizz[44][485] = 9'b111111111;
assign micromatrizz[44][486] = 9'b111111111;
assign micromatrizz[44][487] = 9'b111111111;
assign micromatrizz[44][488] = 9'b111111111;
assign micromatrizz[44][489] = 9'b111111111;
assign micromatrizz[44][490] = 9'b111111111;
assign micromatrizz[44][491] = 9'b111111111;
assign micromatrizz[44][492] = 9'b111111111;
assign micromatrizz[44][493] = 9'b111111111;
assign micromatrizz[44][494] = 9'b111111111;
assign micromatrizz[44][495] = 9'b111111111;
assign micromatrizz[44][496] = 9'b111111111;
assign micromatrizz[44][497] = 9'b111111111;
assign micromatrizz[44][498] = 9'b111111111;
assign micromatrizz[44][499] = 9'b111111111;
assign micromatrizz[44][500] = 9'b111111111;
assign micromatrizz[44][501] = 9'b111111111;
assign micromatrizz[44][502] = 9'b111111111;
assign micromatrizz[44][503] = 9'b111111111;
assign micromatrizz[44][504] = 9'b111111111;
assign micromatrizz[44][505] = 9'b111111111;
assign micromatrizz[44][506] = 9'b111111111;
assign micromatrizz[44][507] = 9'b111111111;
assign micromatrizz[44][508] = 9'b111111111;
assign micromatrizz[44][509] = 9'b111111111;
assign micromatrizz[44][510] = 9'b111111111;
assign micromatrizz[44][511] = 9'b111111111;
assign micromatrizz[44][512] = 9'b111111111;
assign micromatrizz[44][513] = 9'b111111111;
assign micromatrizz[44][514] = 9'b111111111;
assign micromatrizz[44][515] = 9'b111111111;
assign micromatrizz[44][516] = 9'b111111111;
assign micromatrizz[44][517] = 9'b111111111;
assign micromatrizz[44][518] = 9'b111111111;
assign micromatrizz[44][519] = 9'b111111111;
assign micromatrizz[44][520] = 9'b111111111;
assign micromatrizz[44][521] = 9'b111111111;
assign micromatrizz[44][522] = 9'b111111111;
assign micromatrizz[44][523] = 9'b111111111;
assign micromatrizz[44][524] = 9'b111111111;
assign micromatrizz[44][525] = 9'b111111111;
assign micromatrizz[44][526] = 9'b111111111;
assign micromatrizz[44][527] = 9'b111111111;
assign micromatrizz[44][528] = 9'b111111111;
assign micromatrizz[44][529] = 9'b111111111;
assign micromatrizz[44][530] = 9'b111111111;
assign micromatrizz[44][531] = 9'b111111111;
assign micromatrizz[44][532] = 9'b111111111;
assign micromatrizz[44][533] = 9'b111111111;
assign micromatrizz[44][534] = 9'b111111111;
assign micromatrizz[44][535] = 9'b111111111;
assign micromatrizz[44][536] = 9'b111111111;
assign micromatrizz[44][537] = 9'b111111111;
assign micromatrizz[44][538] = 9'b111111111;
assign micromatrizz[44][539] = 9'b111111111;
assign micromatrizz[44][540] = 9'b111111111;
assign micromatrizz[44][541] = 9'b111111111;
assign micromatrizz[44][542] = 9'b111111111;
assign micromatrizz[44][543] = 9'b111111111;
assign micromatrizz[44][544] = 9'b111111111;
assign micromatrizz[44][545] = 9'b111111111;
assign micromatrizz[44][546] = 9'b111111111;
assign micromatrizz[44][547] = 9'b111111111;
assign micromatrizz[44][548] = 9'b111111111;
assign micromatrizz[44][549] = 9'b111111111;
assign micromatrizz[44][550] = 9'b111111111;
assign micromatrizz[44][551] = 9'b111111111;
assign micromatrizz[44][552] = 9'b111111111;
assign micromatrizz[44][553] = 9'b111111111;
assign micromatrizz[44][554] = 9'b111111111;
assign micromatrizz[44][555] = 9'b111111111;
assign micromatrizz[44][556] = 9'b111111111;
assign micromatrizz[44][557] = 9'b111111111;
assign micromatrizz[44][558] = 9'b111111111;
assign micromatrizz[44][559] = 9'b111111111;
assign micromatrizz[44][560] = 9'b111111111;
assign micromatrizz[44][561] = 9'b111111111;
assign micromatrizz[44][562] = 9'b111111111;
assign micromatrizz[44][563] = 9'b111111111;
assign micromatrizz[44][564] = 9'b111111111;
assign micromatrizz[44][565] = 9'b111111111;
assign micromatrizz[44][566] = 9'b111111111;
assign micromatrizz[44][567] = 9'b111111111;
assign micromatrizz[44][568] = 9'b111111111;
assign micromatrizz[44][569] = 9'b111111111;
assign micromatrizz[44][570] = 9'b111111111;
assign micromatrizz[44][571] = 9'b111111111;
assign micromatrizz[44][572] = 9'b111111111;
assign micromatrizz[44][573] = 9'b111111111;
assign micromatrizz[44][574] = 9'b111111111;
assign micromatrizz[44][575] = 9'b111111111;
assign micromatrizz[44][576] = 9'b111111111;
assign micromatrizz[44][577] = 9'b111111111;
assign micromatrizz[44][578] = 9'b111111111;
assign micromatrizz[44][579] = 9'b111111111;
assign micromatrizz[44][580] = 9'b111111111;
assign micromatrizz[44][581] = 9'b111111111;
assign micromatrizz[44][582] = 9'b111111111;
assign micromatrizz[44][583] = 9'b111111111;
assign micromatrizz[44][584] = 9'b111111111;
assign micromatrizz[44][585] = 9'b111111111;
assign micromatrizz[44][586] = 9'b111111111;
assign micromatrizz[44][587] = 9'b111111111;
assign micromatrizz[44][588] = 9'b111111111;
assign micromatrizz[44][589] = 9'b111111111;
assign micromatrizz[44][590] = 9'b111111111;
assign micromatrizz[44][591] = 9'b111111111;
assign micromatrizz[44][592] = 9'b111111111;
assign micromatrizz[44][593] = 9'b111111111;
assign micromatrizz[44][594] = 9'b111111111;
assign micromatrizz[44][595] = 9'b111111111;
assign micromatrizz[44][596] = 9'b111111111;
assign micromatrizz[44][597] = 9'b111111111;
assign micromatrizz[44][598] = 9'b111111111;
assign micromatrizz[44][599] = 9'b111111111;
assign micromatrizz[44][600] = 9'b111111111;
assign micromatrizz[44][601] = 9'b111111111;
assign micromatrizz[44][602] = 9'b111111111;
assign micromatrizz[44][603] = 9'b111111111;
assign micromatrizz[44][604] = 9'b111111111;
assign micromatrizz[44][605] = 9'b111111111;
assign micromatrizz[44][606] = 9'b111111111;
assign micromatrizz[44][607] = 9'b111111111;
assign micromatrizz[44][608] = 9'b111111111;
assign micromatrizz[44][609] = 9'b111111111;
assign micromatrizz[44][610] = 9'b111111111;
assign micromatrizz[44][611] = 9'b111111111;
assign micromatrizz[44][612] = 9'b111111111;
assign micromatrizz[44][613] = 9'b111111111;
assign micromatrizz[44][614] = 9'b111111111;
assign micromatrizz[44][615] = 9'b111111111;
assign micromatrizz[44][616] = 9'b111111111;
assign micromatrizz[44][617] = 9'b111111111;
assign micromatrizz[44][618] = 9'b111111111;
assign micromatrizz[44][619] = 9'b111111111;
assign micromatrizz[44][620] = 9'b111111111;
assign micromatrizz[44][621] = 9'b111111111;
assign micromatrizz[44][622] = 9'b111111111;
assign micromatrizz[44][623] = 9'b111111111;
assign micromatrizz[44][624] = 9'b111111111;
assign micromatrizz[44][625] = 9'b111111111;
assign micromatrizz[44][626] = 9'b111111111;
assign micromatrizz[44][627] = 9'b111111111;
assign micromatrizz[44][628] = 9'b111111111;
assign micromatrizz[44][629] = 9'b111111111;
assign micromatrizz[44][630] = 9'b111111111;
assign micromatrizz[44][631] = 9'b111111111;
assign micromatrizz[44][632] = 9'b111111111;
assign micromatrizz[44][633] = 9'b111111111;
assign micromatrizz[44][634] = 9'b111111111;
assign micromatrizz[44][635] = 9'b111111111;
assign micromatrizz[44][636] = 9'b111111111;
assign micromatrizz[44][637] = 9'b111111111;
assign micromatrizz[44][638] = 9'b111111111;
assign micromatrizz[44][639] = 9'b111111111;
assign micromatrizz[45][0] = 9'b111111111;
assign micromatrizz[45][1] = 9'b111111111;
assign micromatrizz[45][2] = 9'b111111111;
assign micromatrizz[45][3] = 9'b111111111;
assign micromatrizz[45][4] = 9'b111111111;
assign micromatrizz[45][5] = 9'b111111111;
assign micromatrizz[45][6] = 9'b111111111;
assign micromatrizz[45][7] = 9'b111111111;
assign micromatrizz[45][8] = 9'b111111111;
assign micromatrizz[45][9] = 9'b111111111;
assign micromatrizz[45][10] = 9'b111111111;
assign micromatrizz[45][11] = 9'b111111111;
assign micromatrizz[45][12] = 9'b111111111;
assign micromatrizz[45][13] = 9'b111111111;
assign micromatrizz[45][14] = 9'b111111111;
assign micromatrizz[45][15] = 9'b111111111;
assign micromatrizz[45][16] = 9'b111111111;
assign micromatrizz[45][17] = 9'b111111111;
assign micromatrizz[45][18] = 9'b111111111;
assign micromatrizz[45][19] = 9'b111111111;
assign micromatrizz[45][20] = 9'b111111111;
assign micromatrizz[45][21] = 9'b111111111;
assign micromatrizz[45][22] = 9'b111111111;
assign micromatrizz[45][23] = 9'b111111111;
assign micromatrizz[45][24] = 9'b111111111;
assign micromatrizz[45][25] = 9'b111111111;
assign micromatrizz[45][26] = 9'b111111111;
assign micromatrizz[45][27] = 9'b111111111;
assign micromatrizz[45][28] = 9'b111111111;
assign micromatrizz[45][29] = 9'b111111111;
assign micromatrizz[45][30] = 9'b111111111;
assign micromatrizz[45][31] = 9'b111111111;
assign micromatrizz[45][32] = 9'b111111111;
assign micromatrizz[45][33] = 9'b111111111;
assign micromatrizz[45][34] = 9'b111111111;
assign micromatrizz[45][35] = 9'b111111111;
assign micromatrizz[45][36] = 9'b111111111;
assign micromatrizz[45][37] = 9'b111111111;
assign micromatrizz[45][38] = 9'b111111111;
assign micromatrizz[45][39] = 9'b111111111;
assign micromatrizz[45][40] = 9'b111111111;
assign micromatrizz[45][41] = 9'b111111111;
assign micromatrizz[45][42] = 9'b111111111;
assign micromatrizz[45][43] = 9'b111111111;
assign micromatrizz[45][44] = 9'b111111111;
assign micromatrizz[45][45] = 9'b111111111;
assign micromatrizz[45][46] = 9'b111111111;
assign micromatrizz[45][47] = 9'b111111111;
assign micromatrizz[45][48] = 9'b111111111;
assign micromatrizz[45][49] = 9'b111111111;
assign micromatrizz[45][50] = 9'b111111111;
assign micromatrizz[45][51] = 9'b111111111;
assign micromatrizz[45][52] = 9'b111111111;
assign micromatrizz[45][53] = 9'b111111111;
assign micromatrizz[45][54] = 9'b111111111;
assign micromatrizz[45][55] = 9'b111111111;
assign micromatrizz[45][56] = 9'b111111111;
assign micromatrizz[45][57] = 9'b111111111;
assign micromatrizz[45][58] = 9'b111111111;
assign micromatrizz[45][59] = 9'b111111111;
assign micromatrizz[45][60] = 9'b111111111;
assign micromatrizz[45][61] = 9'b111111111;
assign micromatrizz[45][62] = 9'b111111111;
assign micromatrizz[45][63] = 9'b111111111;
assign micromatrizz[45][64] = 9'b111111111;
assign micromatrizz[45][65] = 9'b111111111;
assign micromatrizz[45][66] = 9'b111111111;
assign micromatrizz[45][67] = 9'b111111111;
assign micromatrizz[45][68] = 9'b111111111;
assign micromatrizz[45][69] = 9'b111111111;
assign micromatrizz[45][70] = 9'b111111111;
assign micromatrizz[45][71] = 9'b111111111;
assign micromatrizz[45][72] = 9'b111111111;
assign micromatrizz[45][73] = 9'b111111111;
assign micromatrizz[45][74] = 9'b111111111;
assign micromatrizz[45][75] = 9'b111111111;
assign micromatrizz[45][76] = 9'b111111111;
assign micromatrizz[45][77] = 9'b111111111;
assign micromatrizz[45][78] = 9'b111111111;
assign micromatrizz[45][79] = 9'b111111111;
assign micromatrizz[45][80] = 9'b111111111;
assign micromatrizz[45][81] = 9'b111111111;
assign micromatrizz[45][82] = 9'b111111111;
assign micromatrizz[45][83] = 9'b111111111;
assign micromatrizz[45][84] = 9'b111111111;
assign micromatrizz[45][85] = 9'b111111111;
assign micromatrizz[45][86] = 9'b111111111;
assign micromatrizz[45][87] = 9'b111111111;
assign micromatrizz[45][88] = 9'b111111111;
assign micromatrizz[45][89] = 9'b111111111;
assign micromatrizz[45][90] = 9'b111111111;
assign micromatrizz[45][91] = 9'b111111111;
assign micromatrizz[45][92] = 9'b111111111;
assign micromatrizz[45][93] = 9'b111111111;
assign micromatrizz[45][94] = 9'b111111111;
assign micromatrizz[45][95] = 9'b111111111;
assign micromatrizz[45][96] = 9'b111111111;
assign micromatrizz[45][97] = 9'b111111111;
assign micromatrizz[45][98] = 9'b111111111;
assign micromatrizz[45][99] = 9'b111111111;
assign micromatrizz[45][100] = 9'b111111111;
assign micromatrizz[45][101] = 9'b111111111;
assign micromatrizz[45][102] = 9'b111111111;
assign micromatrizz[45][103] = 9'b111111111;
assign micromatrizz[45][104] = 9'b111111111;
assign micromatrizz[45][105] = 9'b111111111;
assign micromatrizz[45][106] = 9'b111111111;
assign micromatrizz[45][107] = 9'b111111111;
assign micromatrizz[45][108] = 9'b111111111;
assign micromatrizz[45][109] = 9'b111111111;
assign micromatrizz[45][110] = 9'b111111111;
assign micromatrizz[45][111] = 9'b111111111;
assign micromatrizz[45][112] = 9'b111111111;
assign micromatrizz[45][113] = 9'b111111111;
assign micromatrizz[45][114] = 9'b111111111;
assign micromatrizz[45][115] = 9'b111111111;
assign micromatrizz[45][116] = 9'b111111111;
assign micromatrizz[45][117] = 9'b111111111;
assign micromatrizz[45][118] = 9'b111111111;
assign micromatrizz[45][119] = 9'b111111111;
assign micromatrizz[45][120] = 9'b111111111;
assign micromatrizz[45][121] = 9'b111111111;
assign micromatrizz[45][122] = 9'b111111111;
assign micromatrizz[45][123] = 9'b111111111;
assign micromatrizz[45][124] = 9'b111111111;
assign micromatrizz[45][125] = 9'b111111111;
assign micromatrizz[45][126] = 9'b111111111;
assign micromatrizz[45][127] = 9'b111111111;
assign micromatrizz[45][128] = 9'b111111111;
assign micromatrizz[45][129] = 9'b111111111;
assign micromatrizz[45][130] = 9'b111111111;
assign micromatrizz[45][131] = 9'b111111111;
assign micromatrizz[45][132] = 9'b111111111;
assign micromatrizz[45][133] = 9'b111111111;
assign micromatrizz[45][134] = 9'b111111111;
assign micromatrizz[45][135] = 9'b111111111;
assign micromatrizz[45][136] = 9'b111111111;
assign micromatrizz[45][137] = 9'b111111111;
assign micromatrizz[45][138] = 9'b111111111;
assign micromatrizz[45][139] = 9'b111111111;
assign micromatrizz[45][140] = 9'b111111111;
assign micromatrizz[45][141] = 9'b111111111;
assign micromatrizz[45][142] = 9'b111111111;
assign micromatrizz[45][143] = 9'b111111111;
assign micromatrizz[45][144] = 9'b111111111;
assign micromatrizz[45][145] = 9'b111111111;
assign micromatrizz[45][146] = 9'b111110111;
assign micromatrizz[45][147] = 9'b111110010;
assign micromatrizz[45][148] = 9'b111110011;
assign micromatrizz[45][149] = 9'b111110111;
assign micromatrizz[45][150] = 9'b111111111;
assign micromatrizz[45][151] = 9'b111111111;
assign micromatrizz[45][152] = 9'b111111111;
assign micromatrizz[45][153] = 9'b111111111;
assign micromatrizz[45][154] = 9'b111110010;
assign micromatrizz[45][155] = 9'b111111111;
assign micromatrizz[45][156] = 9'b111111111;
assign micromatrizz[45][157] = 9'b111111111;
assign micromatrizz[45][158] = 9'b111111111;
assign micromatrizz[45][159] = 9'b111111111;
assign micromatrizz[45][160] = 9'b111111111;
assign micromatrizz[45][161] = 9'b111111111;
assign micromatrizz[45][162] = 9'b111111111;
assign micromatrizz[45][163] = 9'b111111111;
assign micromatrizz[45][164] = 9'b111111111;
assign micromatrizz[45][165] = 9'b111111111;
assign micromatrizz[45][166] = 9'b111111111;
assign micromatrizz[45][167] = 9'b111111111;
assign micromatrizz[45][168] = 9'b111111111;
assign micromatrizz[45][169] = 9'b111111111;
assign micromatrizz[45][170] = 9'b111111111;
assign micromatrizz[45][171] = 9'b111111111;
assign micromatrizz[45][172] = 9'b111111111;
assign micromatrizz[45][173] = 9'b111111111;
assign micromatrizz[45][174] = 9'b111111111;
assign micromatrizz[45][175] = 9'b111111111;
assign micromatrizz[45][176] = 9'b111111111;
assign micromatrizz[45][177] = 9'b111111111;
assign micromatrizz[45][178] = 9'b111111111;
assign micromatrizz[45][179] = 9'b111111111;
assign micromatrizz[45][180] = 9'b111111111;
assign micromatrizz[45][181] = 9'b111111111;
assign micromatrizz[45][182] = 9'b111111111;
assign micromatrizz[45][183] = 9'b111111111;
assign micromatrizz[45][184] = 9'b111111111;
assign micromatrizz[45][185] = 9'b111111111;
assign micromatrizz[45][186] = 9'b111111111;
assign micromatrizz[45][187] = 9'b111111111;
assign micromatrizz[45][188] = 9'b111111111;
assign micromatrizz[45][189] = 9'b111111111;
assign micromatrizz[45][190] = 9'b111111111;
assign micromatrizz[45][191] = 9'b111111111;
assign micromatrizz[45][192] = 9'b111111111;
assign micromatrizz[45][193] = 9'b111111111;
assign micromatrizz[45][194] = 9'b111111111;
assign micromatrizz[45][195] = 9'b111111111;
assign micromatrizz[45][196] = 9'b111111111;
assign micromatrizz[45][197] = 9'b111111111;
assign micromatrizz[45][198] = 9'b111111111;
assign micromatrizz[45][199] = 9'b111111111;
assign micromatrizz[45][200] = 9'b111111111;
assign micromatrizz[45][201] = 9'b111111111;
assign micromatrizz[45][202] = 9'b111111111;
assign micromatrizz[45][203] = 9'b111111111;
assign micromatrizz[45][204] = 9'b111111111;
assign micromatrizz[45][205] = 9'b111111111;
assign micromatrizz[45][206] = 9'b111111111;
assign micromatrizz[45][207] = 9'b111111111;
assign micromatrizz[45][208] = 9'b111111111;
assign micromatrizz[45][209] = 9'b111111111;
assign micromatrizz[45][210] = 9'b111111111;
assign micromatrizz[45][211] = 9'b111111111;
assign micromatrizz[45][212] = 9'b111111111;
assign micromatrizz[45][213] = 9'b111111111;
assign micromatrizz[45][214] = 9'b111111111;
assign micromatrizz[45][215] = 9'b111111111;
assign micromatrizz[45][216] = 9'b111111111;
assign micromatrizz[45][217] = 9'b111111111;
assign micromatrizz[45][218] = 9'b111111111;
assign micromatrizz[45][219] = 9'b111111111;
assign micromatrizz[45][220] = 9'b111111111;
assign micromatrizz[45][221] = 9'b111111111;
assign micromatrizz[45][222] = 9'b111111111;
assign micromatrizz[45][223] = 9'b111111111;
assign micromatrizz[45][224] = 9'b111111111;
assign micromatrizz[45][225] = 9'b111111111;
assign micromatrizz[45][226] = 9'b111111111;
assign micromatrizz[45][227] = 9'b111111111;
assign micromatrizz[45][228] = 9'b111111111;
assign micromatrizz[45][229] = 9'b111111111;
assign micromatrizz[45][230] = 9'b111111111;
assign micromatrizz[45][231] = 9'b111111111;
assign micromatrizz[45][232] = 9'b111111111;
assign micromatrizz[45][233] = 9'b111111111;
assign micromatrizz[45][234] = 9'b111111111;
assign micromatrizz[45][235] = 9'b111111111;
assign micromatrizz[45][236] = 9'b111111111;
assign micromatrizz[45][237] = 9'b111111111;
assign micromatrizz[45][238] = 9'b111111111;
assign micromatrizz[45][239] = 9'b111111111;
assign micromatrizz[45][240] = 9'b111111111;
assign micromatrizz[45][241] = 9'b111111111;
assign micromatrizz[45][242] = 9'b111111111;
assign micromatrizz[45][243] = 9'b111111111;
assign micromatrizz[45][244] = 9'b111111111;
assign micromatrizz[45][245] = 9'b111111111;
assign micromatrizz[45][246] = 9'b111111111;
assign micromatrizz[45][247] = 9'b111111111;
assign micromatrizz[45][248] = 9'b111111111;
assign micromatrizz[45][249] = 9'b111111111;
assign micromatrizz[45][250] = 9'b111111111;
assign micromatrizz[45][251] = 9'b111111111;
assign micromatrizz[45][252] = 9'b111111111;
assign micromatrizz[45][253] = 9'b111111111;
assign micromatrizz[45][254] = 9'b111111111;
assign micromatrizz[45][255] = 9'b111111111;
assign micromatrizz[45][256] = 9'b111111111;
assign micromatrizz[45][257] = 9'b111111111;
assign micromatrizz[45][258] = 9'b111111111;
assign micromatrizz[45][259] = 9'b111111111;
assign micromatrizz[45][260] = 9'b111111111;
assign micromatrizz[45][261] = 9'b111111111;
assign micromatrizz[45][262] = 9'b111111111;
assign micromatrizz[45][263] = 9'b111111111;
assign micromatrizz[45][264] = 9'b111111111;
assign micromatrizz[45][265] = 9'b111111111;
assign micromatrizz[45][266] = 9'b111111111;
assign micromatrizz[45][267] = 9'b111111111;
assign micromatrizz[45][268] = 9'b111111111;
assign micromatrizz[45][269] = 9'b111111111;
assign micromatrizz[45][270] = 9'b111111111;
assign micromatrizz[45][271] = 9'b111111111;
assign micromatrizz[45][272] = 9'b111111111;
assign micromatrizz[45][273] = 9'b111111111;
assign micromatrizz[45][274] = 9'b111111111;
assign micromatrizz[45][275] = 9'b111111111;
assign micromatrizz[45][276] = 9'b111111111;
assign micromatrizz[45][277] = 9'b111111111;
assign micromatrizz[45][278] = 9'b111111111;
assign micromatrizz[45][279] = 9'b111111111;
assign micromatrizz[45][280] = 9'b111111111;
assign micromatrizz[45][281] = 9'b111111111;
assign micromatrizz[45][282] = 9'b111111111;
assign micromatrizz[45][283] = 9'b111111111;
assign micromatrizz[45][284] = 9'b111111111;
assign micromatrizz[45][285] = 9'b111111111;
assign micromatrizz[45][286] = 9'b111111111;
assign micromatrizz[45][287] = 9'b111111111;
assign micromatrizz[45][288] = 9'b111111111;
assign micromatrizz[45][289] = 9'b111111111;
assign micromatrizz[45][290] = 9'b111111111;
assign micromatrizz[45][291] = 9'b111111111;
assign micromatrizz[45][292] = 9'b111111111;
assign micromatrizz[45][293] = 9'b111111111;
assign micromatrizz[45][294] = 9'b111111111;
assign micromatrizz[45][295] = 9'b111111111;
assign micromatrizz[45][296] = 9'b111111111;
assign micromatrizz[45][297] = 9'b111111111;
assign micromatrizz[45][298] = 9'b111111111;
assign micromatrizz[45][299] = 9'b111111111;
assign micromatrizz[45][300] = 9'b111111111;
assign micromatrizz[45][301] = 9'b111111111;
assign micromatrizz[45][302] = 9'b111111111;
assign micromatrizz[45][303] = 9'b111111111;
assign micromatrizz[45][304] = 9'b111111111;
assign micromatrizz[45][305] = 9'b111111111;
assign micromatrizz[45][306] = 9'b111111111;
assign micromatrizz[45][307] = 9'b111111111;
assign micromatrizz[45][308] = 9'b111111111;
assign micromatrizz[45][309] = 9'b111111111;
assign micromatrizz[45][310] = 9'b111111111;
assign micromatrizz[45][311] = 9'b111111111;
assign micromatrizz[45][312] = 9'b111111111;
assign micromatrizz[45][313] = 9'b111111111;
assign micromatrizz[45][314] = 9'b111111111;
assign micromatrizz[45][315] = 9'b111111111;
assign micromatrizz[45][316] = 9'b111111111;
assign micromatrizz[45][317] = 9'b111111111;
assign micromatrizz[45][318] = 9'b111111111;
assign micromatrizz[45][319] = 9'b111111111;
assign micromatrizz[45][320] = 9'b111111111;
assign micromatrizz[45][321] = 9'b111111111;
assign micromatrizz[45][322] = 9'b111111111;
assign micromatrizz[45][323] = 9'b111111111;
assign micromatrizz[45][324] = 9'b111111111;
assign micromatrizz[45][325] = 9'b111111111;
assign micromatrizz[45][326] = 9'b111111111;
assign micromatrizz[45][327] = 9'b111111111;
assign micromatrizz[45][328] = 9'b111111111;
assign micromatrizz[45][329] = 9'b111111111;
assign micromatrizz[45][330] = 9'b111111111;
assign micromatrizz[45][331] = 9'b111111111;
assign micromatrizz[45][332] = 9'b111111111;
assign micromatrizz[45][333] = 9'b111111111;
assign micromatrizz[45][334] = 9'b111111111;
assign micromatrizz[45][335] = 9'b111111111;
assign micromatrizz[45][336] = 9'b111111111;
assign micromatrizz[45][337] = 9'b111111111;
assign micromatrizz[45][338] = 9'b111111111;
assign micromatrizz[45][339] = 9'b111111111;
assign micromatrizz[45][340] = 9'b111111111;
assign micromatrizz[45][341] = 9'b111111111;
assign micromatrizz[45][342] = 9'b111111111;
assign micromatrizz[45][343] = 9'b111111111;
assign micromatrizz[45][344] = 9'b111111111;
assign micromatrizz[45][345] = 9'b111111111;
assign micromatrizz[45][346] = 9'b111111111;
assign micromatrizz[45][347] = 9'b111111111;
assign micromatrizz[45][348] = 9'b111111111;
assign micromatrizz[45][349] = 9'b111111111;
assign micromatrizz[45][350] = 9'b111111111;
assign micromatrizz[45][351] = 9'b111111111;
assign micromatrizz[45][352] = 9'b111111111;
assign micromatrizz[45][353] = 9'b111111111;
assign micromatrizz[45][354] = 9'b111111111;
assign micromatrizz[45][355] = 9'b111111111;
assign micromatrizz[45][356] = 9'b111111111;
assign micromatrizz[45][357] = 9'b111111111;
assign micromatrizz[45][358] = 9'b111111111;
assign micromatrizz[45][359] = 9'b111111111;
assign micromatrizz[45][360] = 9'b111111111;
assign micromatrizz[45][361] = 9'b111111111;
assign micromatrizz[45][362] = 9'b111111111;
assign micromatrizz[45][363] = 9'b111111111;
assign micromatrizz[45][364] = 9'b111111111;
assign micromatrizz[45][365] = 9'b111111111;
assign micromatrizz[45][366] = 9'b111111111;
assign micromatrizz[45][367] = 9'b111111111;
assign micromatrizz[45][368] = 9'b111111111;
assign micromatrizz[45][369] = 9'b111111111;
assign micromatrizz[45][370] = 9'b111111111;
assign micromatrizz[45][371] = 9'b111111111;
assign micromatrizz[45][372] = 9'b111111111;
assign micromatrizz[45][373] = 9'b111111111;
assign micromatrizz[45][374] = 9'b111111111;
assign micromatrizz[45][375] = 9'b111111111;
assign micromatrizz[45][376] = 9'b111111111;
assign micromatrizz[45][377] = 9'b111111111;
assign micromatrizz[45][378] = 9'b111111111;
assign micromatrizz[45][379] = 9'b111111111;
assign micromatrizz[45][380] = 9'b111111111;
assign micromatrizz[45][381] = 9'b111111111;
assign micromatrizz[45][382] = 9'b111111111;
assign micromatrizz[45][383] = 9'b111111111;
assign micromatrizz[45][384] = 9'b111111111;
assign micromatrizz[45][385] = 9'b111111111;
assign micromatrizz[45][386] = 9'b111111111;
assign micromatrizz[45][387] = 9'b111111111;
assign micromatrizz[45][388] = 9'b111111111;
assign micromatrizz[45][389] = 9'b111111111;
assign micromatrizz[45][390] = 9'b111111111;
assign micromatrizz[45][391] = 9'b111111111;
assign micromatrizz[45][392] = 9'b111111111;
assign micromatrizz[45][393] = 9'b111111111;
assign micromatrizz[45][394] = 9'b111111111;
assign micromatrizz[45][395] = 9'b111111111;
assign micromatrizz[45][396] = 9'b111111111;
assign micromatrizz[45][397] = 9'b111111111;
assign micromatrizz[45][398] = 9'b111111111;
assign micromatrizz[45][399] = 9'b111111111;
assign micromatrizz[45][400] = 9'b111111111;
assign micromatrizz[45][401] = 9'b111111111;
assign micromatrizz[45][402] = 9'b111111111;
assign micromatrizz[45][403] = 9'b111111111;
assign micromatrizz[45][404] = 9'b111111111;
assign micromatrizz[45][405] = 9'b111111111;
assign micromatrizz[45][406] = 9'b111111111;
assign micromatrizz[45][407] = 9'b111111111;
assign micromatrizz[45][408] = 9'b111111111;
assign micromatrizz[45][409] = 9'b111111111;
assign micromatrizz[45][410] = 9'b111111111;
assign micromatrizz[45][411] = 9'b111111111;
assign micromatrizz[45][412] = 9'b111111111;
assign micromatrizz[45][413] = 9'b111111111;
assign micromatrizz[45][414] = 9'b111111111;
assign micromatrizz[45][415] = 9'b111111111;
assign micromatrizz[45][416] = 9'b111111111;
assign micromatrizz[45][417] = 9'b111111111;
assign micromatrizz[45][418] = 9'b111111111;
assign micromatrizz[45][419] = 9'b111111111;
assign micromatrizz[45][420] = 9'b111111111;
assign micromatrizz[45][421] = 9'b111111111;
assign micromatrizz[45][422] = 9'b111111111;
assign micromatrizz[45][423] = 9'b111111111;
assign micromatrizz[45][424] = 9'b111111111;
assign micromatrizz[45][425] = 9'b111111111;
assign micromatrizz[45][426] = 9'b111111111;
assign micromatrizz[45][427] = 9'b111111111;
assign micromatrizz[45][428] = 9'b111111111;
assign micromatrizz[45][429] = 9'b111111111;
assign micromatrizz[45][430] = 9'b111111111;
assign micromatrizz[45][431] = 9'b111111111;
assign micromatrizz[45][432] = 9'b111111111;
assign micromatrizz[45][433] = 9'b111111111;
assign micromatrizz[45][434] = 9'b111111111;
assign micromatrizz[45][435] = 9'b111111111;
assign micromatrizz[45][436] = 9'b111111111;
assign micromatrizz[45][437] = 9'b111111111;
assign micromatrizz[45][438] = 9'b111111111;
assign micromatrizz[45][439] = 9'b111111111;
assign micromatrizz[45][440] = 9'b111111111;
assign micromatrizz[45][441] = 9'b111111111;
assign micromatrizz[45][442] = 9'b111111111;
assign micromatrizz[45][443] = 9'b111111111;
assign micromatrizz[45][444] = 9'b111111111;
assign micromatrizz[45][445] = 9'b111111111;
assign micromatrizz[45][446] = 9'b111111111;
assign micromatrizz[45][447] = 9'b111111111;
assign micromatrizz[45][448] = 9'b111111111;
assign micromatrizz[45][449] = 9'b111111111;
assign micromatrizz[45][450] = 9'b111111111;
assign micromatrizz[45][451] = 9'b111111111;
assign micromatrizz[45][452] = 9'b111111111;
assign micromatrizz[45][453] = 9'b111111111;
assign micromatrizz[45][454] = 9'b111111111;
assign micromatrizz[45][455] = 9'b111111111;
assign micromatrizz[45][456] = 9'b111111111;
assign micromatrizz[45][457] = 9'b111111111;
assign micromatrizz[45][458] = 9'b111111111;
assign micromatrizz[45][459] = 9'b111111111;
assign micromatrizz[45][460] = 9'b111111111;
assign micromatrizz[45][461] = 9'b111111111;
assign micromatrizz[45][462] = 9'b111111111;
assign micromatrizz[45][463] = 9'b111111111;
assign micromatrizz[45][464] = 9'b111111111;
assign micromatrizz[45][465] = 9'b111111111;
assign micromatrizz[45][466] = 9'b111111111;
assign micromatrizz[45][467] = 9'b111111111;
assign micromatrizz[45][468] = 9'b111111111;
assign micromatrizz[45][469] = 9'b111111111;
assign micromatrizz[45][470] = 9'b111111111;
assign micromatrizz[45][471] = 9'b111111111;
assign micromatrizz[45][472] = 9'b111111111;
assign micromatrizz[45][473] = 9'b111111111;
assign micromatrizz[45][474] = 9'b111111111;
assign micromatrizz[45][475] = 9'b111111111;
assign micromatrizz[45][476] = 9'b111111111;
assign micromatrizz[45][477] = 9'b111111111;
assign micromatrizz[45][478] = 9'b111111111;
assign micromatrizz[45][479] = 9'b111111111;
assign micromatrizz[45][480] = 9'b111111111;
assign micromatrizz[45][481] = 9'b111111111;
assign micromatrizz[45][482] = 9'b111111111;
assign micromatrizz[45][483] = 9'b111111111;
assign micromatrizz[45][484] = 9'b111111111;
assign micromatrizz[45][485] = 9'b111111111;
assign micromatrizz[45][486] = 9'b111111111;
assign micromatrizz[45][487] = 9'b111111111;
assign micromatrizz[45][488] = 9'b111111111;
assign micromatrizz[45][489] = 9'b111111111;
assign micromatrizz[45][490] = 9'b111111111;
assign micromatrizz[45][491] = 9'b111111111;
assign micromatrizz[45][492] = 9'b111111111;
assign micromatrizz[45][493] = 9'b111111111;
assign micromatrizz[45][494] = 9'b111111111;
assign micromatrizz[45][495] = 9'b111111111;
assign micromatrizz[45][496] = 9'b111111111;
assign micromatrizz[45][497] = 9'b111111111;
assign micromatrizz[45][498] = 9'b111111111;
assign micromatrizz[45][499] = 9'b111111111;
assign micromatrizz[45][500] = 9'b111111111;
assign micromatrizz[45][501] = 9'b111111111;
assign micromatrizz[45][502] = 9'b111111111;
assign micromatrizz[45][503] = 9'b111111111;
assign micromatrizz[45][504] = 9'b111111111;
assign micromatrizz[45][505] = 9'b111111111;
assign micromatrizz[45][506] = 9'b111111111;
assign micromatrizz[45][507] = 9'b111111111;
assign micromatrizz[45][508] = 9'b111111111;
assign micromatrizz[45][509] = 9'b111111111;
assign micromatrizz[45][510] = 9'b111111111;
assign micromatrizz[45][511] = 9'b111111111;
assign micromatrizz[45][512] = 9'b111111111;
assign micromatrizz[45][513] = 9'b111111111;
assign micromatrizz[45][514] = 9'b111111111;
assign micromatrizz[45][515] = 9'b111111111;
assign micromatrizz[45][516] = 9'b111111111;
assign micromatrizz[45][517] = 9'b111111111;
assign micromatrizz[45][518] = 9'b111111111;
assign micromatrizz[45][519] = 9'b111111111;
assign micromatrizz[45][520] = 9'b111111111;
assign micromatrizz[45][521] = 9'b111111111;
assign micromatrizz[45][522] = 9'b111111111;
assign micromatrizz[45][523] = 9'b111111111;
assign micromatrizz[45][524] = 9'b111111111;
assign micromatrizz[45][525] = 9'b111111111;
assign micromatrizz[45][526] = 9'b111111111;
assign micromatrizz[45][527] = 9'b111111111;
assign micromatrizz[45][528] = 9'b111111111;
assign micromatrizz[45][529] = 9'b111111111;
assign micromatrizz[45][530] = 9'b111111111;
assign micromatrizz[45][531] = 9'b111111111;
assign micromatrizz[45][532] = 9'b111111111;
assign micromatrizz[45][533] = 9'b111111111;
assign micromatrizz[45][534] = 9'b111111111;
assign micromatrizz[45][535] = 9'b111111111;
assign micromatrizz[45][536] = 9'b111111111;
assign micromatrizz[45][537] = 9'b111111111;
assign micromatrizz[45][538] = 9'b111111111;
assign micromatrizz[45][539] = 9'b111111111;
assign micromatrizz[45][540] = 9'b111111111;
assign micromatrizz[45][541] = 9'b111111111;
assign micromatrizz[45][542] = 9'b111111111;
assign micromatrizz[45][543] = 9'b111111111;
assign micromatrizz[45][544] = 9'b111111111;
assign micromatrizz[45][545] = 9'b111111111;
assign micromatrizz[45][546] = 9'b111111111;
assign micromatrizz[45][547] = 9'b111111111;
assign micromatrizz[45][548] = 9'b111111111;
assign micromatrizz[45][549] = 9'b111111111;
assign micromatrizz[45][550] = 9'b111111111;
assign micromatrizz[45][551] = 9'b111111111;
assign micromatrizz[45][552] = 9'b111111111;
assign micromatrizz[45][553] = 9'b111111111;
assign micromatrizz[45][554] = 9'b111111111;
assign micromatrizz[45][555] = 9'b111111111;
assign micromatrizz[45][556] = 9'b111111111;
assign micromatrizz[45][557] = 9'b111111111;
assign micromatrizz[45][558] = 9'b111111111;
assign micromatrizz[45][559] = 9'b111111111;
assign micromatrizz[45][560] = 9'b111111111;
assign micromatrizz[45][561] = 9'b111111111;
assign micromatrizz[45][562] = 9'b111111111;
assign micromatrizz[45][563] = 9'b111111111;
assign micromatrizz[45][564] = 9'b111111111;
assign micromatrizz[45][565] = 9'b111111111;
assign micromatrizz[45][566] = 9'b111111111;
assign micromatrizz[45][567] = 9'b111111111;
assign micromatrizz[45][568] = 9'b111111111;
assign micromatrizz[45][569] = 9'b111111111;
assign micromatrizz[45][570] = 9'b111111111;
assign micromatrizz[45][571] = 9'b111111111;
assign micromatrizz[45][572] = 9'b111111111;
assign micromatrizz[45][573] = 9'b111111111;
assign micromatrizz[45][574] = 9'b111111111;
assign micromatrizz[45][575] = 9'b111111111;
assign micromatrizz[45][576] = 9'b111111111;
assign micromatrizz[45][577] = 9'b111111111;
assign micromatrizz[45][578] = 9'b111111111;
assign micromatrizz[45][579] = 9'b111111111;
assign micromatrizz[45][580] = 9'b111111111;
assign micromatrizz[45][581] = 9'b111111111;
assign micromatrizz[45][582] = 9'b111111111;
assign micromatrizz[45][583] = 9'b111111111;
assign micromatrizz[45][584] = 9'b111111111;
assign micromatrizz[45][585] = 9'b111111111;
assign micromatrizz[45][586] = 9'b111111111;
assign micromatrizz[45][587] = 9'b111111111;
assign micromatrizz[45][588] = 9'b111111111;
assign micromatrizz[45][589] = 9'b111111111;
assign micromatrizz[45][590] = 9'b111111111;
assign micromatrizz[45][591] = 9'b111111111;
assign micromatrizz[45][592] = 9'b111111111;
assign micromatrizz[45][593] = 9'b111111111;
assign micromatrizz[45][594] = 9'b111111111;
assign micromatrizz[45][595] = 9'b111111111;
assign micromatrizz[45][596] = 9'b111111111;
assign micromatrizz[45][597] = 9'b111111111;
assign micromatrizz[45][598] = 9'b111111111;
assign micromatrizz[45][599] = 9'b111111111;
assign micromatrizz[45][600] = 9'b111111111;
assign micromatrizz[45][601] = 9'b111111111;
assign micromatrizz[45][602] = 9'b111111111;
assign micromatrizz[45][603] = 9'b111111111;
assign micromatrizz[45][604] = 9'b111111111;
assign micromatrizz[45][605] = 9'b111111111;
assign micromatrizz[45][606] = 9'b111111111;
assign micromatrizz[45][607] = 9'b111111111;
assign micromatrizz[45][608] = 9'b111111111;
assign micromatrizz[45][609] = 9'b111111111;
assign micromatrizz[45][610] = 9'b111111111;
assign micromatrizz[45][611] = 9'b111111111;
assign micromatrizz[45][612] = 9'b111111111;
assign micromatrizz[45][613] = 9'b111111111;
assign micromatrizz[45][614] = 9'b111111111;
assign micromatrizz[45][615] = 9'b111111111;
assign micromatrizz[45][616] = 9'b111111111;
assign micromatrizz[45][617] = 9'b111111111;
assign micromatrizz[45][618] = 9'b111111111;
assign micromatrizz[45][619] = 9'b111111111;
assign micromatrizz[45][620] = 9'b111111111;
assign micromatrizz[45][621] = 9'b111111111;
assign micromatrizz[45][622] = 9'b111111111;
assign micromatrizz[45][623] = 9'b111111111;
assign micromatrizz[45][624] = 9'b111111111;
assign micromatrizz[45][625] = 9'b111111111;
assign micromatrizz[45][626] = 9'b111111111;
assign micromatrizz[45][627] = 9'b111111111;
assign micromatrizz[45][628] = 9'b111111111;
assign micromatrizz[45][629] = 9'b111111111;
assign micromatrizz[45][630] = 9'b111111111;
assign micromatrizz[45][631] = 9'b111111111;
assign micromatrizz[45][632] = 9'b111111111;
assign micromatrizz[45][633] = 9'b111111111;
assign micromatrizz[45][634] = 9'b111111111;
assign micromatrizz[45][635] = 9'b111111111;
assign micromatrizz[45][636] = 9'b111111111;
assign micromatrizz[45][637] = 9'b111111111;
assign micromatrizz[45][638] = 9'b111111111;
assign micromatrizz[45][639] = 9'b111111111;
assign micromatrizz[46][0] = 9'b111111111;
assign micromatrizz[46][1] = 9'b111111111;
assign micromatrizz[46][2] = 9'b111111111;
assign micromatrizz[46][3] = 9'b111111111;
assign micromatrizz[46][4] = 9'b111111111;
assign micromatrizz[46][5] = 9'b111111111;
assign micromatrizz[46][6] = 9'b111111111;
assign micromatrizz[46][7] = 9'b111111111;
assign micromatrizz[46][8] = 9'b111111111;
assign micromatrizz[46][9] = 9'b111111111;
assign micromatrizz[46][10] = 9'b111111111;
assign micromatrizz[46][11] = 9'b111111111;
assign micromatrizz[46][12] = 9'b111111111;
assign micromatrizz[46][13] = 9'b111111111;
assign micromatrizz[46][14] = 9'b111111111;
assign micromatrizz[46][15] = 9'b111111111;
assign micromatrizz[46][16] = 9'b111111111;
assign micromatrizz[46][17] = 9'b111111111;
assign micromatrizz[46][18] = 9'b111111111;
assign micromatrizz[46][19] = 9'b111111111;
assign micromatrizz[46][20] = 9'b111111111;
assign micromatrizz[46][21] = 9'b111111111;
assign micromatrizz[46][22] = 9'b111111111;
assign micromatrizz[46][23] = 9'b111111111;
assign micromatrizz[46][24] = 9'b111111111;
assign micromatrizz[46][25] = 9'b111111111;
assign micromatrizz[46][26] = 9'b111111111;
assign micromatrizz[46][27] = 9'b111111111;
assign micromatrizz[46][28] = 9'b111111111;
assign micromatrizz[46][29] = 9'b111111111;
assign micromatrizz[46][30] = 9'b111111111;
assign micromatrizz[46][31] = 9'b111111111;
assign micromatrizz[46][32] = 9'b111111111;
assign micromatrizz[46][33] = 9'b111111111;
assign micromatrizz[46][34] = 9'b111111111;
assign micromatrizz[46][35] = 9'b111111111;
assign micromatrizz[46][36] = 9'b111111111;
assign micromatrizz[46][37] = 9'b111111111;
assign micromatrizz[46][38] = 9'b111111111;
assign micromatrizz[46][39] = 9'b111111111;
assign micromatrizz[46][40] = 9'b111111111;
assign micromatrizz[46][41] = 9'b111111111;
assign micromatrizz[46][42] = 9'b111111111;
assign micromatrizz[46][43] = 9'b111111111;
assign micromatrizz[46][44] = 9'b111111111;
assign micromatrizz[46][45] = 9'b111111111;
assign micromatrizz[46][46] = 9'b111111111;
assign micromatrizz[46][47] = 9'b111111111;
assign micromatrizz[46][48] = 9'b111111111;
assign micromatrizz[46][49] = 9'b111111111;
assign micromatrizz[46][50] = 9'b111111111;
assign micromatrizz[46][51] = 9'b111111111;
assign micromatrizz[46][52] = 9'b111111111;
assign micromatrizz[46][53] = 9'b111111111;
assign micromatrizz[46][54] = 9'b111111111;
assign micromatrizz[46][55] = 9'b111111111;
assign micromatrizz[46][56] = 9'b111111111;
assign micromatrizz[46][57] = 9'b111111111;
assign micromatrizz[46][58] = 9'b111111111;
assign micromatrizz[46][59] = 9'b111111111;
assign micromatrizz[46][60] = 9'b111111111;
assign micromatrizz[46][61] = 9'b111111111;
assign micromatrizz[46][62] = 9'b111111111;
assign micromatrizz[46][63] = 9'b111111111;
assign micromatrizz[46][64] = 9'b111111111;
assign micromatrizz[46][65] = 9'b111111111;
assign micromatrizz[46][66] = 9'b111111111;
assign micromatrizz[46][67] = 9'b111111111;
assign micromatrizz[46][68] = 9'b111111111;
assign micromatrizz[46][69] = 9'b111111111;
assign micromatrizz[46][70] = 9'b111111111;
assign micromatrizz[46][71] = 9'b111111111;
assign micromatrizz[46][72] = 9'b111111111;
assign micromatrizz[46][73] = 9'b111111111;
assign micromatrizz[46][74] = 9'b111111111;
assign micromatrizz[46][75] = 9'b111111111;
assign micromatrizz[46][76] = 9'b111111111;
assign micromatrizz[46][77] = 9'b111111111;
assign micromatrizz[46][78] = 9'b111111111;
assign micromatrizz[46][79] = 9'b111111111;
assign micromatrizz[46][80] = 9'b111111111;
assign micromatrizz[46][81] = 9'b111111111;
assign micromatrizz[46][82] = 9'b111111111;
assign micromatrizz[46][83] = 9'b111111111;
assign micromatrizz[46][84] = 9'b111111111;
assign micromatrizz[46][85] = 9'b111111111;
assign micromatrizz[46][86] = 9'b111111111;
assign micromatrizz[46][87] = 9'b111111111;
assign micromatrizz[46][88] = 9'b111111111;
assign micromatrizz[46][89] = 9'b111111111;
assign micromatrizz[46][90] = 9'b111111111;
assign micromatrizz[46][91] = 9'b111111111;
assign micromatrizz[46][92] = 9'b111111111;
assign micromatrizz[46][93] = 9'b111111111;
assign micromatrizz[46][94] = 9'b111111111;
assign micromatrizz[46][95] = 9'b111111111;
assign micromatrizz[46][96] = 9'b111111111;
assign micromatrizz[46][97] = 9'b111111111;
assign micromatrizz[46][98] = 9'b111111111;
assign micromatrizz[46][99] = 9'b111111111;
assign micromatrizz[46][100] = 9'b111111111;
assign micromatrizz[46][101] = 9'b111111111;
assign micromatrizz[46][102] = 9'b111111111;
assign micromatrizz[46][103] = 9'b111111111;
assign micromatrizz[46][104] = 9'b111111111;
assign micromatrizz[46][105] = 9'b111111111;
assign micromatrizz[46][106] = 9'b111111111;
assign micromatrizz[46][107] = 9'b111111111;
assign micromatrizz[46][108] = 9'b111111111;
assign micromatrizz[46][109] = 9'b111111111;
assign micromatrizz[46][110] = 9'b111111111;
assign micromatrizz[46][111] = 9'b111111111;
assign micromatrizz[46][112] = 9'b111111111;
assign micromatrizz[46][113] = 9'b111111111;
assign micromatrizz[46][114] = 9'b111111111;
assign micromatrizz[46][115] = 9'b111111111;
assign micromatrizz[46][116] = 9'b111111111;
assign micromatrizz[46][117] = 9'b111111111;
assign micromatrizz[46][118] = 9'b111111111;
assign micromatrizz[46][119] = 9'b111111111;
assign micromatrizz[46][120] = 9'b111111111;
assign micromatrizz[46][121] = 9'b111111111;
assign micromatrizz[46][122] = 9'b111111111;
assign micromatrizz[46][123] = 9'b111111111;
assign micromatrizz[46][124] = 9'b111111111;
assign micromatrizz[46][125] = 9'b111111111;
assign micromatrizz[46][126] = 9'b111111111;
assign micromatrizz[46][127] = 9'b111111111;
assign micromatrizz[46][128] = 9'b111111111;
assign micromatrizz[46][129] = 9'b111111111;
assign micromatrizz[46][130] = 9'b111111111;
assign micromatrizz[46][131] = 9'b111111111;
assign micromatrizz[46][132] = 9'b111111111;
assign micromatrizz[46][133] = 9'b111111111;
assign micromatrizz[46][134] = 9'b111111111;
assign micromatrizz[46][135] = 9'b111111111;
assign micromatrizz[46][136] = 9'b111111111;
assign micromatrizz[46][137] = 9'b111111111;
assign micromatrizz[46][138] = 9'b111111111;
assign micromatrizz[46][139] = 9'b111111111;
assign micromatrizz[46][140] = 9'b111111111;
assign micromatrizz[46][141] = 9'b111111111;
assign micromatrizz[46][142] = 9'b111111111;
assign micromatrizz[46][143] = 9'b111111111;
assign micromatrizz[46][144] = 9'b111111111;
assign micromatrizz[46][145] = 9'b111110111;
assign micromatrizz[46][146] = 9'b111110010;
assign micromatrizz[46][147] = 9'b111110011;
assign micromatrizz[46][148] = 9'b111110011;
assign micromatrizz[46][149] = 9'b111110010;
assign micromatrizz[46][150] = 9'b111110011;
assign micromatrizz[46][151] = 9'b111110011;
assign micromatrizz[46][152] = 9'b111110111;
assign micromatrizz[46][153] = 9'b111110111;
assign micromatrizz[46][154] = 9'b111111111;
assign micromatrizz[46][155] = 9'b111111111;
assign micromatrizz[46][156] = 9'b111111111;
assign micromatrizz[46][157] = 9'b111111111;
assign micromatrizz[46][158] = 9'b111111111;
assign micromatrizz[46][159] = 9'b111111111;
assign micromatrizz[46][160] = 9'b111111111;
assign micromatrizz[46][161] = 9'b111111111;
assign micromatrizz[46][162] = 9'b111111111;
assign micromatrizz[46][163] = 9'b111111111;
assign micromatrizz[46][164] = 9'b111111111;
assign micromatrizz[46][165] = 9'b111111111;
assign micromatrizz[46][166] = 9'b111111111;
assign micromatrizz[46][167] = 9'b111111111;
assign micromatrizz[46][168] = 9'b111111111;
assign micromatrizz[46][169] = 9'b111111111;
assign micromatrizz[46][170] = 9'b111111111;
assign micromatrizz[46][171] = 9'b111111111;
assign micromatrizz[46][172] = 9'b111111111;
assign micromatrizz[46][173] = 9'b111111111;
assign micromatrizz[46][174] = 9'b111111111;
assign micromatrizz[46][175] = 9'b111111111;
assign micromatrizz[46][176] = 9'b111111111;
assign micromatrizz[46][177] = 9'b111111111;
assign micromatrizz[46][178] = 9'b111111111;
assign micromatrizz[46][179] = 9'b111111111;
assign micromatrizz[46][180] = 9'b111111111;
assign micromatrizz[46][181] = 9'b111111111;
assign micromatrizz[46][182] = 9'b111111111;
assign micromatrizz[46][183] = 9'b111111111;
assign micromatrizz[46][184] = 9'b111111111;
assign micromatrizz[46][185] = 9'b111111111;
assign micromatrizz[46][186] = 9'b111111111;
assign micromatrizz[46][187] = 9'b111111111;
assign micromatrizz[46][188] = 9'b111111111;
assign micromatrizz[46][189] = 9'b111111111;
assign micromatrizz[46][190] = 9'b111111111;
assign micromatrizz[46][191] = 9'b111111111;
assign micromatrizz[46][192] = 9'b111111111;
assign micromatrizz[46][193] = 9'b111111111;
assign micromatrizz[46][194] = 9'b111111111;
assign micromatrizz[46][195] = 9'b111111111;
assign micromatrizz[46][196] = 9'b111111111;
assign micromatrizz[46][197] = 9'b111111111;
assign micromatrizz[46][198] = 9'b111111111;
assign micromatrizz[46][199] = 9'b111111111;
assign micromatrizz[46][200] = 9'b111111111;
assign micromatrizz[46][201] = 9'b111111111;
assign micromatrizz[46][202] = 9'b111111111;
assign micromatrizz[46][203] = 9'b111111111;
assign micromatrizz[46][204] = 9'b111111111;
assign micromatrizz[46][205] = 9'b111111111;
assign micromatrizz[46][206] = 9'b111111111;
assign micromatrizz[46][207] = 9'b111111111;
assign micromatrizz[46][208] = 9'b111111111;
assign micromatrizz[46][209] = 9'b111111111;
assign micromatrizz[46][210] = 9'b111111111;
assign micromatrizz[46][211] = 9'b111111111;
assign micromatrizz[46][212] = 9'b111111111;
assign micromatrizz[46][213] = 9'b111111111;
assign micromatrizz[46][214] = 9'b111111111;
assign micromatrizz[46][215] = 9'b111111111;
assign micromatrizz[46][216] = 9'b111111111;
assign micromatrizz[46][217] = 9'b111111111;
assign micromatrizz[46][218] = 9'b111111111;
assign micromatrizz[46][219] = 9'b111111111;
assign micromatrizz[46][220] = 9'b111111111;
assign micromatrizz[46][221] = 9'b111111111;
assign micromatrizz[46][222] = 9'b111111111;
assign micromatrizz[46][223] = 9'b111111111;
assign micromatrizz[46][224] = 9'b111111111;
assign micromatrizz[46][225] = 9'b111111111;
assign micromatrizz[46][226] = 9'b111111111;
assign micromatrizz[46][227] = 9'b111111111;
assign micromatrizz[46][228] = 9'b111111111;
assign micromatrizz[46][229] = 9'b111111111;
assign micromatrizz[46][230] = 9'b111111111;
assign micromatrizz[46][231] = 9'b111111111;
assign micromatrizz[46][232] = 9'b111111111;
assign micromatrizz[46][233] = 9'b111111111;
assign micromatrizz[46][234] = 9'b111111111;
assign micromatrizz[46][235] = 9'b111111111;
assign micromatrizz[46][236] = 9'b111111111;
assign micromatrizz[46][237] = 9'b111111111;
assign micromatrizz[46][238] = 9'b111111111;
assign micromatrizz[46][239] = 9'b111111111;
assign micromatrizz[46][240] = 9'b111111111;
assign micromatrizz[46][241] = 9'b111111111;
assign micromatrizz[46][242] = 9'b111111111;
assign micromatrizz[46][243] = 9'b111111111;
assign micromatrizz[46][244] = 9'b111111111;
assign micromatrizz[46][245] = 9'b111111111;
assign micromatrizz[46][246] = 9'b111111111;
assign micromatrizz[46][247] = 9'b111111111;
assign micromatrizz[46][248] = 9'b111111111;
assign micromatrizz[46][249] = 9'b111111111;
assign micromatrizz[46][250] = 9'b111111111;
assign micromatrizz[46][251] = 9'b111111111;
assign micromatrizz[46][252] = 9'b111111111;
assign micromatrizz[46][253] = 9'b111111111;
assign micromatrizz[46][254] = 9'b111111111;
assign micromatrizz[46][255] = 9'b111111111;
assign micromatrizz[46][256] = 9'b111111111;
assign micromatrizz[46][257] = 9'b111111111;
assign micromatrizz[46][258] = 9'b111111111;
assign micromatrizz[46][259] = 9'b111111111;
assign micromatrizz[46][260] = 9'b111111111;
assign micromatrizz[46][261] = 9'b111111111;
assign micromatrizz[46][262] = 9'b111111111;
assign micromatrizz[46][263] = 9'b111111111;
assign micromatrizz[46][264] = 9'b111111111;
assign micromatrizz[46][265] = 9'b111111111;
assign micromatrizz[46][266] = 9'b111111111;
assign micromatrizz[46][267] = 9'b111111111;
assign micromatrizz[46][268] = 9'b111111111;
assign micromatrizz[46][269] = 9'b111111111;
assign micromatrizz[46][270] = 9'b111111111;
assign micromatrizz[46][271] = 9'b111111111;
assign micromatrizz[46][272] = 9'b111111111;
assign micromatrizz[46][273] = 9'b111111111;
assign micromatrizz[46][274] = 9'b111111111;
assign micromatrizz[46][275] = 9'b111111111;
assign micromatrizz[46][276] = 9'b111111111;
assign micromatrizz[46][277] = 9'b111111111;
assign micromatrizz[46][278] = 9'b111111111;
assign micromatrizz[46][279] = 9'b111111111;
assign micromatrizz[46][280] = 9'b111111111;
assign micromatrizz[46][281] = 9'b111111111;
assign micromatrizz[46][282] = 9'b111111111;
assign micromatrizz[46][283] = 9'b111111111;
assign micromatrizz[46][284] = 9'b111111111;
assign micromatrizz[46][285] = 9'b111111111;
assign micromatrizz[46][286] = 9'b111111111;
assign micromatrizz[46][287] = 9'b111111111;
assign micromatrizz[46][288] = 9'b111111111;
assign micromatrizz[46][289] = 9'b111111111;
assign micromatrizz[46][290] = 9'b111111111;
assign micromatrizz[46][291] = 9'b111111111;
assign micromatrizz[46][292] = 9'b111111111;
assign micromatrizz[46][293] = 9'b111111111;
assign micromatrizz[46][294] = 9'b111111111;
assign micromatrizz[46][295] = 9'b111111111;
assign micromatrizz[46][296] = 9'b111111111;
assign micromatrizz[46][297] = 9'b111111111;
assign micromatrizz[46][298] = 9'b111111111;
assign micromatrizz[46][299] = 9'b111111111;
assign micromatrizz[46][300] = 9'b111111111;
assign micromatrizz[46][301] = 9'b111111111;
assign micromatrizz[46][302] = 9'b111111111;
assign micromatrizz[46][303] = 9'b111111111;
assign micromatrizz[46][304] = 9'b111111111;
assign micromatrizz[46][305] = 9'b111111111;
assign micromatrizz[46][306] = 9'b111111111;
assign micromatrizz[46][307] = 9'b111111111;
assign micromatrizz[46][308] = 9'b111111111;
assign micromatrizz[46][309] = 9'b111111111;
assign micromatrizz[46][310] = 9'b111111111;
assign micromatrizz[46][311] = 9'b111111111;
assign micromatrizz[46][312] = 9'b111111111;
assign micromatrizz[46][313] = 9'b111111111;
assign micromatrizz[46][314] = 9'b111111111;
assign micromatrizz[46][315] = 9'b111111111;
assign micromatrizz[46][316] = 9'b111111111;
assign micromatrizz[46][317] = 9'b111111111;
assign micromatrizz[46][318] = 9'b111111111;
assign micromatrizz[46][319] = 9'b111111111;
assign micromatrizz[46][320] = 9'b111111111;
assign micromatrizz[46][321] = 9'b111111111;
assign micromatrizz[46][322] = 9'b111111111;
assign micromatrizz[46][323] = 9'b111111111;
assign micromatrizz[46][324] = 9'b111111111;
assign micromatrizz[46][325] = 9'b111111111;
assign micromatrizz[46][326] = 9'b111111111;
assign micromatrizz[46][327] = 9'b111111111;
assign micromatrizz[46][328] = 9'b111111111;
assign micromatrizz[46][329] = 9'b111111111;
assign micromatrizz[46][330] = 9'b111111111;
assign micromatrizz[46][331] = 9'b111111111;
assign micromatrizz[46][332] = 9'b111111111;
assign micromatrizz[46][333] = 9'b111111111;
assign micromatrizz[46][334] = 9'b111111111;
assign micromatrizz[46][335] = 9'b111111111;
assign micromatrizz[46][336] = 9'b111111111;
assign micromatrizz[46][337] = 9'b111111111;
assign micromatrizz[46][338] = 9'b111111111;
assign micromatrizz[46][339] = 9'b111111111;
assign micromatrizz[46][340] = 9'b111111111;
assign micromatrizz[46][341] = 9'b111111111;
assign micromatrizz[46][342] = 9'b111111111;
assign micromatrizz[46][343] = 9'b111111111;
assign micromatrizz[46][344] = 9'b111111111;
assign micromatrizz[46][345] = 9'b111111111;
assign micromatrizz[46][346] = 9'b111111111;
assign micromatrizz[46][347] = 9'b111111111;
assign micromatrizz[46][348] = 9'b111111111;
assign micromatrizz[46][349] = 9'b111111111;
assign micromatrizz[46][350] = 9'b111111111;
assign micromatrizz[46][351] = 9'b111111111;
assign micromatrizz[46][352] = 9'b111111111;
assign micromatrizz[46][353] = 9'b111111111;
assign micromatrizz[46][354] = 9'b111111111;
assign micromatrizz[46][355] = 9'b111111111;
assign micromatrizz[46][356] = 9'b111111111;
assign micromatrizz[46][357] = 9'b111111111;
assign micromatrizz[46][358] = 9'b111111111;
assign micromatrizz[46][359] = 9'b111111111;
assign micromatrizz[46][360] = 9'b111111111;
assign micromatrizz[46][361] = 9'b111111111;
assign micromatrizz[46][362] = 9'b111111111;
assign micromatrizz[46][363] = 9'b111111111;
assign micromatrizz[46][364] = 9'b111111111;
assign micromatrizz[46][365] = 9'b111111111;
assign micromatrizz[46][366] = 9'b111111111;
assign micromatrizz[46][367] = 9'b111111111;
assign micromatrizz[46][368] = 9'b111111111;
assign micromatrizz[46][369] = 9'b111111111;
assign micromatrizz[46][370] = 9'b111111111;
assign micromatrizz[46][371] = 9'b111111111;
assign micromatrizz[46][372] = 9'b111111111;
assign micromatrizz[46][373] = 9'b111111111;
assign micromatrizz[46][374] = 9'b111111111;
assign micromatrizz[46][375] = 9'b111111111;
assign micromatrizz[46][376] = 9'b111111111;
assign micromatrizz[46][377] = 9'b111111111;
assign micromatrizz[46][378] = 9'b111111111;
assign micromatrizz[46][379] = 9'b111111111;
assign micromatrizz[46][380] = 9'b111111111;
assign micromatrizz[46][381] = 9'b111111111;
assign micromatrizz[46][382] = 9'b111111111;
assign micromatrizz[46][383] = 9'b111111111;
assign micromatrizz[46][384] = 9'b111111111;
assign micromatrizz[46][385] = 9'b111111111;
assign micromatrizz[46][386] = 9'b111111111;
assign micromatrizz[46][387] = 9'b111111111;
assign micromatrizz[46][388] = 9'b111111111;
assign micromatrizz[46][389] = 9'b111111111;
assign micromatrizz[46][390] = 9'b111111111;
assign micromatrizz[46][391] = 9'b111111111;
assign micromatrizz[46][392] = 9'b111111111;
assign micromatrizz[46][393] = 9'b111111111;
assign micromatrizz[46][394] = 9'b111111111;
assign micromatrizz[46][395] = 9'b111111111;
assign micromatrizz[46][396] = 9'b111111111;
assign micromatrizz[46][397] = 9'b111111111;
assign micromatrizz[46][398] = 9'b111111111;
assign micromatrizz[46][399] = 9'b111111111;
assign micromatrizz[46][400] = 9'b111111111;
assign micromatrizz[46][401] = 9'b111111111;
assign micromatrizz[46][402] = 9'b111111111;
assign micromatrizz[46][403] = 9'b111111111;
assign micromatrizz[46][404] = 9'b111111111;
assign micromatrizz[46][405] = 9'b111111111;
assign micromatrizz[46][406] = 9'b111111111;
assign micromatrizz[46][407] = 9'b111111111;
assign micromatrizz[46][408] = 9'b111111111;
assign micromatrizz[46][409] = 9'b111111111;
assign micromatrizz[46][410] = 9'b111111111;
assign micromatrizz[46][411] = 9'b111111111;
assign micromatrizz[46][412] = 9'b111111111;
assign micromatrizz[46][413] = 9'b111111111;
assign micromatrizz[46][414] = 9'b111111111;
assign micromatrizz[46][415] = 9'b111111111;
assign micromatrizz[46][416] = 9'b111111111;
assign micromatrizz[46][417] = 9'b111111111;
assign micromatrizz[46][418] = 9'b111111111;
assign micromatrizz[46][419] = 9'b111111111;
assign micromatrizz[46][420] = 9'b111111111;
assign micromatrizz[46][421] = 9'b111111111;
assign micromatrizz[46][422] = 9'b111111111;
assign micromatrizz[46][423] = 9'b111111111;
assign micromatrizz[46][424] = 9'b111111111;
assign micromatrizz[46][425] = 9'b111111111;
assign micromatrizz[46][426] = 9'b111111111;
assign micromatrizz[46][427] = 9'b111111111;
assign micromatrizz[46][428] = 9'b111111111;
assign micromatrizz[46][429] = 9'b111111111;
assign micromatrizz[46][430] = 9'b111111111;
assign micromatrizz[46][431] = 9'b111111111;
assign micromatrizz[46][432] = 9'b111111111;
assign micromatrizz[46][433] = 9'b111111111;
assign micromatrizz[46][434] = 9'b111111111;
assign micromatrizz[46][435] = 9'b111111111;
assign micromatrizz[46][436] = 9'b111111111;
assign micromatrizz[46][437] = 9'b111111111;
assign micromatrizz[46][438] = 9'b111111111;
assign micromatrizz[46][439] = 9'b111111111;
assign micromatrizz[46][440] = 9'b111111111;
assign micromatrizz[46][441] = 9'b111111111;
assign micromatrizz[46][442] = 9'b111111111;
assign micromatrizz[46][443] = 9'b111111111;
assign micromatrizz[46][444] = 9'b111111111;
assign micromatrizz[46][445] = 9'b111111111;
assign micromatrizz[46][446] = 9'b111111111;
assign micromatrizz[46][447] = 9'b111111111;
assign micromatrizz[46][448] = 9'b111111111;
assign micromatrizz[46][449] = 9'b111111111;
assign micromatrizz[46][450] = 9'b111111111;
assign micromatrizz[46][451] = 9'b111111111;
assign micromatrizz[46][452] = 9'b111111111;
assign micromatrizz[46][453] = 9'b111111111;
assign micromatrizz[46][454] = 9'b111111111;
assign micromatrizz[46][455] = 9'b111111111;
assign micromatrizz[46][456] = 9'b111111111;
assign micromatrizz[46][457] = 9'b111111111;
assign micromatrizz[46][458] = 9'b111111111;
assign micromatrizz[46][459] = 9'b111111111;
assign micromatrizz[46][460] = 9'b111111111;
assign micromatrizz[46][461] = 9'b111111111;
assign micromatrizz[46][462] = 9'b111111111;
assign micromatrizz[46][463] = 9'b111111111;
assign micromatrizz[46][464] = 9'b111111111;
assign micromatrizz[46][465] = 9'b111111111;
assign micromatrizz[46][466] = 9'b111111111;
assign micromatrizz[46][467] = 9'b111111111;
assign micromatrizz[46][468] = 9'b111111111;
assign micromatrizz[46][469] = 9'b111111111;
assign micromatrizz[46][470] = 9'b111111111;
assign micromatrizz[46][471] = 9'b111111111;
assign micromatrizz[46][472] = 9'b111111111;
assign micromatrizz[46][473] = 9'b111111111;
assign micromatrizz[46][474] = 9'b111111111;
assign micromatrizz[46][475] = 9'b111111111;
assign micromatrizz[46][476] = 9'b111111111;
assign micromatrizz[46][477] = 9'b111111111;
assign micromatrizz[46][478] = 9'b111111111;
assign micromatrizz[46][479] = 9'b111111111;
assign micromatrizz[46][480] = 9'b111111111;
assign micromatrizz[46][481] = 9'b111111111;
assign micromatrizz[46][482] = 9'b111111111;
assign micromatrizz[46][483] = 9'b111111111;
assign micromatrizz[46][484] = 9'b111111111;
assign micromatrizz[46][485] = 9'b111111111;
assign micromatrizz[46][486] = 9'b111111111;
assign micromatrizz[46][487] = 9'b111111111;
assign micromatrizz[46][488] = 9'b111111111;
assign micromatrizz[46][489] = 9'b111111111;
assign micromatrizz[46][490] = 9'b111111111;
assign micromatrizz[46][491] = 9'b111111111;
assign micromatrizz[46][492] = 9'b111111111;
assign micromatrizz[46][493] = 9'b111111111;
assign micromatrizz[46][494] = 9'b111111111;
assign micromatrizz[46][495] = 9'b111111111;
assign micromatrizz[46][496] = 9'b111111111;
assign micromatrizz[46][497] = 9'b111111111;
assign micromatrizz[46][498] = 9'b111111111;
assign micromatrizz[46][499] = 9'b111111111;
assign micromatrizz[46][500] = 9'b111111111;
assign micromatrizz[46][501] = 9'b111111111;
assign micromatrizz[46][502] = 9'b111111111;
assign micromatrizz[46][503] = 9'b111111111;
assign micromatrizz[46][504] = 9'b111111111;
assign micromatrizz[46][505] = 9'b111111111;
assign micromatrizz[46][506] = 9'b111111111;
assign micromatrizz[46][507] = 9'b111111111;
assign micromatrizz[46][508] = 9'b111111111;
assign micromatrizz[46][509] = 9'b111111111;
assign micromatrizz[46][510] = 9'b111111111;
assign micromatrizz[46][511] = 9'b111111111;
assign micromatrizz[46][512] = 9'b111111111;
assign micromatrizz[46][513] = 9'b111111111;
assign micromatrizz[46][514] = 9'b111111111;
assign micromatrizz[46][515] = 9'b111111111;
assign micromatrizz[46][516] = 9'b111111111;
assign micromatrizz[46][517] = 9'b111111111;
assign micromatrizz[46][518] = 9'b111111111;
assign micromatrizz[46][519] = 9'b111111111;
assign micromatrizz[46][520] = 9'b111111111;
assign micromatrizz[46][521] = 9'b111111111;
assign micromatrizz[46][522] = 9'b111111111;
assign micromatrizz[46][523] = 9'b111111111;
assign micromatrizz[46][524] = 9'b111111111;
assign micromatrizz[46][525] = 9'b111111111;
assign micromatrizz[46][526] = 9'b111111111;
assign micromatrizz[46][527] = 9'b111111111;
assign micromatrizz[46][528] = 9'b111111111;
assign micromatrizz[46][529] = 9'b111111111;
assign micromatrizz[46][530] = 9'b111111111;
assign micromatrizz[46][531] = 9'b111111111;
assign micromatrizz[46][532] = 9'b111111111;
assign micromatrizz[46][533] = 9'b111111111;
assign micromatrizz[46][534] = 9'b111111111;
assign micromatrizz[46][535] = 9'b111111111;
assign micromatrizz[46][536] = 9'b111111111;
assign micromatrizz[46][537] = 9'b111111111;
assign micromatrizz[46][538] = 9'b111111111;
assign micromatrizz[46][539] = 9'b111111111;
assign micromatrizz[46][540] = 9'b111111111;
assign micromatrizz[46][541] = 9'b111111111;
assign micromatrizz[46][542] = 9'b111111111;
assign micromatrizz[46][543] = 9'b111111111;
assign micromatrizz[46][544] = 9'b111111111;
assign micromatrizz[46][545] = 9'b111111111;
assign micromatrizz[46][546] = 9'b111111111;
assign micromatrizz[46][547] = 9'b111111111;
assign micromatrizz[46][548] = 9'b111111111;
assign micromatrizz[46][549] = 9'b111111111;
assign micromatrizz[46][550] = 9'b111111111;
assign micromatrizz[46][551] = 9'b111111111;
assign micromatrizz[46][552] = 9'b111111111;
assign micromatrizz[46][553] = 9'b111111111;
assign micromatrizz[46][554] = 9'b111111111;
assign micromatrizz[46][555] = 9'b111111111;
assign micromatrizz[46][556] = 9'b111111111;
assign micromatrizz[46][557] = 9'b111111111;
assign micromatrizz[46][558] = 9'b111111111;
assign micromatrizz[46][559] = 9'b111111111;
assign micromatrizz[46][560] = 9'b111111111;
assign micromatrizz[46][561] = 9'b111111111;
assign micromatrizz[46][562] = 9'b111111111;
assign micromatrizz[46][563] = 9'b111111111;
assign micromatrizz[46][564] = 9'b111111111;
assign micromatrizz[46][565] = 9'b111111111;
assign micromatrizz[46][566] = 9'b111111111;
assign micromatrizz[46][567] = 9'b111111111;
assign micromatrizz[46][568] = 9'b111111111;
assign micromatrizz[46][569] = 9'b111111111;
assign micromatrizz[46][570] = 9'b111111111;
assign micromatrizz[46][571] = 9'b111111111;
assign micromatrizz[46][572] = 9'b111111111;
assign micromatrizz[46][573] = 9'b111111111;
assign micromatrizz[46][574] = 9'b111111111;
assign micromatrizz[46][575] = 9'b111111111;
assign micromatrizz[46][576] = 9'b111111111;
assign micromatrizz[46][577] = 9'b111111111;
assign micromatrizz[46][578] = 9'b111111111;
assign micromatrizz[46][579] = 9'b111111111;
assign micromatrizz[46][580] = 9'b111111111;
assign micromatrizz[46][581] = 9'b111111111;
assign micromatrizz[46][582] = 9'b111111111;
assign micromatrizz[46][583] = 9'b111111111;
assign micromatrizz[46][584] = 9'b111111111;
assign micromatrizz[46][585] = 9'b111111111;
assign micromatrizz[46][586] = 9'b111111111;
assign micromatrizz[46][587] = 9'b111111111;
assign micromatrizz[46][588] = 9'b111111111;
assign micromatrizz[46][589] = 9'b111111111;
assign micromatrizz[46][590] = 9'b111111111;
assign micromatrizz[46][591] = 9'b111111111;
assign micromatrizz[46][592] = 9'b111111111;
assign micromatrizz[46][593] = 9'b111111111;
assign micromatrizz[46][594] = 9'b111111111;
assign micromatrizz[46][595] = 9'b111111111;
assign micromatrizz[46][596] = 9'b111111111;
assign micromatrizz[46][597] = 9'b111111111;
assign micromatrizz[46][598] = 9'b111111111;
assign micromatrizz[46][599] = 9'b111111111;
assign micromatrizz[46][600] = 9'b111111111;
assign micromatrizz[46][601] = 9'b111111111;
assign micromatrizz[46][602] = 9'b111111111;
assign micromatrizz[46][603] = 9'b111111111;
assign micromatrizz[46][604] = 9'b111111111;
assign micromatrizz[46][605] = 9'b111111111;
assign micromatrizz[46][606] = 9'b111111111;
assign micromatrizz[46][607] = 9'b111111111;
assign micromatrizz[46][608] = 9'b111111111;
assign micromatrizz[46][609] = 9'b111111111;
assign micromatrizz[46][610] = 9'b111111111;
assign micromatrizz[46][611] = 9'b111111111;
assign micromatrizz[46][612] = 9'b111111111;
assign micromatrizz[46][613] = 9'b111111111;
assign micromatrizz[46][614] = 9'b111111111;
assign micromatrizz[46][615] = 9'b111111111;
assign micromatrizz[46][616] = 9'b111111111;
assign micromatrizz[46][617] = 9'b111111111;
assign micromatrizz[46][618] = 9'b111111111;
assign micromatrizz[46][619] = 9'b111111111;
assign micromatrizz[46][620] = 9'b111111111;
assign micromatrizz[46][621] = 9'b111111111;
assign micromatrizz[46][622] = 9'b111111111;
assign micromatrizz[46][623] = 9'b111111111;
assign micromatrizz[46][624] = 9'b111111111;
assign micromatrizz[46][625] = 9'b111111111;
assign micromatrizz[46][626] = 9'b111111111;
assign micromatrizz[46][627] = 9'b111111111;
assign micromatrizz[46][628] = 9'b111111111;
assign micromatrizz[46][629] = 9'b111111111;
assign micromatrizz[46][630] = 9'b111111111;
assign micromatrizz[46][631] = 9'b111111111;
assign micromatrizz[46][632] = 9'b111111111;
assign micromatrizz[46][633] = 9'b111111111;
assign micromatrizz[46][634] = 9'b111111111;
assign micromatrizz[46][635] = 9'b111111111;
assign micromatrizz[46][636] = 9'b111111111;
assign micromatrizz[46][637] = 9'b111111111;
assign micromatrizz[46][638] = 9'b111111111;
assign micromatrizz[46][639] = 9'b111111111;
assign micromatrizz[47][0] = 9'b111111111;
assign micromatrizz[47][1] = 9'b111111111;
assign micromatrizz[47][2] = 9'b111111111;
assign micromatrizz[47][3] = 9'b111111111;
assign micromatrizz[47][4] = 9'b111111111;
assign micromatrizz[47][5] = 9'b111111111;
assign micromatrizz[47][6] = 9'b111111111;
assign micromatrizz[47][7] = 9'b111111111;
assign micromatrizz[47][8] = 9'b111111111;
assign micromatrizz[47][9] = 9'b111111111;
assign micromatrizz[47][10] = 9'b111111111;
assign micromatrizz[47][11] = 9'b111111111;
assign micromatrizz[47][12] = 9'b111111111;
assign micromatrizz[47][13] = 9'b111111111;
assign micromatrizz[47][14] = 9'b111111111;
assign micromatrizz[47][15] = 9'b111111111;
assign micromatrizz[47][16] = 9'b111111111;
assign micromatrizz[47][17] = 9'b111111111;
assign micromatrizz[47][18] = 9'b111111111;
assign micromatrizz[47][19] = 9'b111111111;
assign micromatrizz[47][20] = 9'b111111111;
assign micromatrizz[47][21] = 9'b111111111;
assign micromatrizz[47][22] = 9'b111111111;
assign micromatrizz[47][23] = 9'b111111111;
assign micromatrizz[47][24] = 9'b111111111;
assign micromatrizz[47][25] = 9'b111111111;
assign micromatrizz[47][26] = 9'b111111111;
assign micromatrizz[47][27] = 9'b111111111;
assign micromatrizz[47][28] = 9'b111111111;
assign micromatrizz[47][29] = 9'b111111111;
assign micromatrizz[47][30] = 9'b111111111;
assign micromatrizz[47][31] = 9'b111111111;
assign micromatrizz[47][32] = 9'b111111111;
assign micromatrizz[47][33] = 9'b111111111;
assign micromatrizz[47][34] = 9'b111111111;
assign micromatrizz[47][35] = 9'b111111111;
assign micromatrizz[47][36] = 9'b111111111;
assign micromatrizz[47][37] = 9'b111111111;
assign micromatrizz[47][38] = 9'b111111111;
assign micromatrizz[47][39] = 9'b111111111;
assign micromatrizz[47][40] = 9'b111111111;
assign micromatrizz[47][41] = 9'b111111111;
assign micromatrizz[47][42] = 9'b111111111;
assign micromatrizz[47][43] = 9'b111111111;
assign micromatrizz[47][44] = 9'b111111111;
assign micromatrizz[47][45] = 9'b111111111;
assign micromatrizz[47][46] = 9'b111111111;
assign micromatrizz[47][47] = 9'b111111111;
assign micromatrizz[47][48] = 9'b111111111;
assign micromatrizz[47][49] = 9'b111111111;
assign micromatrizz[47][50] = 9'b111111111;
assign micromatrizz[47][51] = 9'b111111111;
assign micromatrizz[47][52] = 9'b111111111;
assign micromatrizz[47][53] = 9'b111111111;
assign micromatrizz[47][54] = 9'b111111111;
assign micromatrizz[47][55] = 9'b111111111;
assign micromatrizz[47][56] = 9'b111111111;
assign micromatrizz[47][57] = 9'b111111111;
assign micromatrizz[47][58] = 9'b111111111;
assign micromatrizz[47][59] = 9'b111111111;
assign micromatrizz[47][60] = 9'b111111111;
assign micromatrizz[47][61] = 9'b111111111;
assign micromatrizz[47][62] = 9'b111111111;
assign micromatrizz[47][63] = 9'b111111111;
assign micromatrizz[47][64] = 9'b111111111;
assign micromatrizz[47][65] = 9'b111111111;
assign micromatrizz[47][66] = 9'b111111111;
assign micromatrizz[47][67] = 9'b111111111;
assign micromatrizz[47][68] = 9'b111111111;
assign micromatrizz[47][69] = 9'b111111111;
assign micromatrizz[47][70] = 9'b111111111;
assign micromatrizz[47][71] = 9'b111111111;
assign micromatrizz[47][72] = 9'b111111111;
assign micromatrizz[47][73] = 9'b111111111;
assign micromatrizz[47][74] = 9'b111111111;
assign micromatrizz[47][75] = 9'b111111111;
assign micromatrizz[47][76] = 9'b111111111;
assign micromatrizz[47][77] = 9'b111111111;
assign micromatrizz[47][78] = 9'b111111111;
assign micromatrizz[47][79] = 9'b111111111;
assign micromatrizz[47][80] = 9'b111111111;
assign micromatrizz[47][81] = 9'b111111111;
assign micromatrizz[47][82] = 9'b111111111;
assign micromatrizz[47][83] = 9'b111111111;
assign micromatrizz[47][84] = 9'b111111111;
assign micromatrizz[47][85] = 9'b111111111;
assign micromatrizz[47][86] = 9'b111111111;
assign micromatrizz[47][87] = 9'b111111111;
assign micromatrizz[47][88] = 9'b111111111;
assign micromatrizz[47][89] = 9'b111111111;
assign micromatrizz[47][90] = 9'b111111111;
assign micromatrizz[47][91] = 9'b111111111;
assign micromatrizz[47][92] = 9'b111111111;
assign micromatrizz[47][93] = 9'b111111111;
assign micromatrizz[47][94] = 9'b111111111;
assign micromatrizz[47][95] = 9'b111111111;
assign micromatrizz[47][96] = 9'b111111111;
assign micromatrizz[47][97] = 9'b111111111;
assign micromatrizz[47][98] = 9'b111111111;
assign micromatrizz[47][99] = 9'b111111111;
assign micromatrizz[47][100] = 9'b111111111;
assign micromatrizz[47][101] = 9'b111111111;
assign micromatrizz[47][102] = 9'b111111111;
assign micromatrizz[47][103] = 9'b111111111;
assign micromatrizz[47][104] = 9'b111111111;
assign micromatrizz[47][105] = 9'b111111111;
assign micromatrizz[47][106] = 9'b111111111;
assign micromatrizz[47][107] = 9'b111111111;
assign micromatrizz[47][108] = 9'b111111111;
assign micromatrizz[47][109] = 9'b111111111;
assign micromatrizz[47][110] = 9'b111111111;
assign micromatrizz[47][111] = 9'b111111111;
assign micromatrizz[47][112] = 9'b111111111;
assign micromatrizz[47][113] = 9'b111111111;
assign micromatrizz[47][114] = 9'b111111111;
assign micromatrizz[47][115] = 9'b111111111;
assign micromatrizz[47][116] = 9'b111111111;
assign micromatrizz[47][117] = 9'b111111111;
assign micromatrizz[47][118] = 9'b111111111;
assign micromatrizz[47][119] = 9'b111111111;
assign micromatrizz[47][120] = 9'b111111111;
assign micromatrizz[47][121] = 9'b111111111;
assign micromatrizz[47][122] = 9'b111111111;
assign micromatrizz[47][123] = 9'b111111111;
assign micromatrizz[47][124] = 9'b111111111;
assign micromatrizz[47][125] = 9'b111111111;
assign micromatrizz[47][126] = 9'b111111111;
assign micromatrizz[47][127] = 9'b111111111;
assign micromatrizz[47][128] = 9'b111111111;
assign micromatrizz[47][129] = 9'b111111111;
assign micromatrizz[47][130] = 9'b111111111;
assign micromatrizz[47][131] = 9'b111111111;
assign micromatrizz[47][132] = 9'b111111111;
assign micromatrizz[47][133] = 9'b111111111;
assign micromatrizz[47][134] = 9'b111111111;
assign micromatrizz[47][135] = 9'b111111111;
assign micromatrizz[47][136] = 9'b111111111;
assign micromatrizz[47][137] = 9'b111111111;
assign micromatrizz[47][138] = 9'b111111111;
assign micromatrizz[47][139] = 9'b111111111;
assign micromatrizz[47][140] = 9'b111111111;
assign micromatrizz[47][141] = 9'b111111111;
assign micromatrizz[47][142] = 9'b111111111;
assign micromatrizz[47][143] = 9'b111111111;
assign micromatrizz[47][144] = 9'b111111111;
assign micromatrizz[47][145] = 9'b111110010;
assign micromatrizz[47][146] = 9'b111110010;
assign micromatrizz[47][147] = 9'b111110010;
assign micromatrizz[47][148] = 9'b111110011;
assign micromatrizz[47][149] = 9'b111110011;
assign micromatrizz[47][150] = 9'b111110011;
assign micromatrizz[47][151] = 9'b111110010;
assign micromatrizz[47][152] = 9'b111110010;
assign micromatrizz[47][153] = 9'b111110111;
assign micromatrizz[47][154] = 9'b111111111;
assign micromatrizz[47][155] = 9'b111111111;
assign micromatrizz[47][156] = 9'b111111111;
assign micromatrizz[47][157] = 9'b111111111;
assign micromatrizz[47][158] = 9'b111111111;
assign micromatrizz[47][159] = 9'b111111111;
assign micromatrizz[47][160] = 9'b111111111;
assign micromatrizz[47][161] = 9'b111111111;
assign micromatrizz[47][162] = 9'b111111111;
assign micromatrizz[47][163] = 9'b111111111;
assign micromatrizz[47][164] = 9'b111111111;
assign micromatrizz[47][165] = 9'b111111111;
assign micromatrizz[47][166] = 9'b111111111;
assign micromatrizz[47][167] = 9'b111111111;
assign micromatrizz[47][168] = 9'b111111111;
assign micromatrizz[47][169] = 9'b111111111;
assign micromatrizz[47][170] = 9'b111111111;
assign micromatrizz[47][171] = 9'b111111111;
assign micromatrizz[47][172] = 9'b111111111;
assign micromatrizz[47][173] = 9'b111111111;
assign micromatrizz[47][174] = 9'b111111111;
assign micromatrizz[47][175] = 9'b111111111;
assign micromatrizz[47][176] = 9'b111111111;
assign micromatrizz[47][177] = 9'b111111111;
assign micromatrizz[47][178] = 9'b111111111;
assign micromatrizz[47][179] = 9'b111111111;
assign micromatrizz[47][180] = 9'b111111111;
assign micromatrizz[47][181] = 9'b111111111;
assign micromatrizz[47][182] = 9'b111111111;
assign micromatrizz[47][183] = 9'b111111111;
assign micromatrizz[47][184] = 9'b111111111;
assign micromatrizz[47][185] = 9'b111111111;
assign micromatrizz[47][186] = 9'b111111111;
assign micromatrizz[47][187] = 9'b111111111;
assign micromatrizz[47][188] = 9'b111111111;
assign micromatrizz[47][189] = 9'b111111111;
assign micromatrizz[47][190] = 9'b111111111;
assign micromatrizz[47][191] = 9'b111111111;
assign micromatrizz[47][192] = 9'b111111111;
assign micromatrizz[47][193] = 9'b111111111;
assign micromatrizz[47][194] = 9'b111111111;
assign micromatrizz[47][195] = 9'b111111111;
assign micromatrizz[47][196] = 9'b111110111;
assign micromatrizz[47][197] = 9'b111110111;
assign micromatrizz[47][198] = 9'b111110111;
assign micromatrizz[47][199] = 9'b111110111;
assign micromatrizz[47][200] = 9'b111110111;
assign micromatrizz[47][201] = 9'b111110111;
assign micromatrizz[47][202] = 9'b111111111;
assign micromatrizz[47][203] = 9'b111111111;
assign micromatrizz[47][204] = 9'b111111111;
assign micromatrizz[47][205] = 9'b111111111;
assign micromatrizz[47][206] = 9'b111111111;
assign micromatrizz[47][207] = 9'b111111111;
assign micromatrizz[47][208] = 9'b111111111;
assign micromatrizz[47][209] = 9'b111111111;
assign micromatrizz[47][210] = 9'b111111111;
assign micromatrizz[47][211] = 9'b111111111;
assign micromatrizz[47][212] = 9'b111111111;
assign micromatrizz[47][213] = 9'b111111111;
assign micromatrizz[47][214] = 9'b111111111;
assign micromatrizz[47][215] = 9'b111111111;
assign micromatrizz[47][216] = 9'b111111111;
assign micromatrizz[47][217] = 9'b111111111;
assign micromatrizz[47][218] = 9'b111111111;
assign micromatrizz[47][219] = 9'b111111111;
assign micromatrizz[47][220] = 9'b111111111;
assign micromatrizz[47][221] = 9'b111111111;
assign micromatrizz[47][222] = 9'b111111111;
assign micromatrizz[47][223] = 9'b111111111;
assign micromatrizz[47][224] = 9'b111111111;
assign micromatrizz[47][225] = 9'b111111111;
assign micromatrizz[47][226] = 9'b111111111;
assign micromatrizz[47][227] = 9'b111111111;
assign micromatrizz[47][228] = 9'b111111111;
assign micromatrizz[47][229] = 9'b111111111;
assign micromatrizz[47][230] = 9'b111111111;
assign micromatrizz[47][231] = 9'b111111111;
assign micromatrizz[47][232] = 9'b111111111;
assign micromatrizz[47][233] = 9'b111111111;
assign micromatrizz[47][234] = 9'b111111111;
assign micromatrizz[47][235] = 9'b111111111;
assign micromatrizz[47][236] = 9'b111111111;
assign micromatrizz[47][237] = 9'b111111111;
assign micromatrizz[47][238] = 9'b111111111;
assign micromatrizz[47][239] = 9'b111111111;
assign micromatrizz[47][240] = 9'b111111111;
assign micromatrizz[47][241] = 9'b111111111;
assign micromatrizz[47][242] = 9'b111111111;
assign micromatrizz[47][243] = 9'b111111111;
assign micromatrizz[47][244] = 9'b111111111;
assign micromatrizz[47][245] = 9'b111111111;
assign micromatrizz[47][246] = 9'b111111111;
assign micromatrizz[47][247] = 9'b111111111;
assign micromatrizz[47][248] = 9'b111111111;
assign micromatrizz[47][249] = 9'b111111111;
assign micromatrizz[47][250] = 9'b111111111;
assign micromatrizz[47][251] = 9'b111111111;
assign micromatrizz[47][252] = 9'b111111111;
assign micromatrizz[47][253] = 9'b111111111;
assign micromatrizz[47][254] = 9'b111111111;
assign micromatrizz[47][255] = 9'b111111111;
assign micromatrizz[47][256] = 9'b111111111;
assign micromatrizz[47][257] = 9'b111111111;
assign micromatrizz[47][258] = 9'b111111111;
assign micromatrizz[47][259] = 9'b111111111;
assign micromatrizz[47][260] = 9'b111111111;
assign micromatrizz[47][261] = 9'b111111111;
assign micromatrizz[47][262] = 9'b111111111;
assign micromatrizz[47][263] = 9'b111111111;
assign micromatrizz[47][264] = 9'b111111111;
assign micromatrizz[47][265] = 9'b111111111;
assign micromatrizz[47][266] = 9'b111111111;
assign micromatrizz[47][267] = 9'b111111111;
assign micromatrizz[47][268] = 9'b111111111;
assign micromatrizz[47][269] = 9'b111111111;
assign micromatrizz[47][270] = 9'b111111111;
assign micromatrizz[47][271] = 9'b111111111;
assign micromatrizz[47][272] = 9'b111111111;
assign micromatrizz[47][273] = 9'b111111111;
assign micromatrizz[47][274] = 9'b111111111;
assign micromatrizz[47][275] = 9'b111111111;
assign micromatrizz[47][276] = 9'b111111111;
assign micromatrizz[47][277] = 9'b111111111;
assign micromatrizz[47][278] = 9'b111111111;
assign micromatrizz[47][279] = 9'b111111111;
assign micromatrizz[47][280] = 9'b111111111;
assign micromatrizz[47][281] = 9'b111111111;
assign micromatrizz[47][282] = 9'b111111111;
assign micromatrizz[47][283] = 9'b111111111;
assign micromatrizz[47][284] = 9'b111111111;
assign micromatrizz[47][285] = 9'b111111111;
assign micromatrizz[47][286] = 9'b111111111;
assign micromatrizz[47][287] = 9'b111111111;
assign micromatrizz[47][288] = 9'b111111111;
assign micromatrizz[47][289] = 9'b111111111;
assign micromatrizz[47][290] = 9'b111111111;
assign micromatrizz[47][291] = 9'b111111111;
assign micromatrizz[47][292] = 9'b111111111;
assign micromatrizz[47][293] = 9'b111111111;
assign micromatrizz[47][294] = 9'b111111111;
assign micromatrizz[47][295] = 9'b111111111;
assign micromatrizz[47][296] = 9'b111111111;
assign micromatrizz[47][297] = 9'b111111111;
assign micromatrizz[47][298] = 9'b111111111;
assign micromatrizz[47][299] = 9'b111111111;
assign micromatrizz[47][300] = 9'b111111111;
assign micromatrizz[47][301] = 9'b111111111;
assign micromatrizz[47][302] = 9'b111111111;
assign micromatrizz[47][303] = 9'b111111111;
assign micromatrizz[47][304] = 9'b111111111;
assign micromatrizz[47][305] = 9'b111111111;
assign micromatrizz[47][306] = 9'b111111111;
assign micromatrizz[47][307] = 9'b111111111;
assign micromatrizz[47][308] = 9'b111111111;
assign micromatrizz[47][309] = 9'b111111111;
assign micromatrizz[47][310] = 9'b111111111;
assign micromatrizz[47][311] = 9'b111111111;
assign micromatrizz[47][312] = 9'b111111111;
assign micromatrizz[47][313] = 9'b111111111;
assign micromatrizz[47][314] = 9'b111111111;
assign micromatrizz[47][315] = 9'b111111111;
assign micromatrizz[47][316] = 9'b111111111;
assign micromatrizz[47][317] = 9'b111111111;
assign micromatrizz[47][318] = 9'b111111111;
assign micromatrizz[47][319] = 9'b111111111;
assign micromatrizz[47][320] = 9'b111111111;
assign micromatrizz[47][321] = 9'b111111111;
assign micromatrizz[47][322] = 9'b111111111;
assign micromatrizz[47][323] = 9'b111111111;
assign micromatrizz[47][324] = 9'b111111111;
assign micromatrizz[47][325] = 9'b111111111;
assign micromatrizz[47][326] = 9'b111111111;
assign micromatrizz[47][327] = 9'b111111111;
assign micromatrizz[47][328] = 9'b111111111;
assign micromatrizz[47][329] = 9'b111111111;
assign micromatrizz[47][330] = 9'b111111111;
assign micromatrizz[47][331] = 9'b111111111;
assign micromatrizz[47][332] = 9'b111111111;
assign micromatrizz[47][333] = 9'b111111111;
assign micromatrizz[47][334] = 9'b111111111;
assign micromatrizz[47][335] = 9'b111111111;
assign micromatrizz[47][336] = 9'b111111111;
assign micromatrizz[47][337] = 9'b111111111;
assign micromatrizz[47][338] = 9'b111111111;
assign micromatrizz[47][339] = 9'b111111111;
assign micromatrizz[47][340] = 9'b111111111;
assign micromatrizz[47][341] = 9'b111111111;
assign micromatrizz[47][342] = 9'b111111111;
assign micromatrizz[47][343] = 9'b111111111;
assign micromatrizz[47][344] = 9'b111111111;
assign micromatrizz[47][345] = 9'b111111111;
assign micromatrizz[47][346] = 9'b111111111;
assign micromatrizz[47][347] = 9'b111111111;
assign micromatrizz[47][348] = 9'b111111111;
assign micromatrizz[47][349] = 9'b111111111;
assign micromatrizz[47][350] = 9'b111111111;
assign micromatrizz[47][351] = 9'b111111111;
assign micromatrizz[47][352] = 9'b111111111;
assign micromatrizz[47][353] = 9'b111111111;
assign micromatrizz[47][354] = 9'b111111111;
assign micromatrizz[47][355] = 9'b111111111;
assign micromatrizz[47][356] = 9'b111111111;
assign micromatrizz[47][357] = 9'b111111111;
assign micromatrizz[47][358] = 9'b111111111;
assign micromatrizz[47][359] = 9'b111111111;
assign micromatrizz[47][360] = 9'b111111111;
assign micromatrizz[47][361] = 9'b111111111;
assign micromatrizz[47][362] = 9'b111111111;
assign micromatrizz[47][363] = 9'b111111111;
assign micromatrizz[47][364] = 9'b111110111;
assign micromatrizz[47][365] = 9'b111110010;
assign micromatrizz[47][366] = 9'b111111111;
assign micromatrizz[47][367] = 9'b111111111;
assign micromatrizz[47][368] = 9'b111111111;
assign micromatrizz[47][369] = 9'b111111111;
assign micromatrizz[47][370] = 9'b111111111;
assign micromatrizz[47][371] = 9'b111111111;
assign micromatrizz[47][372] = 9'b111111111;
assign micromatrizz[47][373] = 9'b111111111;
assign micromatrizz[47][374] = 9'b111111111;
assign micromatrizz[47][375] = 9'b111111111;
assign micromatrizz[47][376] = 9'b111111111;
assign micromatrizz[47][377] = 9'b111111111;
assign micromatrizz[47][378] = 9'b111111111;
assign micromatrizz[47][379] = 9'b111111111;
assign micromatrizz[47][380] = 9'b111111111;
assign micromatrizz[47][381] = 9'b111111111;
assign micromatrizz[47][382] = 9'b111111111;
assign micromatrizz[47][383] = 9'b111111111;
assign micromatrizz[47][384] = 9'b111111111;
assign micromatrizz[47][385] = 9'b111111111;
assign micromatrizz[47][386] = 9'b111111111;
assign micromatrizz[47][387] = 9'b111111111;
assign micromatrizz[47][388] = 9'b111111111;
assign micromatrizz[47][389] = 9'b111111111;
assign micromatrizz[47][390] = 9'b111111111;
assign micromatrizz[47][391] = 9'b111111111;
assign micromatrizz[47][392] = 9'b111111111;
assign micromatrizz[47][393] = 9'b111111111;
assign micromatrizz[47][394] = 9'b111111111;
assign micromatrizz[47][395] = 9'b111111111;
assign micromatrizz[47][396] = 9'b111111111;
assign micromatrizz[47][397] = 9'b111111111;
assign micromatrizz[47][398] = 9'b111111111;
assign micromatrizz[47][399] = 9'b111111111;
assign micromatrizz[47][400] = 9'b111111111;
assign micromatrizz[47][401] = 9'b111111111;
assign micromatrizz[47][402] = 9'b111111111;
assign micromatrizz[47][403] = 9'b111111111;
assign micromatrizz[47][404] = 9'b111111111;
assign micromatrizz[47][405] = 9'b111111111;
assign micromatrizz[47][406] = 9'b111111111;
assign micromatrizz[47][407] = 9'b111111111;
assign micromatrizz[47][408] = 9'b111111111;
assign micromatrizz[47][409] = 9'b111111111;
assign micromatrizz[47][410] = 9'b111111111;
assign micromatrizz[47][411] = 9'b111111111;
assign micromatrizz[47][412] = 9'b111111111;
assign micromatrizz[47][413] = 9'b111111111;
assign micromatrizz[47][414] = 9'b111111111;
assign micromatrizz[47][415] = 9'b111111111;
assign micromatrizz[47][416] = 9'b111111111;
assign micromatrizz[47][417] = 9'b111111111;
assign micromatrizz[47][418] = 9'b111111111;
assign micromatrizz[47][419] = 9'b111111111;
assign micromatrizz[47][420] = 9'b111111111;
assign micromatrizz[47][421] = 9'b111111111;
assign micromatrizz[47][422] = 9'b111111111;
assign micromatrizz[47][423] = 9'b111111111;
assign micromatrizz[47][424] = 9'b111111111;
assign micromatrizz[47][425] = 9'b111111111;
assign micromatrizz[47][426] = 9'b111111111;
assign micromatrizz[47][427] = 9'b111111111;
assign micromatrizz[47][428] = 9'b111111111;
assign micromatrizz[47][429] = 9'b111111111;
assign micromatrizz[47][430] = 9'b111111111;
assign micromatrizz[47][431] = 9'b111111111;
assign micromatrizz[47][432] = 9'b111111111;
assign micromatrizz[47][433] = 9'b111111111;
assign micromatrizz[47][434] = 9'b111111111;
assign micromatrizz[47][435] = 9'b111111111;
assign micromatrizz[47][436] = 9'b111111111;
assign micromatrizz[47][437] = 9'b111111111;
assign micromatrizz[47][438] = 9'b111111111;
assign micromatrizz[47][439] = 9'b111111111;
assign micromatrizz[47][440] = 9'b111111111;
assign micromatrizz[47][441] = 9'b111111111;
assign micromatrizz[47][442] = 9'b111111111;
assign micromatrizz[47][443] = 9'b111111111;
assign micromatrizz[47][444] = 9'b111111111;
assign micromatrizz[47][445] = 9'b111111111;
assign micromatrizz[47][446] = 9'b111111111;
assign micromatrizz[47][447] = 9'b111111111;
assign micromatrizz[47][448] = 9'b111111111;
assign micromatrizz[47][449] = 9'b111111111;
assign micromatrizz[47][450] = 9'b111111111;
assign micromatrizz[47][451] = 9'b111111111;
assign micromatrizz[47][452] = 9'b111111111;
assign micromatrizz[47][453] = 9'b111111111;
assign micromatrizz[47][454] = 9'b111111111;
assign micromatrizz[47][455] = 9'b111111111;
assign micromatrizz[47][456] = 9'b111111111;
assign micromatrizz[47][457] = 9'b111111111;
assign micromatrizz[47][458] = 9'b111111111;
assign micromatrizz[47][459] = 9'b111111111;
assign micromatrizz[47][460] = 9'b111111111;
assign micromatrizz[47][461] = 9'b111111111;
assign micromatrizz[47][462] = 9'b111111111;
assign micromatrizz[47][463] = 9'b111111111;
assign micromatrizz[47][464] = 9'b111111111;
assign micromatrizz[47][465] = 9'b111111111;
assign micromatrizz[47][466] = 9'b111111111;
assign micromatrizz[47][467] = 9'b111111111;
assign micromatrizz[47][468] = 9'b111111111;
assign micromatrizz[47][469] = 9'b111111111;
assign micromatrizz[47][470] = 9'b111111111;
assign micromatrizz[47][471] = 9'b111111111;
assign micromatrizz[47][472] = 9'b111111111;
assign micromatrizz[47][473] = 9'b111111111;
assign micromatrizz[47][474] = 9'b111111111;
assign micromatrizz[47][475] = 9'b111111111;
assign micromatrizz[47][476] = 9'b111111111;
assign micromatrizz[47][477] = 9'b111111111;
assign micromatrizz[47][478] = 9'b111111111;
assign micromatrizz[47][479] = 9'b111111111;
assign micromatrizz[47][480] = 9'b111111111;
assign micromatrizz[47][481] = 9'b111111111;
assign micromatrizz[47][482] = 9'b111111111;
assign micromatrizz[47][483] = 9'b111111111;
assign micromatrizz[47][484] = 9'b111111111;
assign micromatrizz[47][485] = 9'b111111111;
assign micromatrizz[47][486] = 9'b111111111;
assign micromatrizz[47][487] = 9'b111111111;
assign micromatrizz[47][488] = 9'b111111111;
assign micromatrizz[47][489] = 9'b111111111;
assign micromatrizz[47][490] = 9'b111111111;
assign micromatrizz[47][491] = 9'b111111111;
assign micromatrizz[47][492] = 9'b111111111;
assign micromatrizz[47][493] = 9'b111111111;
assign micromatrizz[47][494] = 9'b111111111;
assign micromatrizz[47][495] = 9'b111111111;
assign micromatrizz[47][496] = 9'b111111111;
assign micromatrizz[47][497] = 9'b111111111;
assign micromatrizz[47][498] = 9'b111111111;
assign micromatrizz[47][499] = 9'b111111111;
assign micromatrizz[47][500] = 9'b111111111;
assign micromatrizz[47][501] = 9'b111111111;
assign micromatrizz[47][502] = 9'b111111111;
assign micromatrizz[47][503] = 9'b111111111;
assign micromatrizz[47][504] = 9'b111111111;
assign micromatrizz[47][505] = 9'b111111111;
assign micromatrizz[47][506] = 9'b111111111;
assign micromatrizz[47][507] = 9'b111111111;
assign micromatrizz[47][508] = 9'b111111111;
assign micromatrizz[47][509] = 9'b111111111;
assign micromatrizz[47][510] = 9'b111111111;
assign micromatrizz[47][511] = 9'b111111111;
assign micromatrizz[47][512] = 9'b111111111;
assign micromatrizz[47][513] = 9'b111111111;
assign micromatrizz[47][514] = 9'b111111111;
assign micromatrizz[47][515] = 9'b111111111;
assign micromatrizz[47][516] = 9'b111111111;
assign micromatrizz[47][517] = 9'b111110111;
assign micromatrizz[47][518] = 9'b111110111;
assign micromatrizz[47][519] = 9'b111110111;
assign micromatrizz[47][520] = 9'b111111111;
assign micromatrizz[47][521] = 9'b111110111;
assign micromatrizz[47][522] = 9'b111110111;
assign micromatrizz[47][523] = 9'b111111111;
assign micromatrizz[47][524] = 9'b111111111;
assign micromatrizz[47][525] = 9'b111111111;
assign micromatrizz[47][526] = 9'b111111111;
assign micromatrizz[47][527] = 9'b111111111;
assign micromatrizz[47][528] = 9'b111111111;
assign micromatrizz[47][529] = 9'b111111111;
assign micromatrizz[47][530] = 9'b111111111;
assign micromatrizz[47][531] = 9'b111111111;
assign micromatrizz[47][532] = 9'b111111111;
assign micromatrizz[47][533] = 9'b111111111;
assign micromatrizz[47][534] = 9'b111111111;
assign micromatrizz[47][535] = 9'b111111111;
assign micromatrizz[47][536] = 9'b111111111;
assign micromatrizz[47][537] = 9'b111111111;
assign micromatrizz[47][538] = 9'b111111111;
assign micromatrizz[47][539] = 9'b111111111;
assign micromatrizz[47][540] = 9'b111111111;
assign micromatrizz[47][541] = 9'b111111111;
assign micromatrizz[47][542] = 9'b111111111;
assign micromatrizz[47][543] = 9'b111111111;
assign micromatrizz[47][544] = 9'b111111111;
assign micromatrizz[47][545] = 9'b111111111;
assign micromatrizz[47][546] = 9'b111111111;
assign micromatrizz[47][547] = 9'b111111111;
assign micromatrizz[47][548] = 9'b111111111;
assign micromatrizz[47][549] = 9'b111111111;
assign micromatrizz[47][550] = 9'b111111111;
assign micromatrizz[47][551] = 9'b111111111;
assign micromatrizz[47][552] = 9'b111111111;
assign micromatrizz[47][553] = 9'b111111111;
assign micromatrizz[47][554] = 9'b111111111;
assign micromatrizz[47][555] = 9'b111111111;
assign micromatrizz[47][556] = 9'b111111111;
assign micromatrizz[47][557] = 9'b111111111;
assign micromatrizz[47][558] = 9'b111110111;
assign micromatrizz[47][559] = 9'b111110111;
assign micromatrizz[47][560] = 9'b111110111;
assign micromatrizz[47][561] = 9'b111110111;
assign micromatrizz[47][562] = 9'b111110111;
assign micromatrizz[47][563] = 9'b111110111;
assign micromatrizz[47][564] = 9'b111110111;
assign micromatrizz[47][565] = 9'b111111111;
assign micromatrizz[47][566] = 9'b111111111;
assign micromatrizz[47][567] = 9'b111111111;
assign micromatrizz[47][568] = 9'b111111111;
assign micromatrizz[47][569] = 9'b111111111;
assign micromatrizz[47][570] = 9'b111111111;
assign micromatrizz[47][571] = 9'b111111111;
assign micromatrizz[47][572] = 9'b111111111;
assign micromatrizz[47][573] = 9'b111111111;
assign micromatrizz[47][574] = 9'b111111111;
assign micromatrizz[47][575] = 9'b111111111;
assign micromatrizz[47][576] = 9'b111111111;
assign micromatrizz[47][577] = 9'b111111111;
assign micromatrizz[47][578] = 9'b111111111;
assign micromatrizz[47][579] = 9'b111111111;
assign micromatrizz[47][580] = 9'b111111111;
assign micromatrizz[47][581] = 9'b111110111;
assign micromatrizz[47][582] = 9'b111110111;
assign micromatrizz[47][583] = 9'b111110111;
assign micromatrizz[47][584] = 9'b111110111;
assign micromatrizz[47][585] = 9'b111110111;
assign micromatrizz[47][586] = 9'b111110111;
assign micromatrizz[47][587] = 9'b111110111;
assign micromatrizz[47][588] = 9'b111111111;
assign micromatrizz[47][589] = 9'b111111111;
assign micromatrizz[47][590] = 9'b111111111;
assign micromatrizz[47][591] = 9'b111111111;
assign micromatrizz[47][592] = 9'b111111111;
assign micromatrizz[47][593] = 9'b111111111;
assign micromatrizz[47][594] = 9'b111111111;
assign micromatrizz[47][595] = 9'b111111111;
assign micromatrizz[47][596] = 9'b111111111;
assign micromatrizz[47][597] = 9'b111111111;
assign micromatrizz[47][598] = 9'b111111111;
assign micromatrizz[47][599] = 9'b111111111;
assign micromatrizz[47][600] = 9'b111111111;
assign micromatrizz[47][601] = 9'b111111111;
assign micromatrizz[47][602] = 9'b111111111;
assign micromatrizz[47][603] = 9'b111111111;
assign micromatrizz[47][604] = 9'b111111111;
assign micromatrizz[47][605] = 9'b111111111;
assign micromatrizz[47][606] = 9'b111111111;
assign micromatrizz[47][607] = 9'b111111111;
assign micromatrizz[47][608] = 9'b111111111;
assign micromatrizz[47][609] = 9'b111111111;
assign micromatrizz[47][610] = 9'b111111111;
assign micromatrizz[47][611] = 9'b111111111;
assign micromatrizz[47][612] = 9'b111111111;
assign micromatrizz[47][613] = 9'b111111111;
assign micromatrizz[47][614] = 9'b111111111;
assign micromatrizz[47][615] = 9'b111111111;
assign micromatrizz[47][616] = 9'b111111111;
assign micromatrizz[47][617] = 9'b111111111;
assign micromatrizz[47][618] = 9'b111111111;
assign micromatrizz[47][619] = 9'b111111111;
assign micromatrizz[47][620] = 9'b111111111;
assign micromatrizz[47][621] = 9'b111111111;
assign micromatrizz[47][622] = 9'b111111111;
assign micromatrizz[47][623] = 9'b111111111;
assign micromatrizz[47][624] = 9'b111111111;
assign micromatrizz[47][625] = 9'b111111111;
assign micromatrizz[47][626] = 9'b111111111;
assign micromatrizz[47][627] = 9'b111111111;
assign micromatrizz[47][628] = 9'b111111111;
assign micromatrizz[47][629] = 9'b111111111;
assign micromatrizz[47][630] = 9'b111111111;
assign micromatrizz[47][631] = 9'b111111111;
assign micromatrizz[47][632] = 9'b111111111;
assign micromatrizz[47][633] = 9'b111111111;
assign micromatrizz[47][634] = 9'b111111111;
assign micromatrizz[47][635] = 9'b111111111;
assign micromatrizz[47][636] = 9'b111111111;
assign micromatrizz[47][637] = 9'b111111111;
assign micromatrizz[47][638] = 9'b111111111;
assign micromatrizz[47][639] = 9'b111111111;
assign micromatrizz[48][0] = 9'b111111111;
assign micromatrizz[48][1] = 9'b111111111;
assign micromatrizz[48][2] = 9'b111111111;
assign micromatrizz[48][3] = 9'b111111111;
assign micromatrizz[48][4] = 9'b111111111;
assign micromatrizz[48][5] = 9'b111111111;
assign micromatrizz[48][6] = 9'b111111111;
assign micromatrizz[48][7] = 9'b111111111;
assign micromatrizz[48][8] = 9'b111111111;
assign micromatrizz[48][9] = 9'b111111111;
assign micromatrizz[48][10] = 9'b111111111;
assign micromatrizz[48][11] = 9'b111111111;
assign micromatrizz[48][12] = 9'b111111111;
assign micromatrizz[48][13] = 9'b111111111;
assign micromatrizz[48][14] = 9'b111111111;
assign micromatrizz[48][15] = 9'b111111111;
assign micromatrizz[48][16] = 9'b111111111;
assign micromatrizz[48][17] = 9'b111111111;
assign micromatrizz[48][18] = 9'b111111111;
assign micromatrizz[48][19] = 9'b111111111;
assign micromatrizz[48][20] = 9'b111111111;
assign micromatrizz[48][21] = 9'b111111111;
assign micromatrizz[48][22] = 9'b111111111;
assign micromatrizz[48][23] = 9'b111111111;
assign micromatrizz[48][24] = 9'b111111111;
assign micromatrizz[48][25] = 9'b111111111;
assign micromatrizz[48][26] = 9'b111111111;
assign micromatrizz[48][27] = 9'b111111111;
assign micromatrizz[48][28] = 9'b111111111;
assign micromatrizz[48][29] = 9'b111111111;
assign micromatrizz[48][30] = 9'b111111111;
assign micromatrizz[48][31] = 9'b111111111;
assign micromatrizz[48][32] = 9'b111111111;
assign micromatrizz[48][33] = 9'b111111111;
assign micromatrizz[48][34] = 9'b111111111;
assign micromatrizz[48][35] = 9'b111111111;
assign micromatrizz[48][36] = 9'b111111111;
assign micromatrizz[48][37] = 9'b111111111;
assign micromatrizz[48][38] = 9'b111111111;
assign micromatrizz[48][39] = 9'b111111111;
assign micromatrizz[48][40] = 9'b111111111;
assign micromatrizz[48][41] = 9'b111111111;
assign micromatrizz[48][42] = 9'b111111111;
assign micromatrizz[48][43] = 9'b111111111;
assign micromatrizz[48][44] = 9'b111111111;
assign micromatrizz[48][45] = 9'b111111111;
assign micromatrizz[48][46] = 9'b111111111;
assign micromatrizz[48][47] = 9'b111111111;
assign micromatrizz[48][48] = 9'b111111111;
assign micromatrizz[48][49] = 9'b111111111;
assign micromatrizz[48][50] = 9'b111111111;
assign micromatrizz[48][51] = 9'b111111111;
assign micromatrizz[48][52] = 9'b111111111;
assign micromatrizz[48][53] = 9'b111111111;
assign micromatrizz[48][54] = 9'b111111111;
assign micromatrizz[48][55] = 9'b111111111;
assign micromatrizz[48][56] = 9'b111111111;
assign micromatrizz[48][57] = 9'b111111111;
assign micromatrizz[48][58] = 9'b111111111;
assign micromatrizz[48][59] = 9'b111111111;
assign micromatrizz[48][60] = 9'b111111111;
assign micromatrizz[48][61] = 9'b111111111;
assign micromatrizz[48][62] = 9'b111111111;
assign micromatrizz[48][63] = 9'b111111111;
assign micromatrizz[48][64] = 9'b111111111;
assign micromatrizz[48][65] = 9'b111111111;
assign micromatrizz[48][66] = 9'b111111111;
assign micromatrizz[48][67] = 9'b111111111;
assign micromatrizz[48][68] = 9'b111111111;
assign micromatrizz[48][69] = 9'b111111111;
assign micromatrizz[48][70] = 9'b111111111;
assign micromatrizz[48][71] = 9'b111111111;
assign micromatrizz[48][72] = 9'b111111111;
assign micromatrizz[48][73] = 9'b111111111;
assign micromatrizz[48][74] = 9'b111111111;
assign micromatrizz[48][75] = 9'b111111111;
assign micromatrizz[48][76] = 9'b111111111;
assign micromatrizz[48][77] = 9'b111111111;
assign micromatrizz[48][78] = 9'b111111111;
assign micromatrizz[48][79] = 9'b111111111;
assign micromatrizz[48][80] = 9'b111111111;
assign micromatrizz[48][81] = 9'b111111111;
assign micromatrizz[48][82] = 9'b111111111;
assign micromatrizz[48][83] = 9'b111111111;
assign micromatrizz[48][84] = 9'b111111111;
assign micromatrizz[48][85] = 9'b111111111;
assign micromatrizz[48][86] = 9'b111111111;
assign micromatrizz[48][87] = 9'b111111111;
assign micromatrizz[48][88] = 9'b111111111;
assign micromatrizz[48][89] = 9'b111111111;
assign micromatrizz[48][90] = 9'b111111111;
assign micromatrizz[48][91] = 9'b111111111;
assign micromatrizz[48][92] = 9'b111111111;
assign micromatrizz[48][93] = 9'b111111111;
assign micromatrizz[48][94] = 9'b111111111;
assign micromatrizz[48][95] = 9'b111111111;
assign micromatrizz[48][96] = 9'b111111111;
assign micromatrizz[48][97] = 9'b111111111;
assign micromatrizz[48][98] = 9'b111111111;
assign micromatrizz[48][99] = 9'b111111111;
assign micromatrizz[48][100] = 9'b111111111;
assign micromatrizz[48][101] = 9'b111111111;
assign micromatrizz[48][102] = 9'b111111111;
assign micromatrizz[48][103] = 9'b111111111;
assign micromatrizz[48][104] = 9'b111111111;
assign micromatrizz[48][105] = 9'b111111111;
assign micromatrizz[48][106] = 9'b111111111;
assign micromatrizz[48][107] = 9'b111111111;
assign micromatrizz[48][108] = 9'b111111111;
assign micromatrizz[48][109] = 9'b111111111;
assign micromatrizz[48][110] = 9'b111111111;
assign micromatrizz[48][111] = 9'b111111111;
assign micromatrizz[48][112] = 9'b111111111;
assign micromatrizz[48][113] = 9'b111111111;
assign micromatrizz[48][114] = 9'b111111111;
assign micromatrizz[48][115] = 9'b111111111;
assign micromatrizz[48][116] = 9'b111111111;
assign micromatrizz[48][117] = 9'b111111111;
assign micromatrizz[48][118] = 9'b111111111;
assign micromatrizz[48][119] = 9'b111111111;
assign micromatrizz[48][120] = 9'b111111111;
assign micromatrizz[48][121] = 9'b111111111;
assign micromatrizz[48][122] = 9'b111111111;
assign micromatrizz[48][123] = 9'b111111111;
assign micromatrizz[48][124] = 9'b111111111;
assign micromatrizz[48][125] = 9'b111111111;
assign micromatrizz[48][126] = 9'b111111111;
assign micromatrizz[48][127] = 9'b111111111;
assign micromatrizz[48][128] = 9'b111111111;
assign micromatrizz[48][129] = 9'b111111111;
assign micromatrizz[48][130] = 9'b111111111;
assign micromatrizz[48][131] = 9'b111111111;
assign micromatrizz[48][132] = 9'b111111111;
assign micromatrizz[48][133] = 9'b111111111;
assign micromatrizz[48][134] = 9'b111111111;
assign micromatrizz[48][135] = 9'b111111111;
assign micromatrizz[48][136] = 9'b111111111;
assign micromatrizz[48][137] = 9'b111111111;
assign micromatrizz[48][138] = 9'b111111111;
assign micromatrizz[48][139] = 9'b111111111;
assign micromatrizz[48][140] = 9'b111111111;
assign micromatrizz[48][141] = 9'b111111111;
assign micromatrizz[48][142] = 9'b111111111;
assign micromatrizz[48][143] = 9'b111111111;
assign micromatrizz[48][144] = 9'b111110010;
assign micromatrizz[48][145] = 9'b111111111;
assign micromatrizz[48][146] = 9'b111111111;
assign micromatrizz[48][147] = 9'b111110111;
assign micromatrizz[48][148] = 9'b111110011;
assign micromatrizz[48][149] = 9'b111110011;
assign micromatrizz[48][150] = 9'b111110011;
assign micromatrizz[48][151] = 9'b111110011;
assign micromatrizz[48][152] = 9'b111110111;
assign micromatrizz[48][153] = 9'b111111111;
assign micromatrizz[48][154] = 9'b111111111;
assign micromatrizz[48][155] = 9'b111111111;
assign micromatrizz[48][156] = 9'b111111111;
assign micromatrizz[48][157] = 9'b111111111;
assign micromatrizz[48][158] = 9'b111111111;
assign micromatrizz[48][159] = 9'b111111111;
assign micromatrizz[48][160] = 9'b111111111;
assign micromatrizz[48][161] = 9'b111111111;
assign micromatrizz[48][162] = 9'b111111111;
assign micromatrizz[48][163] = 9'b111111111;
assign micromatrizz[48][164] = 9'b111111111;
assign micromatrizz[48][165] = 9'b111111111;
assign micromatrizz[48][166] = 9'b111111111;
assign micromatrizz[48][167] = 9'b111111111;
assign micromatrizz[48][168] = 9'b111111111;
assign micromatrizz[48][169] = 9'b111111111;
assign micromatrizz[48][170] = 9'b111111111;
assign micromatrizz[48][171] = 9'b111111111;
assign micromatrizz[48][172] = 9'b111111111;
assign micromatrizz[48][173] = 9'b111111111;
assign micromatrizz[48][174] = 9'b111111111;
assign micromatrizz[48][175] = 9'b111111111;
assign micromatrizz[48][176] = 9'b111111111;
assign micromatrizz[48][177] = 9'b111111111;
assign micromatrizz[48][178] = 9'b111111111;
assign micromatrizz[48][179] = 9'b111111111;
assign micromatrizz[48][180] = 9'b111111111;
assign micromatrizz[48][181] = 9'b111111111;
assign micromatrizz[48][182] = 9'b111111111;
assign micromatrizz[48][183] = 9'b111111111;
assign micromatrizz[48][184] = 9'b111111111;
assign micromatrizz[48][185] = 9'b111111111;
assign micromatrizz[48][186] = 9'b111111111;
assign micromatrizz[48][187] = 9'b111111111;
assign micromatrizz[48][188] = 9'b111111111;
assign micromatrizz[48][189] = 9'b111111111;
assign micromatrizz[48][190] = 9'b111111111;
assign micromatrizz[48][191] = 9'b111111111;
assign micromatrizz[48][192] = 9'b111111111;
assign micromatrizz[48][193] = 9'b111111111;
assign micromatrizz[48][194] = 9'b111111111;
assign micromatrizz[48][195] = 9'b111110110;
assign micromatrizz[48][196] = 9'b111110010;
assign micromatrizz[48][197] = 9'b111110011;
assign micromatrizz[48][198] = 9'b111110010;
assign micromatrizz[48][199] = 9'b111110010;
assign micromatrizz[48][200] = 9'b111110010;
assign micromatrizz[48][201] = 9'b111110010;
assign micromatrizz[48][202] = 9'b111110111;
assign micromatrizz[48][203] = 9'b111111111;
assign micromatrizz[48][204] = 9'b111111111;
assign micromatrizz[48][205] = 9'b111111111;
assign micromatrizz[48][206] = 9'b111111111;
assign micromatrizz[48][207] = 9'b111111111;
assign micromatrizz[48][208] = 9'b111111111;
assign micromatrizz[48][209] = 9'b111111111;
assign micromatrizz[48][210] = 9'b111111111;
assign micromatrizz[48][211] = 9'b111111111;
assign micromatrizz[48][212] = 9'b111111111;
assign micromatrizz[48][213] = 9'b111111111;
assign micromatrizz[48][214] = 9'b111111111;
assign micromatrizz[48][215] = 9'b111111111;
assign micromatrizz[48][216] = 9'b111111111;
assign micromatrizz[48][217] = 9'b111111111;
assign micromatrizz[48][218] = 9'b111111111;
assign micromatrizz[48][219] = 9'b111111111;
assign micromatrizz[48][220] = 9'b111111111;
assign micromatrizz[48][221] = 9'b111111111;
assign micromatrizz[48][222] = 9'b111111111;
assign micromatrizz[48][223] = 9'b111111111;
assign micromatrizz[48][224] = 9'b111111111;
assign micromatrizz[48][225] = 9'b111111111;
assign micromatrizz[48][226] = 9'b111111111;
assign micromatrizz[48][227] = 9'b111111111;
assign micromatrizz[48][228] = 9'b111111111;
assign micromatrizz[48][229] = 9'b111111111;
assign micromatrizz[48][230] = 9'b111111111;
assign micromatrizz[48][231] = 9'b111111111;
assign micromatrizz[48][232] = 9'b111111111;
assign micromatrizz[48][233] = 9'b111111111;
assign micromatrizz[48][234] = 9'b111111111;
assign micromatrizz[48][235] = 9'b111111111;
assign micromatrizz[48][236] = 9'b111111111;
assign micromatrizz[48][237] = 9'b111111111;
assign micromatrizz[48][238] = 9'b111111111;
assign micromatrizz[48][239] = 9'b111111111;
assign micromatrizz[48][240] = 9'b111111111;
assign micromatrizz[48][241] = 9'b111111111;
assign micromatrizz[48][242] = 9'b111111111;
assign micromatrizz[48][243] = 9'b111111111;
assign micromatrizz[48][244] = 9'b111111111;
assign micromatrizz[48][245] = 9'b111111111;
assign micromatrizz[48][246] = 9'b111111111;
assign micromatrizz[48][247] = 9'b111111111;
assign micromatrizz[48][248] = 9'b111111111;
assign micromatrizz[48][249] = 9'b111111111;
assign micromatrizz[48][250] = 9'b111111111;
assign micromatrizz[48][251] = 9'b111111111;
assign micromatrizz[48][252] = 9'b111111111;
assign micromatrizz[48][253] = 9'b111111111;
assign micromatrizz[48][254] = 9'b111111111;
assign micromatrizz[48][255] = 9'b111111111;
assign micromatrizz[48][256] = 9'b111111111;
assign micromatrizz[48][257] = 9'b111111111;
assign micromatrizz[48][258] = 9'b111111111;
assign micromatrizz[48][259] = 9'b111111111;
assign micromatrizz[48][260] = 9'b111111111;
assign micromatrizz[48][261] = 9'b111111111;
assign micromatrizz[48][262] = 9'b111111111;
assign micromatrizz[48][263] = 9'b111111111;
assign micromatrizz[48][264] = 9'b111111111;
assign micromatrizz[48][265] = 9'b111111111;
assign micromatrizz[48][266] = 9'b111111111;
assign micromatrizz[48][267] = 9'b111111111;
assign micromatrizz[48][268] = 9'b111111111;
assign micromatrizz[48][269] = 9'b111111111;
assign micromatrizz[48][270] = 9'b111111111;
assign micromatrizz[48][271] = 9'b111111111;
assign micromatrizz[48][272] = 9'b111111111;
assign micromatrizz[48][273] = 9'b111111111;
assign micromatrizz[48][274] = 9'b111111111;
assign micromatrizz[48][275] = 9'b111111111;
assign micromatrizz[48][276] = 9'b111111111;
assign micromatrizz[48][277] = 9'b111111111;
assign micromatrizz[48][278] = 9'b111111111;
assign micromatrizz[48][279] = 9'b111111111;
assign micromatrizz[48][280] = 9'b111111111;
assign micromatrizz[48][281] = 9'b111111111;
assign micromatrizz[48][282] = 9'b111111111;
assign micromatrizz[48][283] = 9'b111111111;
assign micromatrizz[48][284] = 9'b111111111;
assign micromatrizz[48][285] = 9'b111111111;
assign micromatrizz[48][286] = 9'b111111111;
assign micromatrizz[48][287] = 9'b111111111;
assign micromatrizz[48][288] = 9'b111111111;
assign micromatrizz[48][289] = 9'b111111111;
assign micromatrizz[48][290] = 9'b111111111;
assign micromatrizz[48][291] = 9'b111111111;
assign micromatrizz[48][292] = 9'b111111111;
assign micromatrizz[48][293] = 9'b111111111;
assign micromatrizz[48][294] = 9'b111111111;
assign micromatrizz[48][295] = 9'b111111111;
assign micromatrizz[48][296] = 9'b111111111;
assign micromatrizz[48][297] = 9'b111111111;
assign micromatrizz[48][298] = 9'b111111111;
assign micromatrizz[48][299] = 9'b111111111;
assign micromatrizz[48][300] = 9'b111111111;
assign micromatrizz[48][301] = 9'b111111111;
assign micromatrizz[48][302] = 9'b111111111;
assign micromatrizz[48][303] = 9'b111111111;
assign micromatrizz[48][304] = 9'b111111111;
assign micromatrizz[48][305] = 9'b111111111;
assign micromatrizz[48][306] = 9'b111111111;
assign micromatrizz[48][307] = 9'b111111111;
assign micromatrizz[48][308] = 9'b111111111;
assign micromatrizz[48][309] = 9'b111111111;
assign micromatrizz[48][310] = 9'b111111111;
assign micromatrizz[48][311] = 9'b111111111;
assign micromatrizz[48][312] = 9'b111111111;
assign micromatrizz[48][313] = 9'b111111111;
assign micromatrizz[48][314] = 9'b111111111;
assign micromatrizz[48][315] = 9'b111111111;
assign micromatrizz[48][316] = 9'b111111111;
assign micromatrizz[48][317] = 9'b111111111;
assign micromatrizz[48][318] = 9'b111111111;
assign micromatrizz[48][319] = 9'b111111111;
assign micromatrizz[48][320] = 9'b111111111;
assign micromatrizz[48][321] = 9'b111111111;
assign micromatrizz[48][322] = 9'b111111111;
assign micromatrizz[48][323] = 9'b111111111;
assign micromatrizz[48][324] = 9'b111111111;
assign micromatrizz[48][325] = 9'b111111111;
assign micromatrizz[48][326] = 9'b111111111;
assign micromatrizz[48][327] = 9'b111111111;
assign micromatrizz[48][328] = 9'b111111111;
assign micromatrizz[48][329] = 9'b111111111;
assign micromatrizz[48][330] = 9'b111111111;
assign micromatrizz[48][331] = 9'b111111111;
assign micromatrizz[48][332] = 9'b111111111;
assign micromatrizz[48][333] = 9'b111111111;
assign micromatrizz[48][334] = 9'b111111111;
assign micromatrizz[48][335] = 9'b111111111;
assign micromatrizz[48][336] = 9'b111111111;
assign micromatrizz[48][337] = 9'b111111111;
assign micromatrizz[48][338] = 9'b111111111;
assign micromatrizz[48][339] = 9'b111111111;
assign micromatrizz[48][340] = 9'b111111111;
assign micromatrizz[48][341] = 9'b111111111;
assign micromatrizz[48][342] = 9'b111111111;
assign micromatrizz[48][343] = 9'b111111111;
assign micromatrizz[48][344] = 9'b111111111;
assign micromatrizz[48][345] = 9'b111111111;
assign micromatrizz[48][346] = 9'b111111111;
assign micromatrizz[48][347] = 9'b111111111;
assign micromatrizz[48][348] = 9'b111111111;
assign micromatrizz[48][349] = 9'b111111111;
assign micromatrizz[48][350] = 9'b111111111;
assign micromatrizz[48][351] = 9'b111111111;
assign micromatrizz[48][352] = 9'b111111111;
assign micromatrizz[48][353] = 9'b111111111;
assign micromatrizz[48][354] = 9'b111111111;
assign micromatrizz[48][355] = 9'b111111111;
assign micromatrizz[48][356] = 9'b111111111;
assign micromatrizz[48][357] = 9'b111111111;
assign micromatrizz[48][358] = 9'b111111111;
assign micromatrizz[48][359] = 9'b111111111;
assign micromatrizz[48][360] = 9'b111111111;
assign micromatrizz[48][361] = 9'b111111111;
assign micromatrizz[48][362] = 9'b111110111;
assign micromatrizz[48][363] = 9'b111110010;
assign micromatrizz[48][364] = 9'b111110011;
assign micromatrizz[48][365] = 9'b111110010;
assign micromatrizz[48][366] = 9'b111111111;
assign micromatrizz[48][367] = 9'b111111111;
assign micromatrizz[48][368] = 9'b111111111;
assign micromatrizz[48][369] = 9'b111111111;
assign micromatrizz[48][370] = 9'b111111111;
assign micromatrizz[48][371] = 9'b111111111;
assign micromatrizz[48][372] = 9'b111111111;
assign micromatrizz[48][373] = 9'b111111111;
assign micromatrizz[48][374] = 9'b111111111;
assign micromatrizz[48][375] = 9'b111111111;
assign micromatrizz[48][376] = 9'b111111111;
assign micromatrizz[48][377] = 9'b111111111;
assign micromatrizz[48][378] = 9'b111111111;
assign micromatrizz[48][379] = 9'b111111111;
assign micromatrizz[48][380] = 9'b111111111;
assign micromatrizz[48][381] = 9'b111111111;
assign micromatrizz[48][382] = 9'b111111111;
assign micromatrizz[48][383] = 9'b111111111;
assign micromatrizz[48][384] = 9'b111111111;
assign micromatrizz[48][385] = 9'b111111111;
assign micromatrizz[48][386] = 9'b111111111;
assign micromatrizz[48][387] = 9'b111111111;
assign micromatrizz[48][388] = 9'b111111111;
assign micromatrizz[48][389] = 9'b111111111;
assign micromatrizz[48][390] = 9'b111111111;
assign micromatrizz[48][391] = 9'b111111111;
assign micromatrizz[48][392] = 9'b111111111;
assign micromatrizz[48][393] = 9'b111111111;
assign micromatrizz[48][394] = 9'b111111111;
assign micromatrizz[48][395] = 9'b111111111;
assign micromatrizz[48][396] = 9'b111111111;
assign micromatrizz[48][397] = 9'b111111111;
assign micromatrizz[48][398] = 9'b111111111;
assign micromatrizz[48][399] = 9'b111111111;
assign micromatrizz[48][400] = 9'b111111111;
assign micromatrizz[48][401] = 9'b111111111;
assign micromatrizz[48][402] = 9'b111111111;
assign micromatrizz[48][403] = 9'b111111111;
assign micromatrizz[48][404] = 9'b111111111;
assign micromatrizz[48][405] = 9'b111111111;
assign micromatrizz[48][406] = 9'b111111111;
assign micromatrizz[48][407] = 9'b111111111;
assign micromatrizz[48][408] = 9'b111111111;
assign micromatrizz[48][409] = 9'b111111111;
assign micromatrizz[48][410] = 9'b111111111;
assign micromatrizz[48][411] = 9'b111111111;
assign micromatrizz[48][412] = 9'b111111111;
assign micromatrizz[48][413] = 9'b111111111;
assign micromatrizz[48][414] = 9'b111111111;
assign micromatrizz[48][415] = 9'b111111111;
assign micromatrizz[48][416] = 9'b111111111;
assign micromatrizz[48][417] = 9'b111111111;
assign micromatrizz[48][418] = 9'b111111111;
assign micromatrizz[48][419] = 9'b111111111;
assign micromatrizz[48][420] = 9'b111111111;
assign micromatrizz[48][421] = 9'b111111111;
assign micromatrizz[48][422] = 9'b111111111;
assign micromatrizz[48][423] = 9'b111111111;
assign micromatrizz[48][424] = 9'b111111111;
assign micromatrizz[48][425] = 9'b111111111;
assign micromatrizz[48][426] = 9'b111111111;
assign micromatrizz[48][427] = 9'b111111111;
assign micromatrizz[48][428] = 9'b111111111;
assign micromatrizz[48][429] = 9'b111111111;
assign micromatrizz[48][430] = 9'b111111111;
assign micromatrizz[48][431] = 9'b111111111;
assign micromatrizz[48][432] = 9'b111111111;
assign micromatrizz[48][433] = 9'b111111111;
assign micromatrizz[48][434] = 9'b111111111;
assign micromatrizz[48][435] = 9'b111111111;
assign micromatrizz[48][436] = 9'b111111111;
assign micromatrizz[48][437] = 9'b111111111;
assign micromatrizz[48][438] = 9'b111111111;
assign micromatrizz[48][439] = 9'b111111111;
assign micromatrizz[48][440] = 9'b111111111;
assign micromatrizz[48][441] = 9'b111111111;
assign micromatrizz[48][442] = 9'b111111111;
assign micromatrizz[48][443] = 9'b111111111;
assign micromatrizz[48][444] = 9'b111111111;
assign micromatrizz[48][445] = 9'b111111111;
assign micromatrizz[48][446] = 9'b111111111;
assign micromatrizz[48][447] = 9'b111111111;
assign micromatrizz[48][448] = 9'b111111111;
assign micromatrizz[48][449] = 9'b111111111;
assign micromatrizz[48][450] = 9'b111111111;
assign micromatrizz[48][451] = 9'b111111111;
assign micromatrizz[48][452] = 9'b111111111;
assign micromatrizz[48][453] = 9'b111111111;
assign micromatrizz[48][454] = 9'b111111111;
assign micromatrizz[48][455] = 9'b111111111;
assign micromatrizz[48][456] = 9'b111111111;
assign micromatrizz[48][457] = 9'b111111111;
assign micromatrizz[48][458] = 9'b111111111;
assign micromatrizz[48][459] = 9'b111111111;
assign micromatrizz[48][460] = 9'b111111111;
assign micromatrizz[48][461] = 9'b111111111;
assign micromatrizz[48][462] = 9'b111111111;
assign micromatrizz[48][463] = 9'b111111111;
assign micromatrizz[48][464] = 9'b111111111;
assign micromatrizz[48][465] = 9'b111111111;
assign micromatrizz[48][466] = 9'b111111111;
assign micromatrizz[48][467] = 9'b111111111;
assign micromatrizz[48][468] = 9'b111111111;
assign micromatrizz[48][469] = 9'b111111111;
assign micromatrizz[48][470] = 9'b111111111;
assign micromatrizz[48][471] = 9'b111111111;
assign micromatrizz[48][472] = 9'b111111111;
assign micromatrizz[48][473] = 9'b111111111;
assign micromatrizz[48][474] = 9'b111111111;
assign micromatrizz[48][475] = 9'b111111111;
assign micromatrizz[48][476] = 9'b111111111;
assign micromatrizz[48][477] = 9'b111111111;
assign micromatrizz[48][478] = 9'b111111111;
assign micromatrizz[48][479] = 9'b111111111;
assign micromatrizz[48][480] = 9'b111111111;
assign micromatrizz[48][481] = 9'b111111111;
assign micromatrizz[48][482] = 9'b111111111;
assign micromatrizz[48][483] = 9'b111111111;
assign micromatrizz[48][484] = 9'b111111111;
assign micromatrizz[48][485] = 9'b111111111;
assign micromatrizz[48][486] = 9'b111111111;
assign micromatrizz[48][487] = 9'b111111111;
assign micromatrizz[48][488] = 9'b111111111;
assign micromatrizz[48][489] = 9'b111111111;
assign micromatrizz[48][490] = 9'b111111111;
assign micromatrizz[48][491] = 9'b111111111;
assign micromatrizz[48][492] = 9'b111111111;
assign micromatrizz[48][493] = 9'b111111111;
assign micromatrizz[48][494] = 9'b111111111;
assign micromatrizz[48][495] = 9'b111111111;
assign micromatrizz[48][496] = 9'b111111111;
assign micromatrizz[48][497] = 9'b111111111;
assign micromatrizz[48][498] = 9'b111111111;
assign micromatrizz[48][499] = 9'b111111111;
assign micromatrizz[48][500] = 9'b111111111;
assign micromatrizz[48][501] = 9'b111111111;
assign micromatrizz[48][502] = 9'b111111111;
assign micromatrizz[48][503] = 9'b111111111;
assign micromatrizz[48][504] = 9'b111111111;
assign micromatrizz[48][505] = 9'b111111111;
assign micromatrizz[48][506] = 9'b111111111;
assign micromatrizz[48][507] = 9'b111111111;
assign micromatrizz[48][508] = 9'b111111111;
assign micromatrizz[48][509] = 9'b111111111;
assign micromatrizz[48][510] = 9'b111111111;
assign micromatrizz[48][511] = 9'b111111111;
assign micromatrizz[48][512] = 9'b111111111;
assign micromatrizz[48][513] = 9'b111111111;
assign micromatrizz[48][514] = 9'b111111111;
assign micromatrizz[48][515] = 9'b111111111;
assign micromatrizz[48][516] = 9'b111110110;
assign micromatrizz[48][517] = 9'b111110010;
assign micromatrizz[48][518] = 9'b111110011;
assign micromatrizz[48][519] = 9'b111110010;
assign micromatrizz[48][520] = 9'b111110010;
assign micromatrizz[48][521] = 9'b111110010;
assign micromatrizz[48][522] = 9'b111110010;
assign micromatrizz[48][523] = 9'b111110111;
assign micromatrizz[48][524] = 9'b111111111;
assign micromatrizz[48][525] = 9'b111111111;
assign micromatrizz[48][526] = 9'b111111111;
assign micromatrizz[48][527] = 9'b111111111;
assign micromatrizz[48][528] = 9'b111111111;
assign micromatrizz[48][529] = 9'b111111111;
assign micromatrizz[48][530] = 9'b111111111;
assign micromatrizz[48][531] = 9'b111111111;
assign micromatrizz[48][532] = 9'b111111111;
assign micromatrizz[48][533] = 9'b111111111;
assign micromatrizz[48][534] = 9'b111111111;
assign micromatrizz[48][535] = 9'b111111111;
assign micromatrizz[48][536] = 9'b111111111;
assign micromatrizz[48][537] = 9'b111111111;
assign micromatrizz[48][538] = 9'b111111111;
assign micromatrizz[48][539] = 9'b111111111;
assign micromatrizz[48][540] = 9'b111111111;
assign micromatrizz[48][541] = 9'b111111111;
assign micromatrizz[48][542] = 9'b111111111;
assign micromatrizz[48][543] = 9'b111111111;
assign micromatrizz[48][544] = 9'b111111111;
assign micromatrizz[48][545] = 9'b111111111;
assign micromatrizz[48][546] = 9'b111111111;
assign micromatrizz[48][547] = 9'b111111111;
assign micromatrizz[48][548] = 9'b111111111;
assign micromatrizz[48][549] = 9'b111111111;
assign micromatrizz[48][550] = 9'b111111111;
assign micromatrizz[48][551] = 9'b111111111;
assign micromatrizz[48][552] = 9'b111111111;
assign micromatrizz[48][553] = 9'b111111111;
assign micromatrizz[48][554] = 9'b111111111;
assign micromatrizz[48][555] = 9'b111111111;
assign micromatrizz[48][556] = 9'b111111111;
assign micromatrizz[48][557] = 9'b111111111;
assign micromatrizz[48][558] = 9'b111110010;
assign micromatrizz[48][559] = 9'b111110010;
assign micromatrizz[48][560] = 9'b111110010;
assign micromatrizz[48][561] = 9'b111110010;
assign micromatrizz[48][562] = 9'b111110010;
assign micromatrizz[48][563] = 9'b111110010;
assign micromatrizz[48][564] = 9'b111110010;
assign micromatrizz[48][565] = 9'b111111111;
assign micromatrizz[48][566] = 9'b111111111;
assign micromatrizz[48][567] = 9'b111111111;
assign micromatrizz[48][568] = 9'b111111111;
assign micromatrizz[48][569] = 9'b111111111;
assign micromatrizz[48][570] = 9'b111111111;
assign micromatrizz[48][571] = 9'b111111111;
assign micromatrizz[48][572] = 9'b111111111;
assign micromatrizz[48][573] = 9'b111111111;
assign micromatrizz[48][574] = 9'b111111111;
assign micromatrizz[48][575] = 9'b111111111;
assign micromatrizz[48][576] = 9'b111111111;
assign micromatrizz[48][577] = 9'b111111111;
assign micromatrizz[48][578] = 9'b111111111;
assign micromatrizz[48][579] = 9'b111111111;
assign micromatrizz[48][580] = 9'b111111111;
assign micromatrizz[48][581] = 9'b111110010;
assign micromatrizz[48][582] = 9'b111110010;
assign micromatrizz[48][583] = 9'b111110010;
assign micromatrizz[48][584] = 9'b111110010;
assign micromatrizz[48][585] = 9'b111110010;
assign micromatrizz[48][586] = 9'b111110011;
assign micromatrizz[48][587] = 9'b111110010;
assign micromatrizz[48][588] = 9'b111110111;
assign micromatrizz[48][589] = 9'b111111111;
assign micromatrizz[48][590] = 9'b111111111;
assign micromatrizz[48][591] = 9'b111111111;
assign micromatrizz[48][592] = 9'b111111111;
assign micromatrizz[48][593] = 9'b111111111;
assign micromatrizz[48][594] = 9'b111111111;
assign micromatrizz[48][595] = 9'b111111111;
assign micromatrizz[48][596] = 9'b111111111;
assign micromatrizz[48][597] = 9'b111111111;
assign micromatrizz[48][598] = 9'b111111111;
assign micromatrizz[48][599] = 9'b111111111;
assign micromatrizz[48][600] = 9'b111111111;
assign micromatrizz[48][601] = 9'b111111111;
assign micromatrizz[48][602] = 9'b111111111;
assign micromatrizz[48][603] = 9'b111111111;
assign micromatrizz[48][604] = 9'b111111111;
assign micromatrizz[48][605] = 9'b111111111;
assign micromatrizz[48][606] = 9'b111111111;
assign micromatrizz[48][607] = 9'b111111111;
assign micromatrizz[48][608] = 9'b111111111;
assign micromatrizz[48][609] = 9'b111111111;
assign micromatrizz[48][610] = 9'b111111111;
assign micromatrizz[48][611] = 9'b111111111;
assign micromatrizz[48][612] = 9'b111111111;
assign micromatrizz[48][613] = 9'b111111111;
assign micromatrizz[48][614] = 9'b111111111;
assign micromatrizz[48][615] = 9'b111111111;
assign micromatrizz[48][616] = 9'b111111111;
assign micromatrizz[48][617] = 9'b111111111;
assign micromatrizz[48][618] = 9'b111111111;
assign micromatrizz[48][619] = 9'b111111111;
assign micromatrizz[48][620] = 9'b111111111;
assign micromatrizz[48][621] = 9'b111111111;
assign micromatrizz[48][622] = 9'b111111111;
assign micromatrizz[48][623] = 9'b111111111;
assign micromatrizz[48][624] = 9'b111111111;
assign micromatrizz[48][625] = 9'b111111111;
assign micromatrizz[48][626] = 9'b111111111;
assign micromatrizz[48][627] = 9'b111111111;
assign micromatrizz[48][628] = 9'b111111111;
assign micromatrizz[48][629] = 9'b111111111;
assign micromatrizz[48][630] = 9'b111111111;
assign micromatrizz[48][631] = 9'b111111111;
assign micromatrizz[48][632] = 9'b111111111;
assign micromatrizz[48][633] = 9'b111111111;
assign micromatrizz[48][634] = 9'b111111111;
assign micromatrizz[48][635] = 9'b111111111;
assign micromatrizz[48][636] = 9'b111111111;
assign micromatrizz[48][637] = 9'b111111111;
assign micromatrizz[48][638] = 9'b111111111;
assign micromatrizz[48][639] = 9'b111111111;
assign micromatrizz[49][0] = 9'b111111111;
assign micromatrizz[49][1] = 9'b111111111;
assign micromatrizz[49][2] = 9'b111111111;
assign micromatrizz[49][3] = 9'b111111111;
assign micromatrizz[49][4] = 9'b111111111;
assign micromatrizz[49][5] = 9'b111111111;
assign micromatrizz[49][6] = 9'b111111111;
assign micromatrizz[49][7] = 9'b111111111;
assign micromatrizz[49][8] = 9'b111111111;
assign micromatrizz[49][9] = 9'b111111111;
assign micromatrizz[49][10] = 9'b111111111;
assign micromatrizz[49][11] = 9'b111111111;
assign micromatrizz[49][12] = 9'b111111111;
assign micromatrizz[49][13] = 9'b111111111;
assign micromatrizz[49][14] = 9'b111111111;
assign micromatrizz[49][15] = 9'b111111111;
assign micromatrizz[49][16] = 9'b111111111;
assign micromatrizz[49][17] = 9'b111111111;
assign micromatrizz[49][18] = 9'b111111111;
assign micromatrizz[49][19] = 9'b111111111;
assign micromatrizz[49][20] = 9'b111111111;
assign micromatrizz[49][21] = 9'b111111111;
assign micromatrizz[49][22] = 9'b111111111;
assign micromatrizz[49][23] = 9'b111111111;
assign micromatrizz[49][24] = 9'b111111111;
assign micromatrizz[49][25] = 9'b111111111;
assign micromatrizz[49][26] = 9'b111111111;
assign micromatrizz[49][27] = 9'b111111111;
assign micromatrizz[49][28] = 9'b111111111;
assign micromatrizz[49][29] = 9'b111111111;
assign micromatrizz[49][30] = 9'b111111111;
assign micromatrizz[49][31] = 9'b111111111;
assign micromatrizz[49][32] = 9'b111111111;
assign micromatrizz[49][33] = 9'b111111111;
assign micromatrizz[49][34] = 9'b111111111;
assign micromatrizz[49][35] = 9'b111111111;
assign micromatrizz[49][36] = 9'b111111111;
assign micromatrizz[49][37] = 9'b111111111;
assign micromatrizz[49][38] = 9'b111111111;
assign micromatrizz[49][39] = 9'b111111111;
assign micromatrizz[49][40] = 9'b111111111;
assign micromatrizz[49][41] = 9'b111111111;
assign micromatrizz[49][42] = 9'b111111111;
assign micromatrizz[49][43] = 9'b111111111;
assign micromatrizz[49][44] = 9'b111111111;
assign micromatrizz[49][45] = 9'b111111111;
assign micromatrizz[49][46] = 9'b111111111;
assign micromatrizz[49][47] = 9'b111111111;
assign micromatrizz[49][48] = 9'b111111111;
assign micromatrizz[49][49] = 9'b111111111;
assign micromatrizz[49][50] = 9'b111111111;
assign micromatrizz[49][51] = 9'b111111111;
assign micromatrizz[49][52] = 9'b111111111;
assign micromatrizz[49][53] = 9'b111111111;
assign micromatrizz[49][54] = 9'b111111111;
assign micromatrizz[49][55] = 9'b111111111;
assign micromatrizz[49][56] = 9'b111111111;
assign micromatrizz[49][57] = 9'b111111111;
assign micromatrizz[49][58] = 9'b111111111;
assign micromatrizz[49][59] = 9'b111111111;
assign micromatrizz[49][60] = 9'b111111111;
assign micromatrizz[49][61] = 9'b111111111;
assign micromatrizz[49][62] = 9'b111111111;
assign micromatrizz[49][63] = 9'b111111111;
assign micromatrizz[49][64] = 9'b111111111;
assign micromatrizz[49][65] = 9'b111111111;
assign micromatrizz[49][66] = 9'b111111111;
assign micromatrizz[49][67] = 9'b111111111;
assign micromatrizz[49][68] = 9'b111111111;
assign micromatrizz[49][69] = 9'b111111111;
assign micromatrizz[49][70] = 9'b111111111;
assign micromatrizz[49][71] = 9'b111111111;
assign micromatrizz[49][72] = 9'b111111111;
assign micromatrizz[49][73] = 9'b111111111;
assign micromatrizz[49][74] = 9'b111111111;
assign micromatrizz[49][75] = 9'b111111111;
assign micromatrizz[49][76] = 9'b111111111;
assign micromatrizz[49][77] = 9'b111111111;
assign micromatrizz[49][78] = 9'b111111111;
assign micromatrizz[49][79] = 9'b111111111;
assign micromatrizz[49][80] = 9'b111111111;
assign micromatrizz[49][81] = 9'b111111111;
assign micromatrizz[49][82] = 9'b111111111;
assign micromatrizz[49][83] = 9'b111111111;
assign micromatrizz[49][84] = 9'b111111111;
assign micromatrizz[49][85] = 9'b111111111;
assign micromatrizz[49][86] = 9'b111111111;
assign micromatrizz[49][87] = 9'b111111111;
assign micromatrizz[49][88] = 9'b111111111;
assign micromatrizz[49][89] = 9'b111111111;
assign micromatrizz[49][90] = 9'b111111111;
assign micromatrizz[49][91] = 9'b111111111;
assign micromatrizz[49][92] = 9'b111111111;
assign micromatrizz[49][93] = 9'b111111111;
assign micromatrizz[49][94] = 9'b111111111;
assign micromatrizz[49][95] = 9'b111111111;
assign micromatrizz[49][96] = 9'b111111111;
assign micromatrizz[49][97] = 9'b111111111;
assign micromatrizz[49][98] = 9'b111111111;
assign micromatrizz[49][99] = 9'b111111111;
assign micromatrizz[49][100] = 9'b111111111;
assign micromatrizz[49][101] = 9'b111111111;
assign micromatrizz[49][102] = 9'b111111111;
assign micromatrizz[49][103] = 9'b111111111;
assign micromatrizz[49][104] = 9'b111111111;
assign micromatrizz[49][105] = 9'b111111111;
assign micromatrizz[49][106] = 9'b111111111;
assign micromatrizz[49][107] = 9'b111111111;
assign micromatrizz[49][108] = 9'b111111111;
assign micromatrizz[49][109] = 9'b111111111;
assign micromatrizz[49][110] = 9'b111111111;
assign micromatrizz[49][111] = 9'b111111111;
assign micromatrizz[49][112] = 9'b111111111;
assign micromatrizz[49][113] = 9'b111111111;
assign micromatrizz[49][114] = 9'b111111111;
assign micromatrizz[49][115] = 9'b111111111;
assign micromatrizz[49][116] = 9'b111111111;
assign micromatrizz[49][117] = 9'b111111111;
assign micromatrizz[49][118] = 9'b111111111;
assign micromatrizz[49][119] = 9'b111111111;
assign micromatrizz[49][120] = 9'b111111111;
assign micromatrizz[49][121] = 9'b111111111;
assign micromatrizz[49][122] = 9'b111111111;
assign micromatrizz[49][123] = 9'b111111111;
assign micromatrizz[49][124] = 9'b111111111;
assign micromatrizz[49][125] = 9'b111111111;
assign micromatrizz[49][126] = 9'b111111111;
assign micromatrizz[49][127] = 9'b111111111;
assign micromatrizz[49][128] = 9'b111111111;
assign micromatrizz[49][129] = 9'b111111111;
assign micromatrizz[49][130] = 9'b111111111;
assign micromatrizz[49][131] = 9'b111111111;
assign micromatrizz[49][132] = 9'b111111111;
assign micromatrizz[49][133] = 9'b111111111;
assign micromatrizz[49][134] = 9'b111111111;
assign micromatrizz[49][135] = 9'b111111111;
assign micromatrizz[49][136] = 9'b111111111;
assign micromatrizz[49][137] = 9'b111111111;
assign micromatrizz[49][138] = 9'b111111111;
assign micromatrizz[49][139] = 9'b111111111;
assign micromatrizz[49][140] = 9'b111111111;
assign micromatrizz[49][141] = 9'b111111111;
assign micromatrizz[49][142] = 9'b111111111;
assign micromatrizz[49][143] = 9'b111110110;
assign micromatrizz[49][144] = 9'b111111111;
assign micromatrizz[49][145] = 9'b111111111;
assign micromatrizz[49][146] = 9'b111111111;
assign micromatrizz[49][147] = 9'b111111111;
assign micromatrizz[49][148] = 9'b111111111;
assign micromatrizz[49][149] = 9'b111111111;
assign micromatrizz[49][150] = 9'b111110111;
assign micromatrizz[49][151] = 9'b111110111;
assign micromatrizz[49][152] = 9'b111111111;
assign micromatrizz[49][153] = 9'b111111111;
assign micromatrizz[49][154] = 9'b111111111;
assign micromatrizz[49][155] = 9'b111111111;
assign micromatrizz[49][156] = 9'b111111111;
assign micromatrizz[49][157] = 9'b111111111;
assign micromatrizz[49][158] = 9'b111111111;
assign micromatrizz[49][159] = 9'b111111111;
assign micromatrizz[49][160] = 9'b111111111;
assign micromatrizz[49][161] = 9'b111111111;
assign micromatrizz[49][162] = 9'b111111111;
assign micromatrizz[49][163] = 9'b111111111;
assign micromatrizz[49][164] = 9'b111111111;
assign micromatrizz[49][165] = 9'b111111111;
assign micromatrizz[49][166] = 9'b111111111;
assign micromatrizz[49][167] = 9'b111111111;
assign micromatrizz[49][168] = 9'b111111111;
assign micromatrizz[49][169] = 9'b111111111;
assign micromatrizz[49][170] = 9'b111111111;
assign micromatrizz[49][171] = 9'b111111111;
assign micromatrizz[49][172] = 9'b111111111;
assign micromatrizz[49][173] = 9'b111111111;
assign micromatrizz[49][174] = 9'b111111111;
assign micromatrizz[49][175] = 9'b111111111;
assign micromatrizz[49][176] = 9'b111111111;
assign micromatrizz[49][177] = 9'b111111111;
assign micromatrizz[49][178] = 9'b111111111;
assign micromatrizz[49][179] = 9'b111111111;
assign micromatrizz[49][180] = 9'b111111111;
assign micromatrizz[49][181] = 9'b111111111;
assign micromatrizz[49][182] = 9'b111111111;
assign micromatrizz[49][183] = 9'b111111111;
assign micromatrizz[49][184] = 9'b111111111;
assign micromatrizz[49][185] = 9'b111111111;
assign micromatrizz[49][186] = 9'b111111111;
assign micromatrizz[49][187] = 9'b111111111;
assign micromatrizz[49][188] = 9'b111111111;
assign micromatrizz[49][189] = 9'b111111111;
assign micromatrizz[49][190] = 9'b111111111;
assign micromatrizz[49][191] = 9'b111111111;
assign micromatrizz[49][192] = 9'b111111111;
assign micromatrizz[49][193] = 9'b111111111;
assign micromatrizz[49][194] = 9'b111111111;
assign micromatrizz[49][195] = 9'b111110010;
assign micromatrizz[49][196] = 9'b111110010;
assign micromatrizz[49][197] = 9'b111110011;
assign micromatrizz[49][198] = 9'b111110011;
assign micromatrizz[49][199] = 9'b111110010;
assign micromatrizz[49][200] = 9'b111110010;
assign micromatrizz[49][201] = 9'b111110011;
assign micromatrizz[49][202] = 9'b111110111;
assign micromatrizz[49][203] = 9'b111111111;
assign micromatrizz[49][204] = 9'b111111111;
assign micromatrizz[49][205] = 9'b111111111;
assign micromatrizz[49][206] = 9'b111111111;
assign micromatrizz[49][207] = 9'b111111111;
assign micromatrizz[49][208] = 9'b111111111;
assign micromatrizz[49][209] = 9'b111111111;
assign micromatrizz[49][210] = 9'b111111111;
assign micromatrizz[49][211] = 9'b111111111;
assign micromatrizz[49][212] = 9'b111111111;
assign micromatrizz[49][213] = 9'b111111111;
assign micromatrizz[49][214] = 9'b111111111;
assign micromatrizz[49][215] = 9'b111111111;
assign micromatrizz[49][216] = 9'b111111111;
assign micromatrizz[49][217] = 9'b111111111;
assign micromatrizz[49][218] = 9'b111111111;
assign micromatrizz[49][219] = 9'b111111111;
assign micromatrizz[49][220] = 9'b111111111;
assign micromatrizz[49][221] = 9'b111111111;
assign micromatrizz[49][222] = 9'b111111111;
assign micromatrizz[49][223] = 9'b111111111;
assign micromatrizz[49][224] = 9'b111111111;
assign micromatrizz[49][225] = 9'b111111111;
assign micromatrizz[49][226] = 9'b111111111;
assign micromatrizz[49][227] = 9'b111111111;
assign micromatrizz[49][228] = 9'b111111111;
assign micromatrizz[49][229] = 9'b111111111;
assign micromatrizz[49][230] = 9'b111111111;
assign micromatrizz[49][231] = 9'b111111111;
assign micromatrizz[49][232] = 9'b111111111;
assign micromatrizz[49][233] = 9'b111111111;
assign micromatrizz[49][234] = 9'b111111111;
assign micromatrizz[49][235] = 9'b111111111;
assign micromatrizz[49][236] = 9'b111111111;
assign micromatrizz[49][237] = 9'b111111111;
assign micromatrizz[49][238] = 9'b111111111;
assign micromatrizz[49][239] = 9'b111111111;
assign micromatrizz[49][240] = 9'b111111111;
assign micromatrizz[49][241] = 9'b111111111;
assign micromatrizz[49][242] = 9'b111111111;
assign micromatrizz[49][243] = 9'b111111111;
assign micromatrizz[49][244] = 9'b111111111;
assign micromatrizz[49][245] = 9'b111111111;
assign micromatrizz[49][246] = 9'b111111111;
assign micromatrizz[49][247] = 9'b111111111;
assign micromatrizz[49][248] = 9'b111111111;
assign micromatrizz[49][249] = 9'b111111111;
assign micromatrizz[49][250] = 9'b111111111;
assign micromatrizz[49][251] = 9'b111111111;
assign micromatrizz[49][252] = 9'b111111111;
assign micromatrizz[49][253] = 9'b111111111;
assign micromatrizz[49][254] = 9'b111111111;
assign micromatrizz[49][255] = 9'b111111111;
assign micromatrizz[49][256] = 9'b111111111;
assign micromatrizz[49][257] = 9'b111111111;
assign micromatrizz[49][258] = 9'b111111111;
assign micromatrizz[49][259] = 9'b111111111;
assign micromatrizz[49][260] = 9'b111111111;
assign micromatrizz[49][261] = 9'b111111111;
assign micromatrizz[49][262] = 9'b111111111;
assign micromatrizz[49][263] = 9'b111111111;
assign micromatrizz[49][264] = 9'b111111111;
assign micromatrizz[49][265] = 9'b111111111;
assign micromatrizz[49][266] = 9'b111111111;
assign micromatrizz[49][267] = 9'b111111111;
assign micromatrizz[49][268] = 9'b111111111;
assign micromatrizz[49][269] = 9'b111111111;
assign micromatrizz[49][270] = 9'b111111111;
assign micromatrizz[49][271] = 9'b111111111;
assign micromatrizz[49][272] = 9'b111111111;
assign micromatrizz[49][273] = 9'b111111111;
assign micromatrizz[49][274] = 9'b111111111;
assign micromatrizz[49][275] = 9'b111111111;
assign micromatrizz[49][276] = 9'b111111111;
assign micromatrizz[49][277] = 9'b111111111;
assign micromatrizz[49][278] = 9'b111111111;
assign micromatrizz[49][279] = 9'b111111111;
assign micromatrizz[49][280] = 9'b111111111;
assign micromatrizz[49][281] = 9'b111111111;
assign micromatrizz[49][282] = 9'b111111111;
assign micromatrizz[49][283] = 9'b111111111;
assign micromatrizz[49][284] = 9'b111111111;
assign micromatrizz[49][285] = 9'b111111111;
assign micromatrizz[49][286] = 9'b111111111;
assign micromatrizz[49][287] = 9'b111111111;
assign micromatrizz[49][288] = 9'b111111111;
assign micromatrizz[49][289] = 9'b111111111;
assign micromatrizz[49][290] = 9'b111111111;
assign micromatrizz[49][291] = 9'b111111111;
assign micromatrizz[49][292] = 9'b111111111;
assign micromatrizz[49][293] = 9'b111111111;
assign micromatrizz[49][294] = 9'b111111111;
assign micromatrizz[49][295] = 9'b111111111;
assign micromatrizz[49][296] = 9'b111111111;
assign micromatrizz[49][297] = 9'b111111111;
assign micromatrizz[49][298] = 9'b111111111;
assign micromatrizz[49][299] = 9'b111111111;
assign micromatrizz[49][300] = 9'b111111111;
assign micromatrizz[49][301] = 9'b111111111;
assign micromatrizz[49][302] = 9'b111111111;
assign micromatrizz[49][303] = 9'b111111111;
assign micromatrizz[49][304] = 9'b111111111;
assign micromatrizz[49][305] = 9'b111111111;
assign micromatrizz[49][306] = 9'b111111111;
assign micromatrizz[49][307] = 9'b111111111;
assign micromatrizz[49][308] = 9'b111111111;
assign micromatrizz[49][309] = 9'b111111111;
assign micromatrizz[49][310] = 9'b111111111;
assign micromatrizz[49][311] = 9'b111111111;
assign micromatrizz[49][312] = 9'b111111111;
assign micromatrizz[49][313] = 9'b111111111;
assign micromatrizz[49][314] = 9'b111111111;
assign micromatrizz[49][315] = 9'b111111111;
assign micromatrizz[49][316] = 9'b111111111;
assign micromatrizz[49][317] = 9'b111111111;
assign micromatrizz[49][318] = 9'b111111111;
assign micromatrizz[49][319] = 9'b111111111;
assign micromatrizz[49][320] = 9'b111111111;
assign micromatrizz[49][321] = 9'b111111111;
assign micromatrizz[49][322] = 9'b111111111;
assign micromatrizz[49][323] = 9'b111111111;
assign micromatrizz[49][324] = 9'b111111111;
assign micromatrizz[49][325] = 9'b111111111;
assign micromatrizz[49][326] = 9'b111111111;
assign micromatrizz[49][327] = 9'b111111111;
assign micromatrizz[49][328] = 9'b111111111;
assign micromatrizz[49][329] = 9'b111111111;
assign micromatrizz[49][330] = 9'b111111111;
assign micromatrizz[49][331] = 9'b111111111;
assign micromatrizz[49][332] = 9'b111111111;
assign micromatrizz[49][333] = 9'b111111111;
assign micromatrizz[49][334] = 9'b111111111;
assign micromatrizz[49][335] = 9'b111111111;
assign micromatrizz[49][336] = 9'b111111111;
assign micromatrizz[49][337] = 9'b111111111;
assign micromatrizz[49][338] = 9'b111111111;
assign micromatrizz[49][339] = 9'b111111111;
assign micromatrizz[49][340] = 9'b111111111;
assign micromatrizz[49][341] = 9'b111111111;
assign micromatrizz[49][342] = 9'b111111111;
assign micromatrizz[49][343] = 9'b111111111;
assign micromatrizz[49][344] = 9'b111111111;
assign micromatrizz[49][345] = 9'b111111111;
assign micromatrizz[49][346] = 9'b111111111;
assign micromatrizz[49][347] = 9'b111111111;
assign micromatrizz[49][348] = 9'b111111111;
assign micromatrizz[49][349] = 9'b111111111;
assign micromatrizz[49][350] = 9'b111111111;
assign micromatrizz[49][351] = 9'b111111111;
assign micromatrizz[49][352] = 9'b111111111;
assign micromatrizz[49][353] = 9'b111111111;
assign micromatrizz[49][354] = 9'b111111111;
assign micromatrizz[49][355] = 9'b111111111;
assign micromatrizz[49][356] = 9'b111111111;
assign micromatrizz[49][357] = 9'b111111111;
assign micromatrizz[49][358] = 9'b111111111;
assign micromatrizz[49][359] = 9'b111111111;
assign micromatrizz[49][360] = 9'b111110111;
assign micromatrizz[49][361] = 9'b111110010;
assign micromatrizz[49][362] = 9'b111110010;
assign micromatrizz[49][363] = 9'b111110010;
assign micromatrizz[49][364] = 9'b111110010;
assign micromatrizz[49][365] = 9'b111110010;
assign micromatrizz[49][366] = 9'b111111111;
assign micromatrizz[49][367] = 9'b111111111;
assign micromatrizz[49][368] = 9'b111111111;
assign micromatrizz[49][369] = 9'b111111111;
assign micromatrizz[49][370] = 9'b111111111;
assign micromatrizz[49][371] = 9'b111111111;
assign micromatrizz[49][372] = 9'b111111111;
assign micromatrizz[49][373] = 9'b111111111;
assign micromatrizz[49][374] = 9'b111111111;
assign micromatrizz[49][375] = 9'b111111111;
assign micromatrizz[49][376] = 9'b111111111;
assign micromatrizz[49][377] = 9'b111111111;
assign micromatrizz[49][378] = 9'b111111111;
assign micromatrizz[49][379] = 9'b111111111;
assign micromatrizz[49][380] = 9'b111111111;
assign micromatrizz[49][381] = 9'b111111111;
assign micromatrizz[49][382] = 9'b111111111;
assign micromatrizz[49][383] = 9'b111111111;
assign micromatrizz[49][384] = 9'b111111111;
assign micromatrizz[49][385] = 9'b111111111;
assign micromatrizz[49][386] = 9'b111111111;
assign micromatrizz[49][387] = 9'b111111111;
assign micromatrizz[49][388] = 9'b111111111;
assign micromatrizz[49][389] = 9'b111111111;
assign micromatrizz[49][390] = 9'b111111111;
assign micromatrizz[49][391] = 9'b111111111;
assign micromatrizz[49][392] = 9'b111111111;
assign micromatrizz[49][393] = 9'b111111111;
assign micromatrizz[49][394] = 9'b111111111;
assign micromatrizz[49][395] = 9'b111111111;
assign micromatrizz[49][396] = 9'b111111111;
assign micromatrizz[49][397] = 9'b111111111;
assign micromatrizz[49][398] = 9'b111111111;
assign micromatrizz[49][399] = 9'b111111111;
assign micromatrizz[49][400] = 9'b111111111;
assign micromatrizz[49][401] = 9'b111111111;
assign micromatrizz[49][402] = 9'b111111111;
assign micromatrizz[49][403] = 9'b111111111;
assign micromatrizz[49][404] = 9'b111111111;
assign micromatrizz[49][405] = 9'b111111111;
assign micromatrizz[49][406] = 9'b111111111;
assign micromatrizz[49][407] = 9'b111111111;
assign micromatrizz[49][408] = 9'b111111111;
assign micromatrizz[49][409] = 9'b111111111;
assign micromatrizz[49][410] = 9'b111111111;
assign micromatrizz[49][411] = 9'b111111111;
assign micromatrizz[49][412] = 9'b111111111;
assign micromatrizz[49][413] = 9'b111111111;
assign micromatrizz[49][414] = 9'b111111111;
assign micromatrizz[49][415] = 9'b111111111;
assign micromatrizz[49][416] = 9'b111111111;
assign micromatrizz[49][417] = 9'b111111111;
assign micromatrizz[49][418] = 9'b111111111;
assign micromatrizz[49][419] = 9'b111111111;
assign micromatrizz[49][420] = 9'b111111111;
assign micromatrizz[49][421] = 9'b111111111;
assign micromatrizz[49][422] = 9'b111111111;
assign micromatrizz[49][423] = 9'b111111111;
assign micromatrizz[49][424] = 9'b111111111;
assign micromatrizz[49][425] = 9'b111111111;
assign micromatrizz[49][426] = 9'b111111111;
assign micromatrizz[49][427] = 9'b111111111;
assign micromatrizz[49][428] = 9'b111111111;
assign micromatrizz[49][429] = 9'b111111111;
assign micromatrizz[49][430] = 9'b111111111;
assign micromatrizz[49][431] = 9'b111111111;
assign micromatrizz[49][432] = 9'b111111111;
assign micromatrizz[49][433] = 9'b111111111;
assign micromatrizz[49][434] = 9'b111111111;
assign micromatrizz[49][435] = 9'b111111111;
assign micromatrizz[49][436] = 9'b111111111;
assign micromatrizz[49][437] = 9'b111111111;
assign micromatrizz[49][438] = 9'b111111111;
assign micromatrizz[49][439] = 9'b111111111;
assign micromatrizz[49][440] = 9'b111111111;
assign micromatrizz[49][441] = 9'b111111111;
assign micromatrizz[49][442] = 9'b111111111;
assign micromatrizz[49][443] = 9'b111111111;
assign micromatrizz[49][444] = 9'b111111111;
assign micromatrizz[49][445] = 9'b111111111;
assign micromatrizz[49][446] = 9'b111111111;
assign micromatrizz[49][447] = 9'b111111111;
assign micromatrizz[49][448] = 9'b111111111;
assign micromatrizz[49][449] = 9'b111111111;
assign micromatrizz[49][450] = 9'b111111111;
assign micromatrizz[49][451] = 9'b111111111;
assign micromatrizz[49][452] = 9'b111111111;
assign micromatrizz[49][453] = 9'b111111111;
assign micromatrizz[49][454] = 9'b111111111;
assign micromatrizz[49][455] = 9'b111111111;
assign micromatrizz[49][456] = 9'b111111111;
assign micromatrizz[49][457] = 9'b111111111;
assign micromatrizz[49][458] = 9'b111111111;
assign micromatrizz[49][459] = 9'b111111111;
assign micromatrizz[49][460] = 9'b111111111;
assign micromatrizz[49][461] = 9'b111111111;
assign micromatrizz[49][462] = 9'b111111111;
assign micromatrizz[49][463] = 9'b111111111;
assign micromatrizz[49][464] = 9'b111111111;
assign micromatrizz[49][465] = 9'b111111111;
assign micromatrizz[49][466] = 9'b111111111;
assign micromatrizz[49][467] = 9'b111111111;
assign micromatrizz[49][468] = 9'b111111111;
assign micromatrizz[49][469] = 9'b111111111;
assign micromatrizz[49][470] = 9'b111111111;
assign micromatrizz[49][471] = 9'b111111111;
assign micromatrizz[49][472] = 9'b111111111;
assign micromatrizz[49][473] = 9'b111111111;
assign micromatrizz[49][474] = 9'b111111111;
assign micromatrizz[49][475] = 9'b111111111;
assign micromatrizz[49][476] = 9'b111111111;
assign micromatrizz[49][477] = 9'b111111111;
assign micromatrizz[49][478] = 9'b111111111;
assign micromatrizz[49][479] = 9'b111111111;
assign micromatrizz[49][480] = 9'b111111111;
assign micromatrizz[49][481] = 9'b111111111;
assign micromatrizz[49][482] = 9'b111111111;
assign micromatrizz[49][483] = 9'b111111111;
assign micromatrizz[49][484] = 9'b111111111;
assign micromatrizz[49][485] = 9'b111111111;
assign micromatrizz[49][486] = 9'b111111111;
assign micromatrizz[49][487] = 9'b111111111;
assign micromatrizz[49][488] = 9'b111111111;
assign micromatrizz[49][489] = 9'b111111111;
assign micromatrizz[49][490] = 9'b111111111;
assign micromatrizz[49][491] = 9'b111111111;
assign micromatrizz[49][492] = 9'b111111111;
assign micromatrizz[49][493] = 9'b111111111;
assign micromatrizz[49][494] = 9'b111111111;
assign micromatrizz[49][495] = 9'b111111111;
assign micromatrizz[49][496] = 9'b111111111;
assign micromatrizz[49][497] = 9'b111111111;
assign micromatrizz[49][498] = 9'b111111111;
assign micromatrizz[49][499] = 9'b111111111;
assign micromatrizz[49][500] = 9'b111111111;
assign micromatrizz[49][501] = 9'b111111111;
assign micromatrizz[49][502] = 9'b111111111;
assign micromatrizz[49][503] = 9'b111111111;
assign micromatrizz[49][504] = 9'b111111111;
assign micromatrizz[49][505] = 9'b111111111;
assign micromatrizz[49][506] = 9'b111111111;
assign micromatrizz[49][507] = 9'b111111111;
assign micromatrizz[49][508] = 9'b111111111;
assign micromatrizz[49][509] = 9'b111111111;
assign micromatrizz[49][510] = 9'b111111111;
assign micromatrizz[49][511] = 9'b111111111;
assign micromatrizz[49][512] = 9'b111111111;
assign micromatrizz[49][513] = 9'b111111111;
assign micromatrizz[49][514] = 9'b111111111;
assign micromatrizz[49][515] = 9'b111111111;
assign micromatrizz[49][516] = 9'b111110010;
assign micromatrizz[49][517] = 9'b111110010;
assign micromatrizz[49][518] = 9'b111110011;
assign micromatrizz[49][519] = 9'b111110011;
assign micromatrizz[49][520] = 9'b111110010;
assign micromatrizz[49][521] = 9'b111110010;
assign micromatrizz[49][522] = 9'b111110011;
assign micromatrizz[49][523] = 9'b111110111;
assign micromatrizz[49][524] = 9'b111111111;
assign micromatrizz[49][525] = 9'b111111111;
assign micromatrizz[49][526] = 9'b111111111;
assign micromatrizz[49][527] = 9'b111111111;
assign micromatrizz[49][528] = 9'b111111111;
assign micromatrizz[49][529] = 9'b111111111;
assign micromatrizz[49][530] = 9'b111111111;
assign micromatrizz[49][531] = 9'b111111111;
assign micromatrizz[49][532] = 9'b111111111;
assign micromatrizz[49][533] = 9'b111111111;
assign micromatrizz[49][534] = 9'b111111111;
assign micromatrizz[49][535] = 9'b111111111;
assign micromatrizz[49][536] = 9'b111111111;
assign micromatrizz[49][537] = 9'b111111111;
assign micromatrizz[49][538] = 9'b111111111;
assign micromatrizz[49][539] = 9'b111111111;
assign micromatrizz[49][540] = 9'b111111111;
assign micromatrizz[49][541] = 9'b111111111;
assign micromatrizz[49][542] = 9'b111111111;
assign micromatrizz[49][543] = 9'b111111111;
assign micromatrizz[49][544] = 9'b111111111;
assign micromatrizz[49][545] = 9'b111111111;
assign micromatrizz[49][546] = 9'b111111111;
assign micromatrizz[49][547] = 9'b111111111;
assign micromatrizz[49][548] = 9'b111111111;
assign micromatrizz[49][549] = 9'b111111111;
assign micromatrizz[49][550] = 9'b111111111;
assign micromatrizz[49][551] = 9'b111111111;
assign micromatrizz[49][552] = 9'b111111111;
assign micromatrizz[49][553] = 9'b111111111;
assign micromatrizz[49][554] = 9'b111111111;
assign micromatrizz[49][555] = 9'b111111111;
assign micromatrizz[49][556] = 9'b111111111;
assign micromatrizz[49][557] = 9'b111111111;
assign micromatrizz[49][558] = 9'b111110010;
assign micromatrizz[49][559] = 9'b111110010;
assign micromatrizz[49][560] = 9'b111110011;
assign micromatrizz[49][561] = 9'b111110011;
assign micromatrizz[49][562] = 9'b111110011;
assign micromatrizz[49][563] = 9'b111110011;
assign micromatrizz[49][564] = 9'b111110011;
assign micromatrizz[49][565] = 9'b111111111;
assign micromatrizz[49][566] = 9'b111111111;
assign micromatrizz[49][567] = 9'b111111111;
assign micromatrizz[49][568] = 9'b111111111;
assign micromatrizz[49][569] = 9'b111111111;
assign micromatrizz[49][570] = 9'b111111111;
assign micromatrizz[49][571] = 9'b111111111;
assign micromatrizz[49][572] = 9'b111111111;
assign micromatrizz[49][573] = 9'b111111111;
assign micromatrizz[49][574] = 9'b111111111;
assign micromatrizz[49][575] = 9'b111111111;
assign micromatrizz[49][576] = 9'b111111111;
assign micromatrizz[49][577] = 9'b111111111;
assign micromatrizz[49][578] = 9'b111111111;
assign micromatrizz[49][579] = 9'b111111111;
assign micromatrizz[49][580] = 9'b111111111;
assign micromatrizz[49][581] = 9'b111110010;
assign micromatrizz[49][582] = 9'b111110011;
assign micromatrizz[49][583] = 9'b111110011;
assign micromatrizz[49][584] = 9'b111110010;
assign micromatrizz[49][585] = 9'b111110010;
assign micromatrizz[49][586] = 9'b111110011;
assign micromatrizz[49][587] = 9'b111110011;
assign micromatrizz[49][588] = 9'b111111111;
assign micromatrizz[49][589] = 9'b111111111;
assign micromatrizz[49][590] = 9'b111111111;
assign micromatrizz[49][591] = 9'b111111111;
assign micromatrizz[49][592] = 9'b111111111;
assign micromatrizz[49][593] = 9'b111111111;
assign micromatrizz[49][594] = 9'b111111111;
assign micromatrizz[49][595] = 9'b111111111;
assign micromatrizz[49][596] = 9'b111111111;
assign micromatrizz[49][597] = 9'b111111111;
assign micromatrizz[49][598] = 9'b111111111;
assign micromatrizz[49][599] = 9'b111111111;
assign micromatrizz[49][600] = 9'b111111111;
assign micromatrizz[49][601] = 9'b111111111;
assign micromatrizz[49][602] = 9'b111111111;
assign micromatrizz[49][603] = 9'b111111111;
assign micromatrizz[49][604] = 9'b111111111;
assign micromatrizz[49][605] = 9'b111111111;
assign micromatrizz[49][606] = 9'b111111111;
assign micromatrizz[49][607] = 9'b111111111;
assign micromatrizz[49][608] = 9'b111111111;
assign micromatrizz[49][609] = 9'b111111111;
assign micromatrizz[49][610] = 9'b111111111;
assign micromatrizz[49][611] = 9'b111111111;
assign micromatrizz[49][612] = 9'b111111111;
assign micromatrizz[49][613] = 9'b111111111;
assign micromatrizz[49][614] = 9'b111111111;
assign micromatrizz[49][615] = 9'b111111111;
assign micromatrizz[49][616] = 9'b111111111;
assign micromatrizz[49][617] = 9'b111111111;
assign micromatrizz[49][618] = 9'b111111111;
assign micromatrizz[49][619] = 9'b111111111;
assign micromatrizz[49][620] = 9'b111111111;
assign micromatrizz[49][621] = 9'b111111111;
assign micromatrizz[49][622] = 9'b111111111;
assign micromatrizz[49][623] = 9'b111111111;
assign micromatrizz[49][624] = 9'b111111111;
assign micromatrizz[49][625] = 9'b111111111;
assign micromatrizz[49][626] = 9'b111111111;
assign micromatrizz[49][627] = 9'b111111111;
assign micromatrizz[49][628] = 9'b111111111;
assign micromatrizz[49][629] = 9'b111111111;
assign micromatrizz[49][630] = 9'b111111111;
assign micromatrizz[49][631] = 9'b111111111;
assign micromatrizz[49][632] = 9'b111111111;
assign micromatrizz[49][633] = 9'b111111111;
assign micromatrizz[49][634] = 9'b111111111;
assign micromatrizz[49][635] = 9'b111111111;
assign micromatrizz[49][636] = 9'b111111111;
assign micromatrizz[49][637] = 9'b111111111;
assign micromatrizz[49][638] = 9'b111111111;
assign micromatrizz[49][639] = 9'b111111111;
assign micromatrizz[50][0] = 9'b111111111;
assign micromatrizz[50][1] = 9'b111111111;
assign micromatrizz[50][2] = 9'b111111111;
assign micromatrizz[50][3] = 9'b111111111;
assign micromatrizz[50][4] = 9'b111111111;
assign micromatrizz[50][5] = 9'b111111111;
assign micromatrizz[50][6] = 9'b111111111;
assign micromatrizz[50][7] = 9'b111111111;
assign micromatrizz[50][8] = 9'b111111111;
assign micromatrizz[50][9] = 9'b111111111;
assign micromatrizz[50][10] = 9'b111111111;
assign micromatrizz[50][11] = 9'b111111111;
assign micromatrizz[50][12] = 9'b111111111;
assign micromatrizz[50][13] = 9'b111111111;
assign micromatrizz[50][14] = 9'b111111111;
assign micromatrizz[50][15] = 9'b111111111;
assign micromatrizz[50][16] = 9'b111111111;
assign micromatrizz[50][17] = 9'b111111111;
assign micromatrizz[50][18] = 9'b111111111;
assign micromatrizz[50][19] = 9'b111111111;
assign micromatrizz[50][20] = 9'b111111111;
assign micromatrizz[50][21] = 9'b111111111;
assign micromatrizz[50][22] = 9'b111111111;
assign micromatrizz[50][23] = 9'b111111111;
assign micromatrizz[50][24] = 9'b111111111;
assign micromatrizz[50][25] = 9'b111111111;
assign micromatrizz[50][26] = 9'b111111111;
assign micromatrizz[50][27] = 9'b111111111;
assign micromatrizz[50][28] = 9'b111111111;
assign micromatrizz[50][29] = 9'b111111111;
assign micromatrizz[50][30] = 9'b111111111;
assign micromatrizz[50][31] = 9'b111111111;
assign micromatrizz[50][32] = 9'b111111111;
assign micromatrizz[50][33] = 9'b111111111;
assign micromatrizz[50][34] = 9'b111111111;
assign micromatrizz[50][35] = 9'b111111111;
assign micromatrizz[50][36] = 9'b111111111;
assign micromatrizz[50][37] = 9'b111111111;
assign micromatrizz[50][38] = 9'b111111111;
assign micromatrizz[50][39] = 9'b111111111;
assign micromatrizz[50][40] = 9'b111111111;
assign micromatrizz[50][41] = 9'b111111111;
assign micromatrizz[50][42] = 9'b111111111;
assign micromatrizz[50][43] = 9'b111111111;
assign micromatrizz[50][44] = 9'b111111111;
assign micromatrizz[50][45] = 9'b111111111;
assign micromatrizz[50][46] = 9'b111111111;
assign micromatrizz[50][47] = 9'b111111111;
assign micromatrizz[50][48] = 9'b111111111;
assign micromatrizz[50][49] = 9'b111111111;
assign micromatrizz[50][50] = 9'b111111111;
assign micromatrizz[50][51] = 9'b111111111;
assign micromatrizz[50][52] = 9'b111111111;
assign micromatrizz[50][53] = 9'b111111111;
assign micromatrizz[50][54] = 9'b111111111;
assign micromatrizz[50][55] = 9'b111111111;
assign micromatrizz[50][56] = 9'b111111111;
assign micromatrizz[50][57] = 9'b111111111;
assign micromatrizz[50][58] = 9'b111111111;
assign micromatrizz[50][59] = 9'b111111111;
assign micromatrizz[50][60] = 9'b111111111;
assign micromatrizz[50][61] = 9'b111111111;
assign micromatrizz[50][62] = 9'b111111111;
assign micromatrizz[50][63] = 9'b111111111;
assign micromatrizz[50][64] = 9'b111111111;
assign micromatrizz[50][65] = 9'b111111111;
assign micromatrizz[50][66] = 9'b111111111;
assign micromatrizz[50][67] = 9'b111111111;
assign micromatrizz[50][68] = 9'b111111111;
assign micromatrizz[50][69] = 9'b111111111;
assign micromatrizz[50][70] = 9'b111111111;
assign micromatrizz[50][71] = 9'b111111111;
assign micromatrizz[50][72] = 9'b111111111;
assign micromatrizz[50][73] = 9'b111111111;
assign micromatrizz[50][74] = 9'b111111111;
assign micromatrizz[50][75] = 9'b111111111;
assign micromatrizz[50][76] = 9'b111111111;
assign micromatrizz[50][77] = 9'b111111111;
assign micromatrizz[50][78] = 9'b111111111;
assign micromatrizz[50][79] = 9'b111111111;
assign micromatrizz[50][80] = 9'b111111111;
assign micromatrizz[50][81] = 9'b111111111;
assign micromatrizz[50][82] = 9'b111111111;
assign micromatrizz[50][83] = 9'b111111111;
assign micromatrizz[50][84] = 9'b111111111;
assign micromatrizz[50][85] = 9'b111111111;
assign micromatrizz[50][86] = 9'b111111111;
assign micromatrizz[50][87] = 9'b111111111;
assign micromatrizz[50][88] = 9'b111111111;
assign micromatrizz[50][89] = 9'b111111111;
assign micromatrizz[50][90] = 9'b111111111;
assign micromatrizz[50][91] = 9'b111111111;
assign micromatrizz[50][92] = 9'b111111111;
assign micromatrizz[50][93] = 9'b111111111;
assign micromatrizz[50][94] = 9'b111111111;
assign micromatrizz[50][95] = 9'b111111111;
assign micromatrizz[50][96] = 9'b111111111;
assign micromatrizz[50][97] = 9'b111111111;
assign micromatrizz[50][98] = 9'b111111111;
assign micromatrizz[50][99] = 9'b111111111;
assign micromatrizz[50][100] = 9'b111111111;
assign micromatrizz[50][101] = 9'b111111111;
assign micromatrizz[50][102] = 9'b111111111;
assign micromatrizz[50][103] = 9'b111111111;
assign micromatrizz[50][104] = 9'b111111111;
assign micromatrizz[50][105] = 9'b111111111;
assign micromatrizz[50][106] = 9'b111111111;
assign micromatrizz[50][107] = 9'b111111111;
assign micromatrizz[50][108] = 9'b111111111;
assign micromatrizz[50][109] = 9'b111111111;
assign micromatrizz[50][110] = 9'b111111111;
assign micromatrizz[50][111] = 9'b111111111;
assign micromatrizz[50][112] = 9'b111111111;
assign micromatrizz[50][113] = 9'b111111111;
assign micromatrizz[50][114] = 9'b111111111;
assign micromatrizz[50][115] = 9'b111111111;
assign micromatrizz[50][116] = 9'b111111111;
assign micromatrizz[50][117] = 9'b111111111;
assign micromatrizz[50][118] = 9'b111111111;
assign micromatrizz[50][119] = 9'b111111111;
assign micromatrizz[50][120] = 9'b111111111;
assign micromatrizz[50][121] = 9'b111111111;
assign micromatrizz[50][122] = 9'b111111111;
assign micromatrizz[50][123] = 9'b111111111;
assign micromatrizz[50][124] = 9'b111111111;
assign micromatrizz[50][125] = 9'b111111111;
assign micromatrizz[50][126] = 9'b111111111;
assign micromatrizz[50][127] = 9'b111111111;
assign micromatrizz[50][128] = 9'b111111111;
assign micromatrizz[50][129] = 9'b111111111;
assign micromatrizz[50][130] = 9'b111111111;
assign micromatrizz[50][131] = 9'b111111111;
assign micromatrizz[50][132] = 9'b111111111;
assign micromatrizz[50][133] = 9'b111111111;
assign micromatrizz[50][134] = 9'b111111111;
assign micromatrizz[50][135] = 9'b111111111;
assign micromatrizz[50][136] = 9'b111111111;
assign micromatrizz[50][137] = 9'b111111111;
assign micromatrizz[50][138] = 9'b111111111;
assign micromatrizz[50][139] = 9'b111111111;
assign micromatrizz[50][140] = 9'b111111111;
assign micromatrizz[50][141] = 9'b111111111;
assign micromatrizz[50][142] = 9'b111111111;
assign micromatrizz[50][143] = 9'b111111111;
assign micromatrizz[50][144] = 9'b111111111;
assign micromatrizz[50][145] = 9'b111111111;
assign micromatrizz[50][146] = 9'b111111111;
assign micromatrizz[50][147] = 9'b111111111;
assign micromatrizz[50][148] = 9'b111111111;
assign micromatrizz[50][149] = 9'b111111111;
assign micromatrizz[50][150] = 9'b111111111;
assign micromatrizz[50][151] = 9'b111111111;
assign micromatrizz[50][152] = 9'b111111111;
assign micromatrizz[50][153] = 9'b111111111;
assign micromatrizz[50][154] = 9'b111111111;
assign micromatrizz[50][155] = 9'b111111111;
assign micromatrizz[50][156] = 9'b111111111;
assign micromatrizz[50][157] = 9'b111111111;
assign micromatrizz[50][158] = 9'b111111111;
assign micromatrizz[50][159] = 9'b111111111;
assign micromatrizz[50][160] = 9'b111111111;
assign micromatrizz[50][161] = 9'b111111111;
assign micromatrizz[50][162] = 9'b111111111;
assign micromatrizz[50][163] = 9'b111111111;
assign micromatrizz[50][164] = 9'b111111111;
assign micromatrizz[50][165] = 9'b111111111;
assign micromatrizz[50][166] = 9'b111111111;
assign micromatrizz[50][167] = 9'b111111111;
assign micromatrizz[50][168] = 9'b111111111;
assign micromatrizz[50][169] = 9'b111111111;
assign micromatrizz[50][170] = 9'b111111111;
assign micromatrizz[50][171] = 9'b111111111;
assign micromatrizz[50][172] = 9'b111111111;
assign micromatrizz[50][173] = 9'b111111111;
assign micromatrizz[50][174] = 9'b111111111;
assign micromatrizz[50][175] = 9'b111111111;
assign micromatrizz[50][176] = 9'b111111111;
assign micromatrizz[50][177] = 9'b111111111;
assign micromatrizz[50][178] = 9'b111111111;
assign micromatrizz[50][179] = 9'b111111111;
assign micromatrizz[50][180] = 9'b111111111;
assign micromatrizz[50][181] = 9'b111111111;
assign micromatrizz[50][182] = 9'b111111111;
assign micromatrizz[50][183] = 9'b111111111;
assign micromatrizz[50][184] = 9'b111111111;
assign micromatrizz[50][185] = 9'b111111111;
assign micromatrizz[50][186] = 9'b111111111;
assign micromatrizz[50][187] = 9'b111111111;
assign micromatrizz[50][188] = 9'b111111111;
assign micromatrizz[50][189] = 9'b111111111;
assign micromatrizz[50][190] = 9'b111111111;
assign micromatrizz[50][191] = 9'b111111111;
assign micromatrizz[50][192] = 9'b111111111;
assign micromatrizz[50][193] = 9'b111111111;
assign micromatrizz[50][194] = 9'b111111111;
assign micromatrizz[50][195] = 9'b111110010;
assign micromatrizz[50][196] = 9'b111110010;
assign micromatrizz[50][197] = 9'b111110011;
assign micromatrizz[50][198] = 9'b111110011;
assign micromatrizz[50][199] = 9'b111110010;
assign micromatrizz[50][200] = 9'b111110010;
assign micromatrizz[50][201] = 9'b111110011;
assign micromatrizz[50][202] = 9'b111110111;
assign micromatrizz[50][203] = 9'b111111111;
assign micromatrizz[50][204] = 9'b111111111;
assign micromatrizz[50][205] = 9'b111111111;
assign micromatrizz[50][206] = 9'b111111111;
assign micromatrizz[50][207] = 9'b111111111;
assign micromatrizz[50][208] = 9'b111111111;
assign micromatrizz[50][209] = 9'b111111111;
assign micromatrizz[50][210] = 9'b111111111;
assign micromatrizz[50][211] = 9'b111111111;
assign micromatrizz[50][212] = 9'b111111111;
assign micromatrizz[50][213] = 9'b111111111;
assign micromatrizz[50][214] = 9'b111111111;
assign micromatrizz[50][215] = 9'b111111111;
assign micromatrizz[50][216] = 9'b111111111;
assign micromatrizz[50][217] = 9'b111111111;
assign micromatrizz[50][218] = 9'b111111111;
assign micromatrizz[50][219] = 9'b111111111;
assign micromatrizz[50][220] = 9'b111111111;
assign micromatrizz[50][221] = 9'b111111111;
assign micromatrizz[50][222] = 9'b111111111;
assign micromatrizz[50][223] = 9'b111111111;
assign micromatrizz[50][224] = 9'b111111111;
assign micromatrizz[50][225] = 9'b111111111;
assign micromatrizz[50][226] = 9'b111111111;
assign micromatrizz[50][227] = 9'b111111111;
assign micromatrizz[50][228] = 9'b111111111;
assign micromatrizz[50][229] = 9'b111111111;
assign micromatrizz[50][230] = 9'b111111111;
assign micromatrizz[50][231] = 9'b111111111;
assign micromatrizz[50][232] = 9'b111111111;
assign micromatrizz[50][233] = 9'b111111111;
assign micromatrizz[50][234] = 9'b111111111;
assign micromatrizz[50][235] = 9'b111111111;
assign micromatrizz[50][236] = 9'b111111111;
assign micromatrizz[50][237] = 9'b111111111;
assign micromatrizz[50][238] = 9'b111111111;
assign micromatrizz[50][239] = 9'b111111111;
assign micromatrizz[50][240] = 9'b111111111;
assign micromatrizz[50][241] = 9'b111111111;
assign micromatrizz[50][242] = 9'b111111111;
assign micromatrizz[50][243] = 9'b111111111;
assign micromatrizz[50][244] = 9'b111111111;
assign micromatrizz[50][245] = 9'b111111111;
assign micromatrizz[50][246] = 9'b111111111;
assign micromatrizz[50][247] = 9'b111111111;
assign micromatrizz[50][248] = 9'b111111111;
assign micromatrizz[50][249] = 9'b111111111;
assign micromatrizz[50][250] = 9'b111111111;
assign micromatrizz[50][251] = 9'b111111111;
assign micromatrizz[50][252] = 9'b111111111;
assign micromatrizz[50][253] = 9'b111111111;
assign micromatrizz[50][254] = 9'b111111111;
assign micromatrizz[50][255] = 9'b111111111;
assign micromatrizz[50][256] = 9'b111111111;
assign micromatrizz[50][257] = 9'b111111111;
assign micromatrizz[50][258] = 9'b111111111;
assign micromatrizz[50][259] = 9'b111111111;
assign micromatrizz[50][260] = 9'b111111111;
assign micromatrizz[50][261] = 9'b111111111;
assign micromatrizz[50][262] = 9'b111111111;
assign micromatrizz[50][263] = 9'b111111111;
assign micromatrizz[50][264] = 9'b111111111;
assign micromatrizz[50][265] = 9'b111111111;
assign micromatrizz[50][266] = 9'b111111111;
assign micromatrizz[50][267] = 9'b111111111;
assign micromatrizz[50][268] = 9'b111111111;
assign micromatrizz[50][269] = 9'b111111111;
assign micromatrizz[50][270] = 9'b111111111;
assign micromatrizz[50][271] = 9'b111111111;
assign micromatrizz[50][272] = 9'b111111111;
assign micromatrizz[50][273] = 9'b111111111;
assign micromatrizz[50][274] = 9'b111111111;
assign micromatrizz[50][275] = 9'b111111111;
assign micromatrizz[50][276] = 9'b111111111;
assign micromatrizz[50][277] = 9'b111111111;
assign micromatrizz[50][278] = 9'b111111111;
assign micromatrizz[50][279] = 9'b111111111;
assign micromatrizz[50][280] = 9'b111111111;
assign micromatrizz[50][281] = 9'b111111111;
assign micromatrizz[50][282] = 9'b111111111;
assign micromatrizz[50][283] = 9'b111111111;
assign micromatrizz[50][284] = 9'b111111111;
assign micromatrizz[50][285] = 9'b111111111;
assign micromatrizz[50][286] = 9'b111111111;
assign micromatrizz[50][287] = 9'b111111111;
assign micromatrizz[50][288] = 9'b111111111;
assign micromatrizz[50][289] = 9'b111111111;
assign micromatrizz[50][290] = 9'b111111111;
assign micromatrizz[50][291] = 9'b111111111;
assign micromatrizz[50][292] = 9'b111111111;
assign micromatrizz[50][293] = 9'b111111111;
assign micromatrizz[50][294] = 9'b111111111;
assign micromatrizz[50][295] = 9'b111111111;
assign micromatrizz[50][296] = 9'b111111111;
assign micromatrizz[50][297] = 9'b111111111;
assign micromatrizz[50][298] = 9'b111111111;
assign micromatrizz[50][299] = 9'b111111111;
assign micromatrizz[50][300] = 9'b111111111;
assign micromatrizz[50][301] = 9'b111111111;
assign micromatrizz[50][302] = 9'b111111111;
assign micromatrizz[50][303] = 9'b111111111;
assign micromatrizz[50][304] = 9'b111111111;
assign micromatrizz[50][305] = 9'b111111111;
assign micromatrizz[50][306] = 9'b111111111;
assign micromatrizz[50][307] = 9'b111111111;
assign micromatrizz[50][308] = 9'b111111111;
assign micromatrizz[50][309] = 9'b111111111;
assign micromatrizz[50][310] = 9'b111111111;
assign micromatrizz[50][311] = 9'b111111111;
assign micromatrizz[50][312] = 9'b111111111;
assign micromatrizz[50][313] = 9'b111111111;
assign micromatrizz[50][314] = 9'b111111111;
assign micromatrizz[50][315] = 9'b111111111;
assign micromatrizz[50][316] = 9'b111111111;
assign micromatrizz[50][317] = 9'b111111111;
assign micromatrizz[50][318] = 9'b111111111;
assign micromatrizz[50][319] = 9'b111111111;
assign micromatrizz[50][320] = 9'b111111111;
assign micromatrizz[50][321] = 9'b111111111;
assign micromatrizz[50][322] = 9'b111111111;
assign micromatrizz[50][323] = 9'b111111111;
assign micromatrizz[50][324] = 9'b111111111;
assign micromatrizz[50][325] = 9'b111111111;
assign micromatrizz[50][326] = 9'b111111111;
assign micromatrizz[50][327] = 9'b111111111;
assign micromatrizz[50][328] = 9'b111111111;
assign micromatrizz[50][329] = 9'b111111111;
assign micromatrizz[50][330] = 9'b111111111;
assign micromatrizz[50][331] = 9'b111111111;
assign micromatrizz[50][332] = 9'b111111111;
assign micromatrizz[50][333] = 9'b111111111;
assign micromatrizz[50][334] = 9'b111111111;
assign micromatrizz[50][335] = 9'b111111111;
assign micromatrizz[50][336] = 9'b111111111;
assign micromatrizz[50][337] = 9'b111111111;
assign micromatrizz[50][338] = 9'b111111111;
assign micromatrizz[50][339] = 9'b111111111;
assign micromatrizz[50][340] = 9'b111111111;
assign micromatrizz[50][341] = 9'b111111111;
assign micromatrizz[50][342] = 9'b111111111;
assign micromatrizz[50][343] = 9'b111111111;
assign micromatrizz[50][344] = 9'b111111111;
assign micromatrizz[50][345] = 9'b111111111;
assign micromatrizz[50][346] = 9'b111111111;
assign micromatrizz[50][347] = 9'b111111111;
assign micromatrizz[50][348] = 9'b111111111;
assign micromatrizz[50][349] = 9'b111111111;
assign micromatrizz[50][350] = 9'b111111111;
assign micromatrizz[50][351] = 9'b111111111;
assign micromatrizz[50][352] = 9'b111111111;
assign micromatrizz[50][353] = 9'b111111111;
assign micromatrizz[50][354] = 9'b111111111;
assign micromatrizz[50][355] = 9'b111111111;
assign micromatrizz[50][356] = 9'b111111111;
assign micromatrizz[50][357] = 9'b111111111;
assign micromatrizz[50][358] = 9'b111111111;
assign micromatrizz[50][359] = 9'b111110010;
assign micromatrizz[50][360] = 9'b111110010;
assign micromatrizz[50][361] = 9'b111110010;
assign micromatrizz[50][362] = 9'b111110010;
assign micromatrizz[50][363] = 9'b111110011;
assign micromatrizz[50][364] = 9'b111110011;
assign micromatrizz[50][365] = 9'b111110010;
assign micromatrizz[50][366] = 9'b111111111;
assign micromatrizz[50][367] = 9'b111111111;
assign micromatrizz[50][368] = 9'b111111111;
assign micromatrizz[50][369] = 9'b111111111;
assign micromatrizz[50][370] = 9'b111111111;
assign micromatrizz[50][371] = 9'b111111111;
assign micromatrizz[50][372] = 9'b111111111;
assign micromatrizz[50][373] = 9'b111111111;
assign micromatrizz[50][374] = 9'b111111111;
assign micromatrizz[50][375] = 9'b111111111;
assign micromatrizz[50][376] = 9'b111111111;
assign micromatrizz[50][377] = 9'b111111111;
assign micromatrizz[50][378] = 9'b111111111;
assign micromatrizz[50][379] = 9'b111111111;
assign micromatrizz[50][380] = 9'b111111111;
assign micromatrizz[50][381] = 9'b111111111;
assign micromatrizz[50][382] = 9'b111111111;
assign micromatrizz[50][383] = 9'b111111111;
assign micromatrizz[50][384] = 9'b111111111;
assign micromatrizz[50][385] = 9'b111111111;
assign micromatrizz[50][386] = 9'b111111111;
assign micromatrizz[50][387] = 9'b111111111;
assign micromatrizz[50][388] = 9'b111111111;
assign micromatrizz[50][389] = 9'b111111111;
assign micromatrizz[50][390] = 9'b111111111;
assign micromatrizz[50][391] = 9'b111111111;
assign micromatrizz[50][392] = 9'b111111111;
assign micromatrizz[50][393] = 9'b111111111;
assign micromatrizz[50][394] = 9'b111111111;
assign micromatrizz[50][395] = 9'b111111111;
assign micromatrizz[50][396] = 9'b111111111;
assign micromatrizz[50][397] = 9'b111111111;
assign micromatrizz[50][398] = 9'b111111111;
assign micromatrizz[50][399] = 9'b111111111;
assign micromatrizz[50][400] = 9'b111111111;
assign micromatrizz[50][401] = 9'b111111111;
assign micromatrizz[50][402] = 9'b111111111;
assign micromatrizz[50][403] = 9'b111111111;
assign micromatrizz[50][404] = 9'b111111111;
assign micromatrizz[50][405] = 9'b111111111;
assign micromatrizz[50][406] = 9'b111111111;
assign micromatrizz[50][407] = 9'b111111111;
assign micromatrizz[50][408] = 9'b111111111;
assign micromatrizz[50][409] = 9'b111111111;
assign micromatrizz[50][410] = 9'b111111111;
assign micromatrizz[50][411] = 9'b111111111;
assign micromatrizz[50][412] = 9'b111111111;
assign micromatrizz[50][413] = 9'b111111111;
assign micromatrizz[50][414] = 9'b111111111;
assign micromatrizz[50][415] = 9'b111111111;
assign micromatrizz[50][416] = 9'b111111111;
assign micromatrizz[50][417] = 9'b111111111;
assign micromatrizz[50][418] = 9'b111111111;
assign micromatrizz[50][419] = 9'b111111111;
assign micromatrizz[50][420] = 9'b111111111;
assign micromatrizz[50][421] = 9'b111111111;
assign micromatrizz[50][422] = 9'b111111111;
assign micromatrizz[50][423] = 9'b111111111;
assign micromatrizz[50][424] = 9'b111111111;
assign micromatrizz[50][425] = 9'b111111111;
assign micromatrizz[50][426] = 9'b111111111;
assign micromatrizz[50][427] = 9'b111111111;
assign micromatrizz[50][428] = 9'b111111111;
assign micromatrizz[50][429] = 9'b111111111;
assign micromatrizz[50][430] = 9'b111111111;
assign micromatrizz[50][431] = 9'b111111111;
assign micromatrizz[50][432] = 9'b111111111;
assign micromatrizz[50][433] = 9'b111111111;
assign micromatrizz[50][434] = 9'b111111111;
assign micromatrizz[50][435] = 9'b111111111;
assign micromatrizz[50][436] = 9'b111111111;
assign micromatrizz[50][437] = 9'b111111111;
assign micromatrizz[50][438] = 9'b111111111;
assign micromatrizz[50][439] = 9'b111111111;
assign micromatrizz[50][440] = 9'b111111111;
assign micromatrizz[50][441] = 9'b111111111;
assign micromatrizz[50][442] = 9'b111111111;
assign micromatrizz[50][443] = 9'b111111111;
assign micromatrizz[50][444] = 9'b111111111;
assign micromatrizz[50][445] = 9'b111111111;
assign micromatrizz[50][446] = 9'b111111111;
assign micromatrizz[50][447] = 9'b111111111;
assign micromatrizz[50][448] = 9'b111111111;
assign micromatrizz[50][449] = 9'b111111111;
assign micromatrizz[50][450] = 9'b111111111;
assign micromatrizz[50][451] = 9'b111111111;
assign micromatrizz[50][452] = 9'b111111111;
assign micromatrizz[50][453] = 9'b111111111;
assign micromatrizz[50][454] = 9'b111111111;
assign micromatrizz[50][455] = 9'b111111111;
assign micromatrizz[50][456] = 9'b111111111;
assign micromatrizz[50][457] = 9'b111111111;
assign micromatrizz[50][458] = 9'b111111111;
assign micromatrizz[50][459] = 9'b111111111;
assign micromatrizz[50][460] = 9'b111111111;
assign micromatrizz[50][461] = 9'b111111111;
assign micromatrizz[50][462] = 9'b111111111;
assign micromatrizz[50][463] = 9'b111111111;
assign micromatrizz[50][464] = 9'b111111111;
assign micromatrizz[50][465] = 9'b111111111;
assign micromatrizz[50][466] = 9'b111111111;
assign micromatrizz[50][467] = 9'b111111111;
assign micromatrizz[50][468] = 9'b111111111;
assign micromatrizz[50][469] = 9'b111111111;
assign micromatrizz[50][470] = 9'b111111111;
assign micromatrizz[50][471] = 9'b111111111;
assign micromatrizz[50][472] = 9'b111111111;
assign micromatrizz[50][473] = 9'b111111111;
assign micromatrizz[50][474] = 9'b111111111;
assign micromatrizz[50][475] = 9'b111111111;
assign micromatrizz[50][476] = 9'b111111111;
assign micromatrizz[50][477] = 9'b111111111;
assign micromatrizz[50][478] = 9'b111111111;
assign micromatrizz[50][479] = 9'b111111111;
assign micromatrizz[50][480] = 9'b111111111;
assign micromatrizz[50][481] = 9'b111111111;
assign micromatrizz[50][482] = 9'b111111111;
assign micromatrizz[50][483] = 9'b111111111;
assign micromatrizz[50][484] = 9'b111111111;
assign micromatrizz[50][485] = 9'b111111111;
assign micromatrizz[50][486] = 9'b111111111;
assign micromatrizz[50][487] = 9'b111111111;
assign micromatrizz[50][488] = 9'b111111111;
assign micromatrizz[50][489] = 9'b111111111;
assign micromatrizz[50][490] = 9'b111111111;
assign micromatrizz[50][491] = 9'b111111111;
assign micromatrizz[50][492] = 9'b111111111;
assign micromatrizz[50][493] = 9'b111111111;
assign micromatrizz[50][494] = 9'b111111111;
assign micromatrizz[50][495] = 9'b111111111;
assign micromatrizz[50][496] = 9'b111111111;
assign micromatrizz[50][497] = 9'b111111111;
assign micromatrizz[50][498] = 9'b111111111;
assign micromatrizz[50][499] = 9'b111111111;
assign micromatrizz[50][500] = 9'b111111111;
assign micromatrizz[50][501] = 9'b111111111;
assign micromatrizz[50][502] = 9'b111111111;
assign micromatrizz[50][503] = 9'b111111111;
assign micromatrizz[50][504] = 9'b111111111;
assign micromatrizz[50][505] = 9'b111111111;
assign micromatrizz[50][506] = 9'b111111111;
assign micromatrizz[50][507] = 9'b111111111;
assign micromatrizz[50][508] = 9'b111111111;
assign micromatrizz[50][509] = 9'b111111111;
assign micromatrizz[50][510] = 9'b111111111;
assign micromatrizz[50][511] = 9'b111111111;
assign micromatrizz[50][512] = 9'b111111111;
assign micromatrizz[50][513] = 9'b111111111;
assign micromatrizz[50][514] = 9'b111111111;
assign micromatrizz[50][515] = 9'b111111111;
assign micromatrizz[50][516] = 9'b111110111;
assign micromatrizz[50][517] = 9'b111110011;
assign micromatrizz[50][518] = 9'b111110011;
assign micromatrizz[50][519] = 9'b111110011;
assign micromatrizz[50][520] = 9'b111110010;
assign micromatrizz[50][521] = 9'b111110010;
assign micromatrizz[50][522] = 9'b111110011;
assign micromatrizz[50][523] = 9'b111110111;
assign micromatrizz[50][524] = 9'b111111111;
assign micromatrizz[50][525] = 9'b111111111;
assign micromatrizz[50][526] = 9'b111111111;
assign micromatrizz[50][527] = 9'b111111111;
assign micromatrizz[50][528] = 9'b111111111;
assign micromatrizz[50][529] = 9'b111111111;
assign micromatrizz[50][530] = 9'b111111111;
assign micromatrizz[50][531] = 9'b111111111;
assign micromatrizz[50][532] = 9'b111111111;
assign micromatrizz[50][533] = 9'b111111111;
assign micromatrizz[50][534] = 9'b111111111;
assign micromatrizz[50][535] = 9'b111111111;
assign micromatrizz[50][536] = 9'b111111111;
assign micromatrizz[50][537] = 9'b111111111;
assign micromatrizz[50][538] = 9'b111111111;
assign micromatrizz[50][539] = 9'b111111111;
assign micromatrizz[50][540] = 9'b111111111;
assign micromatrizz[50][541] = 9'b111111111;
assign micromatrizz[50][542] = 9'b111111111;
assign micromatrizz[50][543] = 9'b111111111;
assign micromatrizz[50][544] = 9'b111111111;
assign micromatrizz[50][545] = 9'b111111111;
assign micromatrizz[50][546] = 9'b111111111;
assign micromatrizz[50][547] = 9'b111111111;
assign micromatrizz[50][548] = 9'b111111111;
assign micromatrizz[50][549] = 9'b111111111;
assign micromatrizz[50][550] = 9'b111111111;
assign micromatrizz[50][551] = 9'b111111111;
assign micromatrizz[50][552] = 9'b111111111;
assign micromatrizz[50][553] = 9'b111111111;
assign micromatrizz[50][554] = 9'b111111111;
assign micromatrizz[50][555] = 9'b111111111;
assign micromatrizz[50][556] = 9'b111111111;
assign micromatrizz[50][557] = 9'b111111111;
assign micromatrizz[50][558] = 9'b111110010;
assign micromatrizz[50][559] = 9'b111110010;
assign micromatrizz[50][560] = 9'b111110010;
assign micromatrizz[50][561] = 9'b111110010;
assign micromatrizz[50][562] = 9'b111110011;
assign micromatrizz[50][563] = 9'b111110011;
assign micromatrizz[50][564] = 9'b111110011;
assign micromatrizz[50][565] = 9'b111111111;
assign micromatrizz[50][566] = 9'b111111111;
assign micromatrizz[50][567] = 9'b111111111;
assign micromatrizz[50][568] = 9'b111111111;
assign micromatrizz[50][569] = 9'b111111111;
assign micromatrizz[50][570] = 9'b111111111;
assign micromatrizz[50][571] = 9'b111111111;
assign micromatrizz[50][572] = 9'b111111111;
assign micromatrizz[50][573] = 9'b111111111;
assign micromatrizz[50][574] = 9'b111111111;
assign micromatrizz[50][575] = 9'b111111111;
assign micromatrizz[50][576] = 9'b111111111;
assign micromatrizz[50][577] = 9'b111111111;
assign micromatrizz[50][578] = 9'b111111111;
assign micromatrizz[50][579] = 9'b111111111;
assign micromatrizz[50][580] = 9'b111111111;
assign micromatrizz[50][581] = 9'b111110010;
assign micromatrizz[50][582] = 9'b111110011;
assign micromatrizz[50][583] = 9'b111110011;
assign micromatrizz[50][584] = 9'b111110010;
assign micromatrizz[50][585] = 9'b111110010;
assign micromatrizz[50][586] = 9'b111110010;
assign micromatrizz[50][587] = 9'b111110011;
assign micromatrizz[50][588] = 9'b111111111;
assign micromatrizz[50][589] = 9'b111111111;
assign micromatrizz[50][590] = 9'b111111111;
assign micromatrizz[50][591] = 9'b111111111;
assign micromatrizz[50][592] = 9'b111111111;
assign micromatrizz[50][593] = 9'b111111111;
assign micromatrizz[50][594] = 9'b111111111;
assign micromatrizz[50][595] = 9'b111111111;
assign micromatrizz[50][596] = 9'b111111111;
assign micromatrizz[50][597] = 9'b111111111;
assign micromatrizz[50][598] = 9'b111111111;
assign micromatrizz[50][599] = 9'b111111111;
assign micromatrizz[50][600] = 9'b111111111;
assign micromatrizz[50][601] = 9'b111111111;
assign micromatrizz[50][602] = 9'b111111111;
assign micromatrizz[50][603] = 9'b111111111;
assign micromatrizz[50][604] = 9'b111111111;
assign micromatrizz[50][605] = 9'b111111111;
assign micromatrizz[50][606] = 9'b111111111;
assign micromatrizz[50][607] = 9'b111111111;
assign micromatrizz[50][608] = 9'b111111111;
assign micromatrizz[50][609] = 9'b111111111;
assign micromatrizz[50][610] = 9'b111111111;
assign micromatrizz[50][611] = 9'b111111111;
assign micromatrizz[50][612] = 9'b111111111;
assign micromatrizz[50][613] = 9'b111111111;
assign micromatrizz[50][614] = 9'b111111111;
assign micromatrizz[50][615] = 9'b111111111;
assign micromatrizz[50][616] = 9'b111111111;
assign micromatrizz[50][617] = 9'b111111111;
assign micromatrizz[50][618] = 9'b111111111;
assign micromatrizz[50][619] = 9'b111111111;
assign micromatrizz[50][620] = 9'b111111111;
assign micromatrizz[50][621] = 9'b111111111;
assign micromatrizz[50][622] = 9'b111111111;
assign micromatrizz[50][623] = 9'b111111111;
assign micromatrizz[50][624] = 9'b111111111;
assign micromatrizz[50][625] = 9'b111111111;
assign micromatrizz[50][626] = 9'b111111111;
assign micromatrizz[50][627] = 9'b111111111;
assign micromatrizz[50][628] = 9'b111111111;
assign micromatrizz[50][629] = 9'b111111111;
assign micromatrizz[50][630] = 9'b111111111;
assign micromatrizz[50][631] = 9'b111111111;
assign micromatrizz[50][632] = 9'b111111111;
assign micromatrizz[50][633] = 9'b111111111;
assign micromatrizz[50][634] = 9'b111111111;
assign micromatrizz[50][635] = 9'b111111111;
assign micromatrizz[50][636] = 9'b111111111;
assign micromatrizz[50][637] = 9'b111111111;
assign micromatrizz[50][638] = 9'b111111111;
assign micromatrizz[50][639] = 9'b111111111;
assign micromatrizz[51][0] = 9'b111111111;
assign micromatrizz[51][1] = 9'b111111111;
assign micromatrizz[51][2] = 9'b111111111;
assign micromatrizz[51][3] = 9'b111111111;
assign micromatrizz[51][4] = 9'b111111111;
assign micromatrizz[51][5] = 9'b111111111;
assign micromatrizz[51][6] = 9'b111111111;
assign micromatrizz[51][7] = 9'b111111111;
assign micromatrizz[51][8] = 9'b111111111;
assign micromatrizz[51][9] = 9'b111111111;
assign micromatrizz[51][10] = 9'b111111111;
assign micromatrizz[51][11] = 9'b111111111;
assign micromatrizz[51][12] = 9'b111111111;
assign micromatrizz[51][13] = 9'b111111111;
assign micromatrizz[51][14] = 9'b111111111;
assign micromatrizz[51][15] = 9'b111111111;
assign micromatrizz[51][16] = 9'b111111111;
assign micromatrizz[51][17] = 9'b111111111;
assign micromatrizz[51][18] = 9'b111111111;
assign micromatrizz[51][19] = 9'b111111111;
assign micromatrizz[51][20] = 9'b111111111;
assign micromatrizz[51][21] = 9'b111111111;
assign micromatrizz[51][22] = 9'b111111111;
assign micromatrizz[51][23] = 9'b111111111;
assign micromatrizz[51][24] = 9'b111111111;
assign micromatrizz[51][25] = 9'b111111111;
assign micromatrizz[51][26] = 9'b111111111;
assign micromatrizz[51][27] = 9'b111111111;
assign micromatrizz[51][28] = 9'b111111111;
assign micromatrizz[51][29] = 9'b111111111;
assign micromatrizz[51][30] = 9'b111111111;
assign micromatrizz[51][31] = 9'b111111111;
assign micromatrizz[51][32] = 9'b111111111;
assign micromatrizz[51][33] = 9'b111111111;
assign micromatrizz[51][34] = 9'b111111111;
assign micromatrizz[51][35] = 9'b111111111;
assign micromatrizz[51][36] = 9'b111111111;
assign micromatrizz[51][37] = 9'b111111111;
assign micromatrizz[51][38] = 9'b111111111;
assign micromatrizz[51][39] = 9'b111111111;
assign micromatrizz[51][40] = 9'b111111111;
assign micromatrizz[51][41] = 9'b111111111;
assign micromatrizz[51][42] = 9'b111111111;
assign micromatrizz[51][43] = 9'b111111111;
assign micromatrizz[51][44] = 9'b111111111;
assign micromatrizz[51][45] = 9'b111111111;
assign micromatrizz[51][46] = 9'b111111111;
assign micromatrizz[51][47] = 9'b111111111;
assign micromatrizz[51][48] = 9'b111111111;
assign micromatrizz[51][49] = 9'b111111111;
assign micromatrizz[51][50] = 9'b111111111;
assign micromatrizz[51][51] = 9'b111111111;
assign micromatrizz[51][52] = 9'b111111111;
assign micromatrizz[51][53] = 9'b111111111;
assign micromatrizz[51][54] = 9'b111111111;
assign micromatrizz[51][55] = 9'b111111111;
assign micromatrizz[51][56] = 9'b111111111;
assign micromatrizz[51][57] = 9'b111111111;
assign micromatrizz[51][58] = 9'b111111111;
assign micromatrizz[51][59] = 9'b111111111;
assign micromatrizz[51][60] = 9'b111111111;
assign micromatrizz[51][61] = 9'b111111111;
assign micromatrizz[51][62] = 9'b111111111;
assign micromatrizz[51][63] = 9'b111111111;
assign micromatrizz[51][64] = 9'b111111111;
assign micromatrizz[51][65] = 9'b111111111;
assign micromatrizz[51][66] = 9'b111111111;
assign micromatrizz[51][67] = 9'b111111111;
assign micromatrizz[51][68] = 9'b111111111;
assign micromatrizz[51][69] = 9'b111111111;
assign micromatrizz[51][70] = 9'b111111111;
assign micromatrizz[51][71] = 9'b111111111;
assign micromatrizz[51][72] = 9'b111111111;
assign micromatrizz[51][73] = 9'b111111111;
assign micromatrizz[51][74] = 9'b111111111;
assign micromatrizz[51][75] = 9'b111111111;
assign micromatrizz[51][76] = 9'b111111111;
assign micromatrizz[51][77] = 9'b111111111;
assign micromatrizz[51][78] = 9'b111111111;
assign micromatrizz[51][79] = 9'b111111111;
assign micromatrizz[51][80] = 9'b111111111;
assign micromatrizz[51][81] = 9'b111111111;
assign micromatrizz[51][82] = 9'b111111111;
assign micromatrizz[51][83] = 9'b111111111;
assign micromatrizz[51][84] = 9'b111111111;
assign micromatrizz[51][85] = 9'b111111111;
assign micromatrizz[51][86] = 9'b111111111;
assign micromatrizz[51][87] = 9'b111111111;
assign micromatrizz[51][88] = 9'b111111111;
assign micromatrizz[51][89] = 9'b111111111;
assign micromatrizz[51][90] = 9'b111111111;
assign micromatrizz[51][91] = 9'b111111111;
assign micromatrizz[51][92] = 9'b111111111;
assign micromatrizz[51][93] = 9'b111111111;
assign micromatrizz[51][94] = 9'b111111111;
assign micromatrizz[51][95] = 9'b111111111;
assign micromatrizz[51][96] = 9'b111111111;
assign micromatrizz[51][97] = 9'b111111111;
assign micromatrizz[51][98] = 9'b111111111;
assign micromatrizz[51][99] = 9'b111111111;
assign micromatrizz[51][100] = 9'b111111111;
assign micromatrizz[51][101] = 9'b111111111;
assign micromatrizz[51][102] = 9'b111111111;
assign micromatrizz[51][103] = 9'b111111111;
assign micromatrizz[51][104] = 9'b111111111;
assign micromatrizz[51][105] = 9'b111111111;
assign micromatrizz[51][106] = 9'b111111111;
assign micromatrizz[51][107] = 9'b111111111;
assign micromatrizz[51][108] = 9'b111111111;
assign micromatrizz[51][109] = 9'b111111111;
assign micromatrizz[51][110] = 9'b111111111;
assign micromatrizz[51][111] = 9'b111111111;
assign micromatrizz[51][112] = 9'b111111111;
assign micromatrizz[51][113] = 9'b111111111;
assign micromatrizz[51][114] = 9'b111111111;
assign micromatrizz[51][115] = 9'b111111111;
assign micromatrizz[51][116] = 9'b111111111;
assign micromatrizz[51][117] = 9'b111111111;
assign micromatrizz[51][118] = 9'b111111111;
assign micromatrizz[51][119] = 9'b111111111;
assign micromatrizz[51][120] = 9'b111111111;
assign micromatrizz[51][121] = 9'b111111111;
assign micromatrizz[51][122] = 9'b111111111;
assign micromatrizz[51][123] = 9'b111111111;
assign micromatrizz[51][124] = 9'b111111111;
assign micromatrizz[51][125] = 9'b111111111;
assign micromatrizz[51][126] = 9'b111111111;
assign micromatrizz[51][127] = 9'b111111111;
assign micromatrizz[51][128] = 9'b111111111;
assign micromatrizz[51][129] = 9'b111111111;
assign micromatrizz[51][130] = 9'b111111111;
assign micromatrizz[51][131] = 9'b111111111;
assign micromatrizz[51][132] = 9'b111111111;
assign micromatrizz[51][133] = 9'b111111111;
assign micromatrizz[51][134] = 9'b111111111;
assign micromatrizz[51][135] = 9'b111111111;
assign micromatrizz[51][136] = 9'b111111111;
assign micromatrizz[51][137] = 9'b111111111;
assign micromatrizz[51][138] = 9'b111111111;
assign micromatrizz[51][139] = 9'b111111111;
assign micromatrizz[51][140] = 9'b111111111;
assign micromatrizz[51][141] = 9'b111111111;
assign micromatrizz[51][142] = 9'b111111111;
assign micromatrizz[51][143] = 9'b111111111;
assign micromatrizz[51][144] = 9'b111111111;
assign micromatrizz[51][145] = 9'b111111111;
assign micromatrizz[51][146] = 9'b111111111;
assign micromatrizz[51][147] = 9'b111111111;
assign micromatrizz[51][148] = 9'b111111111;
assign micromatrizz[51][149] = 9'b111111111;
assign micromatrizz[51][150] = 9'b111111111;
assign micromatrizz[51][151] = 9'b111111111;
assign micromatrizz[51][152] = 9'b111111111;
assign micromatrizz[51][153] = 9'b111111111;
assign micromatrizz[51][154] = 9'b111111111;
assign micromatrizz[51][155] = 9'b111111111;
assign micromatrizz[51][156] = 9'b111111111;
assign micromatrizz[51][157] = 9'b111111111;
assign micromatrizz[51][158] = 9'b111111111;
assign micromatrizz[51][159] = 9'b111111111;
assign micromatrizz[51][160] = 9'b111111111;
assign micromatrizz[51][161] = 9'b111111111;
assign micromatrizz[51][162] = 9'b111111111;
assign micromatrizz[51][163] = 9'b111111111;
assign micromatrizz[51][164] = 9'b111111111;
assign micromatrizz[51][165] = 9'b111111111;
assign micromatrizz[51][166] = 9'b111111111;
assign micromatrizz[51][167] = 9'b111111111;
assign micromatrizz[51][168] = 9'b111111111;
assign micromatrizz[51][169] = 9'b111111111;
assign micromatrizz[51][170] = 9'b111111111;
assign micromatrizz[51][171] = 9'b111111111;
assign micromatrizz[51][172] = 9'b111111111;
assign micromatrizz[51][173] = 9'b111111111;
assign micromatrizz[51][174] = 9'b111111111;
assign micromatrizz[51][175] = 9'b111111111;
assign micromatrizz[51][176] = 9'b111111111;
assign micromatrizz[51][177] = 9'b111111111;
assign micromatrizz[51][178] = 9'b111111111;
assign micromatrizz[51][179] = 9'b111111111;
assign micromatrizz[51][180] = 9'b111111111;
assign micromatrizz[51][181] = 9'b111111111;
assign micromatrizz[51][182] = 9'b111111111;
assign micromatrizz[51][183] = 9'b111111111;
assign micromatrizz[51][184] = 9'b111111111;
assign micromatrizz[51][185] = 9'b111111111;
assign micromatrizz[51][186] = 9'b111111111;
assign micromatrizz[51][187] = 9'b111111111;
assign micromatrizz[51][188] = 9'b111111111;
assign micromatrizz[51][189] = 9'b111111111;
assign micromatrizz[51][190] = 9'b111111111;
assign micromatrizz[51][191] = 9'b111111111;
assign micromatrizz[51][192] = 9'b111111111;
assign micromatrizz[51][193] = 9'b111111111;
assign micromatrizz[51][194] = 9'b111111111;
assign micromatrizz[51][195] = 9'b111110010;
assign micromatrizz[51][196] = 9'b111110010;
assign micromatrizz[51][197] = 9'b111110011;
assign micromatrizz[51][198] = 9'b111110011;
assign micromatrizz[51][199] = 9'b111110010;
assign micromatrizz[51][200] = 9'b111110010;
assign micromatrizz[51][201] = 9'b111110011;
assign micromatrizz[51][202] = 9'b111110111;
assign micromatrizz[51][203] = 9'b111111111;
assign micromatrizz[51][204] = 9'b111111111;
assign micromatrizz[51][205] = 9'b111111111;
assign micromatrizz[51][206] = 9'b111111111;
assign micromatrizz[51][207] = 9'b111111111;
assign micromatrizz[51][208] = 9'b111111111;
assign micromatrizz[51][209] = 9'b111111111;
assign micromatrizz[51][210] = 9'b111111111;
assign micromatrizz[51][211] = 9'b111111111;
assign micromatrizz[51][212] = 9'b111111111;
assign micromatrizz[51][213] = 9'b111111111;
assign micromatrizz[51][214] = 9'b111111111;
assign micromatrizz[51][215] = 9'b111111111;
assign micromatrizz[51][216] = 9'b111111111;
assign micromatrizz[51][217] = 9'b111111111;
assign micromatrizz[51][218] = 9'b111111111;
assign micromatrizz[51][219] = 9'b111111111;
assign micromatrizz[51][220] = 9'b111111111;
assign micromatrizz[51][221] = 9'b111111111;
assign micromatrizz[51][222] = 9'b111111111;
assign micromatrizz[51][223] = 9'b111111111;
assign micromatrizz[51][224] = 9'b111111111;
assign micromatrizz[51][225] = 9'b111111111;
assign micromatrizz[51][226] = 9'b111111111;
assign micromatrizz[51][227] = 9'b111111111;
assign micromatrizz[51][228] = 9'b111111111;
assign micromatrizz[51][229] = 9'b111111111;
assign micromatrizz[51][230] = 9'b111111111;
assign micromatrizz[51][231] = 9'b111111111;
assign micromatrizz[51][232] = 9'b111111111;
assign micromatrizz[51][233] = 9'b111111111;
assign micromatrizz[51][234] = 9'b111111111;
assign micromatrizz[51][235] = 9'b111111111;
assign micromatrizz[51][236] = 9'b111111111;
assign micromatrizz[51][237] = 9'b111111111;
assign micromatrizz[51][238] = 9'b111111111;
assign micromatrizz[51][239] = 9'b111111111;
assign micromatrizz[51][240] = 9'b111111111;
assign micromatrizz[51][241] = 9'b111111111;
assign micromatrizz[51][242] = 9'b111111111;
assign micromatrizz[51][243] = 9'b111111111;
assign micromatrizz[51][244] = 9'b111111111;
assign micromatrizz[51][245] = 9'b111111111;
assign micromatrizz[51][246] = 9'b111111111;
assign micromatrizz[51][247] = 9'b111111111;
assign micromatrizz[51][248] = 9'b111111111;
assign micromatrizz[51][249] = 9'b111111111;
assign micromatrizz[51][250] = 9'b111111111;
assign micromatrizz[51][251] = 9'b111111111;
assign micromatrizz[51][252] = 9'b111111111;
assign micromatrizz[51][253] = 9'b111111111;
assign micromatrizz[51][254] = 9'b111111111;
assign micromatrizz[51][255] = 9'b111111111;
assign micromatrizz[51][256] = 9'b111111111;
assign micromatrizz[51][257] = 9'b111111111;
assign micromatrizz[51][258] = 9'b111111111;
assign micromatrizz[51][259] = 9'b111111111;
assign micromatrizz[51][260] = 9'b111111111;
assign micromatrizz[51][261] = 9'b111111111;
assign micromatrizz[51][262] = 9'b111111111;
assign micromatrizz[51][263] = 9'b111111111;
assign micromatrizz[51][264] = 9'b111111111;
assign micromatrizz[51][265] = 9'b111111111;
assign micromatrizz[51][266] = 9'b111111111;
assign micromatrizz[51][267] = 9'b111111111;
assign micromatrizz[51][268] = 9'b111111111;
assign micromatrizz[51][269] = 9'b111111111;
assign micromatrizz[51][270] = 9'b111111111;
assign micromatrizz[51][271] = 9'b111111111;
assign micromatrizz[51][272] = 9'b111111111;
assign micromatrizz[51][273] = 9'b111111111;
assign micromatrizz[51][274] = 9'b111111111;
assign micromatrizz[51][275] = 9'b111111111;
assign micromatrizz[51][276] = 9'b111111111;
assign micromatrizz[51][277] = 9'b111111111;
assign micromatrizz[51][278] = 9'b111111111;
assign micromatrizz[51][279] = 9'b111111111;
assign micromatrizz[51][280] = 9'b111111111;
assign micromatrizz[51][281] = 9'b111111111;
assign micromatrizz[51][282] = 9'b111111111;
assign micromatrizz[51][283] = 9'b111111111;
assign micromatrizz[51][284] = 9'b111111111;
assign micromatrizz[51][285] = 9'b111111111;
assign micromatrizz[51][286] = 9'b111111111;
assign micromatrizz[51][287] = 9'b111111111;
assign micromatrizz[51][288] = 9'b111111111;
assign micromatrizz[51][289] = 9'b111111111;
assign micromatrizz[51][290] = 9'b111111111;
assign micromatrizz[51][291] = 9'b111111111;
assign micromatrizz[51][292] = 9'b111111111;
assign micromatrizz[51][293] = 9'b111111111;
assign micromatrizz[51][294] = 9'b111111111;
assign micromatrizz[51][295] = 9'b111111111;
assign micromatrizz[51][296] = 9'b111111111;
assign micromatrizz[51][297] = 9'b111111111;
assign micromatrizz[51][298] = 9'b111111111;
assign micromatrizz[51][299] = 9'b111111111;
assign micromatrizz[51][300] = 9'b111111111;
assign micromatrizz[51][301] = 9'b111111111;
assign micromatrizz[51][302] = 9'b111111111;
assign micromatrizz[51][303] = 9'b111111111;
assign micromatrizz[51][304] = 9'b111111111;
assign micromatrizz[51][305] = 9'b111111111;
assign micromatrizz[51][306] = 9'b111111111;
assign micromatrizz[51][307] = 9'b111111111;
assign micromatrizz[51][308] = 9'b111111111;
assign micromatrizz[51][309] = 9'b111111111;
assign micromatrizz[51][310] = 9'b111111111;
assign micromatrizz[51][311] = 9'b111111111;
assign micromatrizz[51][312] = 9'b111111111;
assign micromatrizz[51][313] = 9'b111111111;
assign micromatrizz[51][314] = 9'b111111111;
assign micromatrizz[51][315] = 9'b111111111;
assign micromatrizz[51][316] = 9'b111111111;
assign micromatrizz[51][317] = 9'b111111111;
assign micromatrizz[51][318] = 9'b111111111;
assign micromatrizz[51][319] = 9'b111111111;
assign micromatrizz[51][320] = 9'b111111111;
assign micromatrizz[51][321] = 9'b111111111;
assign micromatrizz[51][322] = 9'b111111111;
assign micromatrizz[51][323] = 9'b111111111;
assign micromatrizz[51][324] = 9'b111111111;
assign micromatrizz[51][325] = 9'b111111111;
assign micromatrizz[51][326] = 9'b111111111;
assign micromatrizz[51][327] = 9'b111111111;
assign micromatrizz[51][328] = 9'b111111111;
assign micromatrizz[51][329] = 9'b111111111;
assign micromatrizz[51][330] = 9'b111111111;
assign micromatrizz[51][331] = 9'b111111111;
assign micromatrizz[51][332] = 9'b111111111;
assign micromatrizz[51][333] = 9'b111111111;
assign micromatrizz[51][334] = 9'b111111111;
assign micromatrizz[51][335] = 9'b111111111;
assign micromatrizz[51][336] = 9'b111111111;
assign micromatrizz[51][337] = 9'b111111111;
assign micromatrizz[51][338] = 9'b111111111;
assign micromatrizz[51][339] = 9'b111111111;
assign micromatrizz[51][340] = 9'b111111111;
assign micromatrizz[51][341] = 9'b111111111;
assign micromatrizz[51][342] = 9'b111111111;
assign micromatrizz[51][343] = 9'b111111111;
assign micromatrizz[51][344] = 9'b111111111;
assign micromatrizz[51][345] = 9'b111111111;
assign micromatrizz[51][346] = 9'b111111111;
assign micromatrizz[51][347] = 9'b111111111;
assign micromatrizz[51][348] = 9'b111111111;
assign micromatrizz[51][349] = 9'b111111111;
assign micromatrizz[51][350] = 9'b111111111;
assign micromatrizz[51][351] = 9'b111111111;
assign micromatrizz[51][352] = 9'b111111111;
assign micromatrizz[51][353] = 9'b111111111;
assign micromatrizz[51][354] = 9'b111111111;
assign micromatrizz[51][355] = 9'b111111111;
assign micromatrizz[51][356] = 9'b111111111;
assign micromatrizz[51][357] = 9'b111111111;
assign micromatrizz[51][358] = 9'b111110111;
assign micromatrizz[51][359] = 9'b111110010;
assign micromatrizz[51][360] = 9'b111110011;
assign micromatrizz[51][361] = 9'b111110011;
assign micromatrizz[51][362] = 9'b111110010;
assign micromatrizz[51][363] = 9'b111110010;
assign micromatrizz[51][364] = 9'b111110011;
assign micromatrizz[51][365] = 9'b111110010;
assign micromatrizz[51][366] = 9'b111111111;
assign micromatrizz[51][367] = 9'b111111111;
assign micromatrizz[51][368] = 9'b111111111;
assign micromatrizz[51][369] = 9'b111111111;
assign micromatrizz[51][370] = 9'b111111111;
assign micromatrizz[51][371] = 9'b111111111;
assign micromatrizz[51][372] = 9'b111111111;
assign micromatrizz[51][373] = 9'b111111111;
assign micromatrizz[51][374] = 9'b111111111;
assign micromatrizz[51][375] = 9'b111111111;
assign micromatrizz[51][376] = 9'b111111111;
assign micromatrizz[51][377] = 9'b111111111;
assign micromatrizz[51][378] = 9'b111111111;
assign micromatrizz[51][379] = 9'b111111111;
assign micromatrizz[51][380] = 9'b111111111;
assign micromatrizz[51][381] = 9'b111111111;
assign micromatrizz[51][382] = 9'b111111111;
assign micromatrizz[51][383] = 9'b111111111;
assign micromatrizz[51][384] = 9'b111111111;
assign micromatrizz[51][385] = 9'b111111111;
assign micromatrizz[51][386] = 9'b111111111;
assign micromatrizz[51][387] = 9'b111111111;
assign micromatrizz[51][388] = 9'b111111111;
assign micromatrizz[51][389] = 9'b111111111;
assign micromatrizz[51][390] = 9'b111111111;
assign micromatrizz[51][391] = 9'b111111111;
assign micromatrizz[51][392] = 9'b111111111;
assign micromatrizz[51][393] = 9'b111111111;
assign micromatrizz[51][394] = 9'b111111111;
assign micromatrizz[51][395] = 9'b111111111;
assign micromatrizz[51][396] = 9'b111111111;
assign micromatrizz[51][397] = 9'b111111111;
assign micromatrizz[51][398] = 9'b111111111;
assign micromatrizz[51][399] = 9'b111111111;
assign micromatrizz[51][400] = 9'b111111111;
assign micromatrizz[51][401] = 9'b111111111;
assign micromatrizz[51][402] = 9'b111111111;
assign micromatrizz[51][403] = 9'b111111111;
assign micromatrizz[51][404] = 9'b111111111;
assign micromatrizz[51][405] = 9'b111111111;
assign micromatrizz[51][406] = 9'b111111111;
assign micromatrizz[51][407] = 9'b111111111;
assign micromatrizz[51][408] = 9'b111111111;
assign micromatrizz[51][409] = 9'b111111111;
assign micromatrizz[51][410] = 9'b111111111;
assign micromatrizz[51][411] = 9'b111111111;
assign micromatrizz[51][412] = 9'b111111111;
assign micromatrizz[51][413] = 9'b111111111;
assign micromatrizz[51][414] = 9'b111111111;
assign micromatrizz[51][415] = 9'b111111111;
assign micromatrizz[51][416] = 9'b111111111;
assign micromatrizz[51][417] = 9'b111111111;
assign micromatrizz[51][418] = 9'b111111111;
assign micromatrizz[51][419] = 9'b111111111;
assign micromatrizz[51][420] = 9'b111111111;
assign micromatrizz[51][421] = 9'b111111111;
assign micromatrizz[51][422] = 9'b111111111;
assign micromatrizz[51][423] = 9'b111111111;
assign micromatrizz[51][424] = 9'b111111111;
assign micromatrizz[51][425] = 9'b111111111;
assign micromatrizz[51][426] = 9'b111111111;
assign micromatrizz[51][427] = 9'b111111111;
assign micromatrizz[51][428] = 9'b111111111;
assign micromatrizz[51][429] = 9'b111111111;
assign micromatrizz[51][430] = 9'b111111111;
assign micromatrizz[51][431] = 9'b111111111;
assign micromatrizz[51][432] = 9'b111111111;
assign micromatrizz[51][433] = 9'b111111111;
assign micromatrizz[51][434] = 9'b111111111;
assign micromatrizz[51][435] = 9'b111111111;
assign micromatrizz[51][436] = 9'b111111111;
assign micromatrizz[51][437] = 9'b111111111;
assign micromatrizz[51][438] = 9'b111111111;
assign micromatrizz[51][439] = 9'b111111111;
assign micromatrizz[51][440] = 9'b111111111;
assign micromatrizz[51][441] = 9'b111111111;
assign micromatrizz[51][442] = 9'b111111111;
assign micromatrizz[51][443] = 9'b111111111;
assign micromatrizz[51][444] = 9'b111111111;
assign micromatrizz[51][445] = 9'b111111111;
assign micromatrizz[51][446] = 9'b111111111;
assign micromatrizz[51][447] = 9'b111111111;
assign micromatrizz[51][448] = 9'b111111111;
assign micromatrizz[51][449] = 9'b111111111;
assign micromatrizz[51][450] = 9'b111111111;
assign micromatrizz[51][451] = 9'b111111111;
assign micromatrizz[51][452] = 9'b111111111;
assign micromatrizz[51][453] = 9'b111111111;
assign micromatrizz[51][454] = 9'b111111111;
assign micromatrizz[51][455] = 9'b111111111;
assign micromatrizz[51][456] = 9'b111111111;
assign micromatrizz[51][457] = 9'b111111111;
assign micromatrizz[51][458] = 9'b111111111;
assign micromatrizz[51][459] = 9'b111111111;
assign micromatrizz[51][460] = 9'b111111111;
assign micromatrizz[51][461] = 9'b111111111;
assign micromatrizz[51][462] = 9'b111111111;
assign micromatrizz[51][463] = 9'b111111111;
assign micromatrizz[51][464] = 9'b111111111;
assign micromatrizz[51][465] = 9'b111111111;
assign micromatrizz[51][466] = 9'b111111111;
assign micromatrizz[51][467] = 9'b111111111;
assign micromatrizz[51][468] = 9'b111111111;
assign micromatrizz[51][469] = 9'b111111111;
assign micromatrizz[51][470] = 9'b111111111;
assign micromatrizz[51][471] = 9'b111111111;
assign micromatrizz[51][472] = 9'b111111111;
assign micromatrizz[51][473] = 9'b111111111;
assign micromatrizz[51][474] = 9'b111111111;
assign micromatrizz[51][475] = 9'b111111111;
assign micromatrizz[51][476] = 9'b111111111;
assign micromatrizz[51][477] = 9'b111111111;
assign micromatrizz[51][478] = 9'b111111111;
assign micromatrizz[51][479] = 9'b111111111;
assign micromatrizz[51][480] = 9'b111111111;
assign micromatrizz[51][481] = 9'b111111111;
assign micromatrizz[51][482] = 9'b111111111;
assign micromatrizz[51][483] = 9'b111111111;
assign micromatrizz[51][484] = 9'b111111111;
assign micromatrizz[51][485] = 9'b111111111;
assign micromatrizz[51][486] = 9'b111111111;
assign micromatrizz[51][487] = 9'b111111111;
assign micromatrizz[51][488] = 9'b111111111;
assign micromatrizz[51][489] = 9'b111111111;
assign micromatrizz[51][490] = 9'b111111111;
assign micromatrizz[51][491] = 9'b111111111;
assign micromatrizz[51][492] = 9'b111111111;
assign micromatrizz[51][493] = 9'b111111111;
assign micromatrizz[51][494] = 9'b111111111;
assign micromatrizz[51][495] = 9'b111111111;
assign micromatrizz[51][496] = 9'b111111111;
assign micromatrizz[51][497] = 9'b111111111;
assign micromatrizz[51][498] = 9'b111111111;
assign micromatrizz[51][499] = 9'b111111111;
assign micromatrizz[51][500] = 9'b111111111;
assign micromatrizz[51][501] = 9'b111111111;
assign micromatrizz[51][502] = 9'b111111111;
assign micromatrizz[51][503] = 9'b111111111;
assign micromatrizz[51][504] = 9'b111111111;
assign micromatrizz[51][505] = 9'b111111111;
assign micromatrizz[51][506] = 9'b111111111;
assign micromatrizz[51][507] = 9'b111111111;
assign micromatrizz[51][508] = 9'b111111111;
assign micromatrizz[51][509] = 9'b111111111;
assign micromatrizz[51][510] = 9'b111111111;
assign micromatrizz[51][511] = 9'b111111111;
assign micromatrizz[51][512] = 9'b111111111;
assign micromatrizz[51][513] = 9'b111111111;
assign micromatrizz[51][514] = 9'b111111111;
assign micromatrizz[51][515] = 9'b111111111;
assign micromatrizz[51][516] = 9'b111110111;
assign micromatrizz[51][517] = 9'b111110010;
assign micromatrizz[51][518] = 9'b111110011;
assign micromatrizz[51][519] = 9'b111110011;
assign micromatrizz[51][520] = 9'b111110010;
assign micromatrizz[51][521] = 9'b111110010;
assign micromatrizz[51][522] = 9'b111110011;
assign micromatrizz[51][523] = 9'b111110111;
assign micromatrizz[51][524] = 9'b111111111;
assign micromatrizz[51][525] = 9'b111111111;
assign micromatrizz[51][526] = 9'b111111111;
assign micromatrizz[51][527] = 9'b111111111;
assign micromatrizz[51][528] = 9'b111111111;
assign micromatrizz[51][529] = 9'b111111111;
assign micromatrizz[51][530] = 9'b111111111;
assign micromatrizz[51][531] = 9'b111111111;
assign micromatrizz[51][532] = 9'b111111111;
assign micromatrizz[51][533] = 9'b111111111;
assign micromatrizz[51][534] = 9'b111111111;
assign micromatrizz[51][535] = 9'b111111111;
assign micromatrizz[51][536] = 9'b111111111;
assign micromatrizz[51][537] = 9'b111111111;
assign micromatrizz[51][538] = 9'b111111111;
assign micromatrizz[51][539] = 9'b111111111;
assign micromatrizz[51][540] = 9'b111111111;
assign micromatrizz[51][541] = 9'b111111111;
assign micromatrizz[51][542] = 9'b111111111;
assign micromatrizz[51][543] = 9'b111111111;
assign micromatrizz[51][544] = 9'b111111111;
assign micromatrizz[51][545] = 9'b111111111;
assign micromatrizz[51][546] = 9'b111111111;
assign micromatrizz[51][547] = 9'b111111111;
assign micromatrizz[51][548] = 9'b111111111;
assign micromatrizz[51][549] = 9'b111111111;
assign micromatrizz[51][550] = 9'b111111111;
assign micromatrizz[51][551] = 9'b111111111;
assign micromatrizz[51][552] = 9'b111111111;
assign micromatrizz[51][553] = 9'b111111111;
assign micromatrizz[51][554] = 9'b111111111;
assign micromatrizz[51][555] = 9'b111111111;
assign micromatrizz[51][556] = 9'b111111111;
assign micromatrizz[51][557] = 9'b111111111;
assign micromatrizz[51][558] = 9'b111110010;
assign micromatrizz[51][559] = 9'b111110010;
assign micromatrizz[51][560] = 9'b111110010;
assign micromatrizz[51][561] = 9'b111110010;
assign micromatrizz[51][562] = 9'b111110011;
assign micromatrizz[51][563] = 9'b111110011;
assign micromatrizz[51][564] = 9'b111110011;
assign micromatrizz[51][565] = 9'b111111111;
assign micromatrizz[51][566] = 9'b111111111;
assign micromatrizz[51][567] = 9'b111111111;
assign micromatrizz[51][568] = 9'b111111111;
assign micromatrizz[51][569] = 9'b111111111;
assign micromatrizz[51][570] = 9'b111111111;
assign micromatrizz[51][571] = 9'b111111111;
assign micromatrizz[51][572] = 9'b111111111;
assign micromatrizz[51][573] = 9'b111111111;
assign micromatrizz[51][574] = 9'b111111111;
assign micromatrizz[51][575] = 9'b111111111;
assign micromatrizz[51][576] = 9'b111111111;
assign micromatrizz[51][577] = 9'b111111111;
assign micromatrizz[51][578] = 9'b111111111;
assign micromatrizz[51][579] = 9'b111111111;
assign micromatrizz[51][580] = 9'b111111111;
assign micromatrizz[51][581] = 9'b111110010;
assign micromatrizz[51][582] = 9'b111110011;
assign micromatrizz[51][583] = 9'b111110011;
assign micromatrizz[51][584] = 9'b111110010;
assign micromatrizz[51][585] = 9'b111110010;
assign micromatrizz[51][586] = 9'b111110011;
assign micromatrizz[51][587] = 9'b111110011;
assign micromatrizz[51][588] = 9'b111111111;
assign micromatrizz[51][589] = 9'b111111111;
assign micromatrizz[51][590] = 9'b111111111;
assign micromatrizz[51][591] = 9'b111111111;
assign micromatrizz[51][592] = 9'b111111111;
assign micromatrizz[51][593] = 9'b111111111;
assign micromatrizz[51][594] = 9'b111111111;
assign micromatrizz[51][595] = 9'b111111111;
assign micromatrizz[51][596] = 9'b111111111;
assign micromatrizz[51][597] = 9'b111111111;
assign micromatrizz[51][598] = 9'b111111111;
assign micromatrizz[51][599] = 9'b111111111;
assign micromatrizz[51][600] = 9'b111111111;
assign micromatrizz[51][601] = 9'b111111111;
assign micromatrizz[51][602] = 9'b111111111;
assign micromatrizz[51][603] = 9'b111111111;
assign micromatrizz[51][604] = 9'b111111111;
assign micromatrizz[51][605] = 9'b111111111;
assign micromatrizz[51][606] = 9'b111111111;
assign micromatrizz[51][607] = 9'b111111111;
assign micromatrizz[51][608] = 9'b111111111;
assign micromatrizz[51][609] = 9'b111111111;
assign micromatrizz[51][610] = 9'b111111111;
assign micromatrizz[51][611] = 9'b111111111;
assign micromatrizz[51][612] = 9'b111111111;
assign micromatrizz[51][613] = 9'b111111111;
assign micromatrizz[51][614] = 9'b111111111;
assign micromatrizz[51][615] = 9'b111111111;
assign micromatrizz[51][616] = 9'b111111111;
assign micromatrizz[51][617] = 9'b111111111;
assign micromatrizz[51][618] = 9'b111111111;
assign micromatrizz[51][619] = 9'b111111111;
assign micromatrizz[51][620] = 9'b111111111;
assign micromatrizz[51][621] = 9'b111111111;
assign micromatrizz[51][622] = 9'b111111111;
assign micromatrizz[51][623] = 9'b111111111;
assign micromatrizz[51][624] = 9'b111111111;
assign micromatrizz[51][625] = 9'b111111111;
assign micromatrizz[51][626] = 9'b111111111;
assign micromatrizz[51][627] = 9'b111111111;
assign micromatrizz[51][628] = 9'b111111111;
assign micromatrizz[51][629] = 9'b111111111;
assign micromatrizz[51][630] = 9'b111111111;
assign micromatrizz[51][631] = 9'b111111111;
assign micromatrizz[51][632] = 9'b111111111;
assign micromatrizz[51][633] = 9'b111111111;
assign micromatrizz[51][634] = 9'b111111111;
assign micromatrizz[51][635] = 9'b111111111;
assign micromatrizz[51][636] = 9'b111111111;
assign micromatrizz[51][637] = 9'b111111111;
assign micromatrizz[51][638] = 9'b111111111;
assign micromatrizz[51][639] = 9'b111111111;
assign micromatrizz[52][0] = 9'b111111111;
assign micromatrizz[52][1] = 9'b111111111;
assign micromatrizz[52][2] = 9'b111111111;
assign micromatrizz[52][3] = 9'b111111111;
assign micromatrizz[52][4] = 9'b111111111;
assign micromatrizz[52][5] = 9'b111111111;
assign micromatrizz[52][6] = 9'b111111111;
assign micromatrizz[52][7] = 9'b111111111;
assign micromatrizz[52][8] = 9'b111111111;
assign micromatrizz[52][9] = 9'b111111111;
assign micromatrizz[52][10] = 9'b111111111;
assign micromatrizz[52][11] = 9'b111111111;
assign micromatrizz[52][12] = 9'b111110111;
assign micromatrizz[52][13] = 9'b111110111;
assign micromatrizz[52][14] = 9'b111110111;
assign micromatrizz[52][15] = 9'b111111111;
assign micromatrizz[52][16] = 9'b111110111;
assign micromatrizz[52][17] = 9'b111110111;
assign micromatrizz[52][18] = 9'b111111111;
assign micromatrizz[52][19] = 9'b111111111;
assign micromatrizz[52][20] = 9'b111111111;
assign micromatrizz[52][21] = 9'b111111111;
assign micromatrizz[52][22] = 9'b111111111;
assign micromatrizz[52][23] = 9'b111110111;
assign micromatrizz[52][24] = 9'b111110010;
assign micromatrizz[52][25] = 9'b111110010;
assign micromatrizz[52][26] = 9'b111110010;
assign micromatrizz[52][27] = 9'b111110011;
assign micromatrizz[52][28] = 9'b111110011;
assign micromatrizz[52][29] = 9'b111110011;
assign micromatrizz[52][30] = 9'b111110010;
assign micromatrizz[52][31] = 9'b111111111;
assign micromatrizz[52][32] = 9'b111111111;
assign micromatrizz[52][33] = 9'b111111111;
assign micromatrizz[52][34] = 9'b111111111;
assign micromatrizz[52][35] = 9'b111110111;
assign micromatrizz[52][36] = 9'b111110010;
assign micromatrizz[52][37] = 9'b111110010;
assign micromatrizz[52][38] = 9'b111110010;
assign micromatrizz[52][39] = 9'b111110010;
assign micromatrizz[52][40] = 9'b111110011;
assign micromatrizz[52][41] = 9'b111110011;
assign micromatrizz[52][42] = 9'b111110011;
assign micromatrizz[52][43] = 9'b111111111;
assign micromatrizz[52][44] = 9'b111111111;
assign micromatrizz[52][45] = 9'b111111111;
assign micromatrizz[52][46] = 9'b111111111;
assign micromatrizz[52][47] = 9'b111110110;
assign micromatrizz[52][48] = 9'b111110010;
assign micromatrizz[52][49] = 9'b111110010;
assign micromatrizz[52][50] = 9'b111110010;
assign micromatrizz[52][51] = 9'b111110011;
assign micromatrizz[52][52] = 9'b111110010;
assign micromatrizz[52][53] = 9'b111110010;
assign micromatrizz[52][54] = 9'b111110111;
assign micromatrizz[52][55] = 9'b111111111;
assign micromatrizz[52][56] = 9'b111111111;
assign micromatrizz[52][57] = 9'b111110111;
assign micromatrizz[52][58] = 9'b111110011;
assign micromatrizz[52][59] = 9'b111110011;
assign micromatrizz[52][60] = 9'b111110010;
assign micromatrizz[52][61] = 9'b111110011;
assign micromatrizz[52][62] = 9'b111110111;
assign micromatrizz[52][63] = 9'b111111111;
assign micromatrizz[52][64] = 9'b111111111;
assign micromatrizz[52][65] = 9'b111111111;
assign micromatrizz[52][66] = 9'b111111111;
assign micromatrizz[52][67] = 9'b111111111;
assign micromatrizz[52][68] = 9'b111111111;
assign micromatrizz[52][69] = 9'b111111111;
assign micromatrizz[52][70] = 9'b111111111;
assign micromatrizz[52][71] = 9'b111111111;
assign micromatrizz[52][72] = 9'b111111111;
assign micromatrizz[52][73] = 9'b111111111;
assign micromatrizz[52][74] = 9'b111110111;
assign micromatrizz[52][75] = 9'b111110111;
assign micromatrizz[52][76] = 9'b111110111;
assign micromatrizz[52][77] = 9'b111110111;
assign micromatrizz[52][78] = 9'b111110111;
assign micromatrizz[52][79] = 9'b111110111;
assign micromatrizz[52][80] = 9'b111111111;
assign micromatrizz[52][81] = 9'b111111111;
assign micromatrizz[52][82] = 9'b111111111;
assign micromatrizz[52][83] = 9'b111111111;
assign micromatrizz[52][84] = 9'b111111111;
assign micromatrizz[52][85] = 9'b111111111;
assign micromatrizz[52][86] = 9'b111111111;
assign micromatrizz[52][87] = 9'b111111111;
assign micromatrizz[52][88] = 9'b111110110;
assign micromatrizz[52][89] = 9'b111110010;
assign micromatrizz[52][90] = 9'b111110011;
assign micromatrizz[52][91] = 9'b111110010;
assign micromatrizz[52][92] = 9'b111110010;
assign micromatrizz[52][93] = 9'b111110011;
assign micromatrizz[52][94] = 9'b111110010;
assign micromatrizz[52][95] = 9'b111110111;
assign micromatrizz[52][96] = 9'b111111111;
assign micromatrizz[52][97] = 9'b111111111;
assign micromatrizz[52][98] = 9'b111111111;
assign micromatrizz[52][99] = 9'b111110111;
assign micromatrizz[52][100] = 9'b111110010;
assign micromatrizz[52][101] = 9'b111110011;
assign micromatrizz[52][102] = 9'b111111111;
assign micromatrizz[52][103] = 9'b111111111;
assign micromatrizz[52][104] = 9'b111111111;
assign micromatrizz[52][105] = 9'b111111111;
assign micromatrizz[52][106] = 9'b111111111;
assign micromatrizz[52][107] = 9'b111111111;
assign micromatrizz[52][108] = 9'b111110111;
assign micromatrizz[52][109] = 9'b111110111;
assign micromatrizz[52][110] = 9'b111110111;
assign micromatrizz[52][111] = 9'b111111111;
assign micromatrizz[52][112] = 9'b111110111;
assign micromatrizz[52][113] = 9'b111110111;
assign micromatrizz[52][114] = 9'b111111111;
assign micromatrizz[52][115] = 9'b111111111;
assign micromatrizz[52][116] = 9'b111111111;
assign micromatrizz[52][117] = 9'b111111111;
assign micromatrizz[52][118] = 9'b111111111;
assign micromatrizz[52][119] = 9'b111111111;
assign micromatrizz[52][120] = 9'b111111111;
assign micromatrizz[52][121] = 9'b111111111;
assign micromatrizz[52][122] = 9'b111111111;
assign micromatrizz[52][123] = 9'b111111111;
assign micromatrizz[52][124] = 9'b111111111;
assign micromatrizz[52][125] = 9'b111110111;
assign micromatrizz[52][126] = 9'b111110011;
assign micromatrizz[52][127] = 9'b111110111;
assign micromatrizz[52][128] = 9'b111110111;
assign micromatrizz[52][129] = 9'b111110111;
assign micromatrizz[52][130] = 9'b111111111;
assign micromatrizz[52][131] = 9'b111111111;
assign micromatrizz[52][132] = 9'b111111111;
assign micromatrizz[52][133] = 9'b111111111;
assign micromatrizz[52][134] = 9'b111111111;
assign micromatrizz[52][135] = 9'b111111111;
assign micromatrizz[52][136] = 9'b111111111;
assign micromatrizz[52][137] = 9'b111111111;
assign micromatrizz[52][138] = 9'b111110111;
assign micromatrizz[52][139] = 9'b111110010;
assign micromatrizz[52][140] = 9'b111110010;
assign micromatrizz[52][141] = 9'b111110011;
assign micromatrizz[52][142] = 9'b111110010;
assign micromatrizz[52][143] = 9'b111110110;
assign micromatrizz[52][144] = 9'b111110010;
assign micromatrizz[52][145] = 9'b111110111;
assign micromatrizz[52][146] = 9'b111111111;
assign micromatrizz[52][147] = 9'b111111111;
assign micromatrizz[52][148] = 9'b111111111;
assign micromatrizz[52][149] = 9'b111110111;
assign micromatrizz[52][150] = 9'b111110111;
assign micromatrizz[52][151] = 9'b111110010;
assign micromatrizz[52][152] = 9'b111110010;
assign micromatrizz[52][153] = 9'b111110010;
assign micromatrizz[52][154] = 9'b111110111;
assign micromatrizz[52][155] = 9'b111111111;
assign micromatrizz[52][156] = 9'b111111111;
assign micromatrizz[52][157] = 9'b111111111;
assign micromatrizz[52][158] = 9'b111111111;
assign micromatrizz[52][159] = 9'b111111111;
assign micromatrizz[52][160] = 9'b111111111;
assign micromatrizz[52][161] = 9'b111111111;
assign micromatrizz[52][162] = 9'b111111111;
assign micromatrizz[52][163] = 9'b111111111;
assign micromatrizz[52][164] = 9'b111111111;
assign micromatrizz[52][165] = 9'b111111111;
assign micromatrizz[52][166] = 9'b111110111;
assign micromatrizz[52][167] = 9'b111110111;
assign micromatrizz[52][168] = 9'b111110111;
assign micromatrizz[52][169] = 9'b111110111;
assign micromatrizz[52][170] = 9'b111110111;
assign micromatrizz[52][171] = 9'b111110110;
assign micromatrizz[52][172] = 9'b111110010;
assign micromatrizz[52][173] = 9'b111110111;
assign micromatrizz[52][174] = 9'b111110111;
assign micromatrizz[52][175] = 9'b111111111;
assign micromatrizz[52][176] = 9'b111111111;
assign micromatrizz[52][177] = 9'b111111111;
assign micromatrizz[52][178] = 9'b111111111;
assign micromatrizz[52][179] = 9'b111111111;
assign micromatrizz[52][180] = 9'b111111111;
assign micromatrizz[52][181] = 9'b111111111;
assign micromatrizz[52][182] = 9'b111111111;
assign micromatrizz[52][183] = 9'b111111111;
assign micromatrizz[52][184] = 9'b111111111;
assign micromatrizz[52][185] = 9'b111111111;
assign micromatrizz[52][186] = 9'b111111111;
assign micromatrizz[52][187] = 9'b111111111;
assign micromatrizz[52][188] = 9'b111110011;
assign micromatrizz[52][189] = 9'b111110011;
assign micromatrizz[52][190] = 9'b111110011;
assign micromatrizz[52][191] = 9'b111110011;
assign micromatrizz[52][192] = 9'b111111111;
assign micromatrizz[52][193] = 9'b111111111;
assign micromatrizz[52][194] = 9'b111111111;
assign micromatrizz[52][195] = 9'b111110010;
assign micromatrizz[52][196] = 9'b111110010;
assign micromatrizz[52][197] = 9'b111110011;
assign micromatrizz[52][198] = 9'b111110011;
assign micromatrizz[52][199] = 9'b111110010;
assign micromatrizz[52][200] = 9'b111110010;
assign micromatrizz[52][201] = 9'b111110011;
assign micromatrizz[52][202] = 9'b111110111;
assign micromatrizz[52][203] = 9'b111111111;
assign micromatrizz[52][204] = 9'b111111111;
assign micromatrizz[52][205] = 9'b111111111;
assign micromatrizz[52][206] = 9'b111111111;
assign micromatrizz[52][207] = 9'b111111111;
assign micromatrizz[52][208] = 9'b111111111;
assign micromatrizz[52][209] = 9'b111111111;
assign micromatrizz[52][210] = 9'b111111111;
assign micromatrizz[52][211] = 9'b111110111;
assign micromatrizz[52][212] = 9'b111110111;
assign micromatrizz[52][213] = 9'b111110111;
assign micromatrizz[52][214] = 9'b111110111;
assign micromatrizz[52][215] = 9'b111110111;
assign micromatrizz[52][216] = 9'b111110111;
assign micromatrizz[52][217] = 9'b111111111;
assign micromatrizz[52][218] = 9'b111111111;
assign micromatrizz[52][219] = 9'b111111111;
assign micromatrizz[52][220] = 9'b111111111;
assign micromatrizz[52][221] = 9'b111111111;
assign micromatrizz[52][222] = 9'b111111111;
assign micromatrizz[52][223] = 9'b111111111;
assign micromatrizz[52][224] = 9'b111111111;
assign micromatrizz[52][225] = 9'b111110111;
assign micromatrizz[52][226] = 9'b111110010;
assign micromatrizz[52][227] = 9'b111110010;
assign micromatrizz[52][228] = 9'b111110010;
assign micromatrizz[52][229] = 9'b111110010;
assign micromatrizz[52][230] = 9'b111110010;
assign micromatrizz[52][231] = 9'b111110010;
assign micromatrizz[52][232] = 9'b111110111;
assign micromatrizz[52][233] = 9'b111111111;
assign micromatrizz[52][234] = 9'b111111111;
assign micromatrizz[52][235] = 9'b111111111;
assign micromatrizz[52][236] = 9'b111110111;
assign micromatrizz[52][237] = 9'b111110010;
assign micromatrizz[52][238] = 9'b111110010;
assign micromatrizz[52][239] = 9'b111110111;
assign micromatrizz[52][240] = 9'b111111111;
assign micromatrizz[52][241] = 9'b111111111;
assign micromatrizz[52][242] = 9'b111111111;
assign micromatrizz[52][243] = 9'b111111111;
assign micromatrizz[52][244] = 9'b111111111;
assign micromatrizz[52][245] = 9'b111111111;
assign micromatrizz[52][246] = 9'b111110111;
assign micromatrizz[52][247] = 9'b111110111;
assign micromatrizz[52][248] = 9'b111110111;
assign micromatrizz[52][249] = 9'b111110111;
assign micromatrizz[52][250] = 9'b111110111;
assign micromatrizz[52][251] = 9'b111110111;
assign micromatrizz[52][252] = 9'b111111111;
assign micromatrizz[52][253] = 9'b111111111;
assign micromatrizz[52][254] = 9'b111111111;
assign micromatrizz[52][255] = 9'b111111111;
assign micromatrizz[52][256] = 9'b111111111;
assign micromatrizz[52][257] = 9'b111111111;
assign micromatrizz[52][258] = 9'b111111111;
assign micromatrizz[52][259] = 9'b111111111;
assign micromatrizz[52][260] = 9'b111111111;
assign micromatrizz[52][261] = 9'b111111111;
assign micromatrizz[52][262] = 9'b111111111;
assign micromatrizz[52][263] = 9'b111110111;
assign micromatrizz[52][264] = 9'b111110111;
assign micromatrizz[52][265] = 9'b111110111;
assign micromatrizz[52][266] = 9'b111110111;
assign micromatrizz[52][267] = 9'b111110111;
assign micromatrizz[52][268] = 9'b111110111;
assign micromatrizz[52][269] = 9'b111110111;
assign micromatrizz[52][270] = 9'b111111111;
assign micromatrizz[52][271] = 9'b111111111;
assign micromatrizz[52][272] = 9'b111111111;
assign micromatrizz[52][273] = 9'b111111111;
assign micromatrizz[52][274] = 9'b111111111;
assign micromatrizz[52][275] = 9'b111111111;
assign micromatrizz[52][276] = 9'b111111111;
assign micromatrizz[52][277] = 9'b111111111;
assign micromatrizz[52][278] = 9'b111111111;
assign micromatrizz[52][279] = 9'b111111111;
assign micromatrizz[52][280] = 9'b111110111;
assign micromatrizz[52][281] = 9'b111110111;
assign micromatrizz[52][282] = 9'b111111111;
assign micromatrizz[52][283] = 9'b111111111;
assign micromatrizz[52][284] = 9'b111110111;
assign micromatrizz[52][285] = 9'b111110010;
assign micromatrizz[52][286] = 9'b111110011;
assign micromatrizz[52][287] = 9'b111110111;
assign micromatrizz[52][288] = 9'b111110111;
assign micromatrizz[52][289] = 9'b111111111;
assign micromatrizz[52][290] = 9'b111111111;
assign micromatrizz[52][291] = 9'b111111111;
assign micromatrizz[52][292] = 9'b111111111;
assign micromatrizz[52][293] = 9'b111111111;
assign micromatrizz[52][294] = 9'b111111111;
assign micromatrizz[52][295] = 9'b111110110;
assign micromatrizz[52][296] = 9'b111110010;
assign micromatrizz[52][297] = 9'b111110011;
assign micromatrizz[52][298] = 9'b111110010;
assign micromatrizz[52][299] = 9'b111110010;
assign micromatrizz[52][300] = 9'b111110011;
assign micromatrizz[52][301] = 9'b111110010;
assign micromatrizz[52][302] = 9'b111110011;
assign micromatrizz[52][303] = 9'b111110011;
assign micromatrizz[52][304] = 9'b111111111;
assign micromatrizz[52][305] = 9'b111111111;
assign micromatrizz[52][306] = 9'b111111111;
assign micromatrizz[52][307] = 9'b111111111;
assign micromatrizz[52][308] = 9'b111111111;
assign micromatrizz[52][309] = 9'b111111111;
assign micromatrizz[52][310] = 9'b111111111;
assign micromatrizz[52][311] = 9'b111111111;
assign micromatrizz[52][312] = 9'b111111111;
assign micromatrizz[52][313] = 9'b111110111;
assign micromatrizz[52][314] = 9'b111110111;
assign micromatrizz[52][315] = 9'b111111111;
assign micromatrizz[52][316] = 9'b111111111;
assign micromatrizz[52][317] = 9'b111111111;
assign micromatrizz[52][318] = 9'b111111111;
assign micromatrizz[52][319] = 9'b111111111;
assign micromatrizz[52][320] = 9'b111111111;
assign micromatrizz[52][321] = 9'b111110111;
assign micromatrizz[52][322] = 9'b111110111;
assign micromatrizz[52][323] = 9'b111110111;
assign micromatrizz[52][324] = 9'b111110111;
assign micromatrizz[52][325] = 9'b111110111;
assign micromatrizz[52][326] = 9'b111110111;
assign micromatrizz[52][327] = 9'b111111111;
assign micromatrizz[52][328] = 9'b111111111;
assign micromatrizz[52][329] = 9'b111111111;
assign micromatrizz[52][330] = 9'b111111111;
assign micromatrizz[52][331] = 9'b111111111;
assign micromatrizz[52][332] = 9'b111111111;
assign micromatrizz[52][333] = 9'b111111111;
assign micromatrizz[52][334] = 9'b111111111;
assign micromatrizz[52][335] = 9'b111110010;
assign micromatrizz[52][336] = 9'b111110010;
assign micromatrizz[52][337] = 9'b111110011;
assign micromatrizz[52][338] = 9'b111110011;
assign micromatrizz[52][339] = 9'b111110011;
assign micromatrizz[52][340] = 9'b111110011;
assign micromatrizz[52][341] = 9'b111110011;
assign micromatrizz[52][342] = 9'b111110111;
assign micromatrizz[52][343] = 9'b111111111;
assign micromatrizz[52][344] = 9'b111111111;
assign micromatrizz[52][345] = 9'b111111111;
assign micromatrizz[52][346] = 9'b111110111;
assign micromatrizz[52][347] = 9'b111110011;
assign micromatrizz[52][348] = 9'b111110010;
assign micromatrizz[52][349] = 9'b111110010;
assign micromatrizz[52][350] = 9'b111110011;
assign micromatrizz[52][351] = 9'b111110111;
assign micromatrizz[52][352] = 9'b111111111;
assign micromatrizz[52][353] = 9'b111111111;
assign micromatrizz[52][354] = 9'b111111111;
assign micromatrizz[52][355] = 9'b111111111;
assign micromatrizz[52][356] = 9'b111111111;
assign micromatrizz[52][357] = 9'b111111111;
assign micromatrizz[52][358] = 9'b111110111;
assign micromatrizz[52][359] = 9'b111110010;
assign micromatrizz[52][360] = 9'b111110011;
assign micromatrizz[52][361] = 9'b111110010;
assign micromatrizz[52][362] = 9'b111110010;
assign micromatrizz[52][363] = 9'b111110010;
assign micromatrizz[52][364] = 9'b111110011;
assign micromatrizz[52][365] = 9'b111110011;
assign micromatrizz[52][366] = 9'b111110111;
assign micromatrizz[52][367] = 9'b111111111;
assign micromatrizz[52][368] = 9'b111110111;
assign micromatrizz[52][369] = 9'b111111111;
assign micromatrizz[52][370] = 9'b111111111;
assign micromatrizz[52][371] = 9'b111111111;
assign micromatrizz[52][372] = 9'b111110010;
assign micromatrizz[52][373] = 9'b111110010;
assign micromatrizz[52][374] = 9'b111110010;
assign micromatrizz[52][375] = 9'b111110011;
assign micromatrizz[52][376] = 9'b111110011;
assign micromatrizz[52][377] = 9'b111110011;
assign micromatrizz[52][378] = 9'b111110010;
assign micromatrizz[52][379] = 9'b111111111;
assign micromatrizz[52][380] = 9'b111111111;
assign micromatrizz[52][381] = 9'b111111111;
assign micromatrizz[52][382] = 9'b111111111;
assign micromatrizz[52][383] = 9'b111110111;
assign micromatrizz[52][384] = 9'b111110010;
assign micromatrizz[52][385] = 9'b111110010;
assign micromatrizz[52][386] = 9'b111110010;
assign micromatrizz[52][387] = 9'b111110011;
assign micromatrizz[52][388] = 9'b111110011;
assign micromatrizz[52][389] = 9'b111110011;
assign micromatrizz[52][390] = 9'b111110010;
assign micromatrizz[52][391] = 9'b111111111;
assign micromatrizz[52][392] = 9'b111111111;
assign micromatrizz[52][393] = 9'b111111111;
assign micromatrizz[52][394] = 9'b111111111;
assign micromatrizz[52][395] = 9'b111110111;
assign micromatrizz[52][396] = 9'b111110010;
assign micromatrizz[52][397] = 9'b111110010;
assign micromatrizz[52][398] = 9'b111110111;
assign micromatrizz[52][399] = 9'b111110010;
assign micromatrizz[52][400] = 9'b111110010;
assign micromatrizz[52][401] = 9'b111110011;
assign micromatrizz[52][402] = 9'b111110111;
assign micromatrizz[52][403] = 9'b111111111;
assign micromatrizz[52][404] = 9'b111111111;
assign micromatrizz[52][405] = 9'b111111111;
assign micromatrizz[52][406] = 9'b111110111;
assign micromatrizz[52][407] = 9'b111110010;
assign micromatrizz[52][408] = 9'b111110010;
assign micromatrizz[52][409] = 9'b111110111;
assign micromatrizz[52][410] = 9'b111111111;
assign micromatrizz[52][411] = 9'b111111111;
assign micromatrizz[52][412] = 9'b111111111;
assign micromatrizz[52][413] = 9'b111111111;
assign micromatrizz[52][414] = 9'b111111111;
assign micromatrizz[52][415] = 9'b111111111;
assign micromatrizz[52][416] = 9'b111111111;
assign micromatrizz[52][417] = 9'b111110111;
assign micromatrizz[52][418] = 9'b111110111;
assign micromatrizz[52][419] = 9'b111110111;
assign micromatrizz[52][420] = 9'b111110111;
assign micromatrizz[52][421] = 9'b111110111;
assign micromatrizz[52][422] = 9'b111111111;
assign micromatrizz[52][423] = 9'b111111111;
assign micromatrizz[52][424] = 9'b111111111;
assign micromatrizz[52][425] = 9'b111111111;
assign micromatrizz[52][426] = 9'b111111111;
assign micromatrizz[52][427] = 9'b111111111;
assign micromatrizz[52][428] = 9'b111111111;
assign micromatrizz[52][429] = 9'b111111111;
assign micromatrizz[52][430] = 9'b111110111;
assign micromatrizz[52][431] = 9'b111110010;
assign micromatrizz[52][432] = 9'b111110010;
assign micromatrizz[52][433] = 9'b111110010;
assign micromatrizz[52][434] = 9'b111110010;
assign micromatrizz[52][435] = 9'b111110011;
assign micromatrizz[52][436] = 9'b111110010;
assign micromatrizz[52][437] = 9'b111110111;
assign micromatrizz[52][438] = 9'b111111111;
assign micromatrizz[52][439] = 9'b111111111;
assign micromatrizz[52][440] = 9'b111111111;
assign micromatrizz[52][441] = 9'b111110111;
assign micromatrizz[52][442] = 9'b111110010;
assign micromatrizz[52][443] = 9'b111110010;
assign micromatrizz[52][444] = 9'b111110111;
assign micromatrizz[52][445] = 9'b111111111;
assign micromatrizz[52][446] = 9'b111111111;
assign micromatrizz[52][447] = 9'b111111111;
assign micromatrizz[52][448] = 9'b111111111;
assign micromatrizz[52][449] = 9'b111111111;
assign micromatrizz[52][450] = 9'b111111111;
assign micromatrizz[52][451] = 9'b111111111;
assign micromatrizz[52][452] = 9'b111110111;
assign micromatrizz[52][453] = 9'b111110111;
assign micromatrizz[52][454] = 9'b111110111;
assign micromatrizz[52][455] = 9'b111110111;
assign micromatrizz[52][456] = 9'b111110111;
assign micromatrizz[52][457] = 9'b111111111;
assign micromatrizz[52][458] = 9'b111111111;
assign micromatrizz[52][459] = 9'b111111111;
assign micromatrizz[52][460] = 9'b111111111;
assign micromatrizz[52][461] = 9'b111111111;
assign micromatrizz[52][462] = 9'b111111111;
assign micromatrizz[52][463] = 9'b111111111;
assign micromatrizz[52][464] = 9'b111111111;
assign micromatrizz[52][465] = 9'b111111111;
assign micromatrizz[52][466] = 9'b111111111;
assign micromatrizz[52][467] = 9'b111111111;
assign micromatrizz[52][468] = 9'b111111111;
assign micromatrizz[52][469] = 9'b111110111;
assign micromatrizz[52][470] = 9'b111110110;
assign micromatrizz[52][471] = 9'b111110111;
assign micromatrizz[52][472] = 9'b111110111;
assign micromatrizz[52][473] = 9'b111110111;
assign micromatrizz[52][474] = 9'b111110111;
assign micromatrizz[52][475] = 9'b111111111;
assign micromatrizz[52][476] = 9'b111111111;
assign micromatrizz[52][477] = 9'b111111111;
assign micromatrizz[52][478] = 9'b111111111;
assign micromatrizz[52][479] = 9'b111111111;
assign micromatrizz[52][480] = 9'b111111111;
assign micromatrizz[52][481] = 9'b111110110;
assign micromatrizz[52][482] = 9'b111110010;
assign micromatrizz[52][483] = 9'b111110010;
assign micromatrizz[52][484] = 9'b111110010;
assign micromatrizz[52][485] = 9'b111110010;
assign micromatrizz[52][486] = 9'b111110010;
assign micromatrizz[52][487] = 9'b111110011;
assign micromatrizz[52][488] = 9'b111110111;
assign micromatrizz[52][489] = 9'b111111111;
assign micromatrizz[52][490] = 9'b111111111;
assign micromatrizz[52][491] = 9'b111111111;
assign micromatrizz[52][492] = 9'b111110111;
assign micromatrizz[52][493] = 9'b111110010;
assign micromatrizz[52][494] = 9'b111110010;
assign micromatrizz[52][495] = 9'b111111111;
assign micromatrizz[52][496] = 9'b111111111;
assign micromatrizz[52][497] = 9'b111111111;
assign micromatrizz[52][498] = 9'b111111111;
assign micromatrizz[52][499] = 9'b111111111;
assign micromatrizz[52][500] = 9'b111111111;
assign micromatrizz[52][501] = 9'b111111111;
assign micromatrizz[52][502] = 9'b111110111;
assign micromatrizz[52][503] = 9'b111110011;
assign micromatrizz[52][504] = 9'b111110111;
assign micromatrizz[52][505] = 9'b111110111;
assign micromatrizz[52][506] = 9'b111110111;
assign micromatrizz[52][507] = 9'b111110111;
assign micromatrizz[52][508] = 9'b111111111;
assign micromatrizz[52][509] = 9'b111111111;
assign micromatrizz[52][510] = 9'b111111111;
assign micromatrizz[52][511] = 9'b111111111;
assign micromatrizz[52][512] = 9'b111111111;
assign micromatrizz[52][513] = 9'b111111111;
assign micromatrizz[52][514] = 9'b111111111;
assign micromatrizz[52][515] = 9'b111111111;
assign micromatrizz[52][516] = 9'b111110111;
assign micromatrizz[52][517] = 9'b111110011;
assign micromatrizz[52][518] = 9'b111110011;
assign micromatrizz[52][519] = 9'b111110011;
assign micromatrizz[52][520] = 9'b111110010;
assign micromatrizz[52][521] = 9'b111110010;
assign micromatrizz[52][522] = 9'b111110011;
assign micromatrizz[52][523] = 9'b111110111;
assign micromatrizz[52][524] = 9'b111111111;
assign micromatrizz[52][525] = 9'b111111111;
assign micromatrizz[52][526] = 9'b111110111;
assign micromatrizz[52][527] = 9'b111110010;
assign micromatrizz[52][528] = 9'b111110010;
assign micromatrizz[52][529] = 9'b111110010;
assign micromatrizz[52][530] = 9'b111110111;
assign micromatrizz[52][531] = 9'b111111111;
assign micromatrizz[52][532] = 9'b111111111;
assign micromatrizz[52][533] = 9'b111111111;
assign micromatrizz[52][534] = 9'b111111111;
assign micromatrizz[52][535] = 9'b111111111;
assign micromatrizz[52][536] = 9'b111111111;
assign micromatrizz[52][537] = 9'b111111111;
assign micromatrizz[52][538] = 9'b111111111;
assign micromatrizz[52][539] = 9'b111111111;
assign micromatrizz[52][540] = 9'b111111111;
assign micromatrizz[52][541] = 9'b111111111;
assign micromatrizz[52][542] = 9'b111111111;
assign micromatrizz[52][543] = 9'b111111111;
assign micromatrizz[52][544] = 9'b111110111;
assign micromatrizz[52][545] = 9'b111110011;
assign micromatrizz[52][546] = 9'b111110111;
assign micromatrizz[52][547] = 9'b111110111;
assign micromatrizz[52][548] = 9'b111110111;
assign micromatrizz[52][549] = 9'b111110111;
assign micromatrizz[52][550] = 9'b111111111;
assign micromatrizz[52][551] = 9'b111111111;
assign micromatrizz[52][552] = 9'b111111111;
assign micromatrizz[52][553] = 9'b111111111;
assign micromatrizz[52][554] = 9'b111111111;
assign micromatrizz[52][555] = 9'b111111111;
assign micromatrizz[52][556] = 9'b111111111;
assign micromatrizz[52][557] = 9'b111111111;
assign micromatrizz[52][558] = 9'b111110010;
assign micromatrizz[52][559] = 9'b111110010;
assign micromatrizz[52][560] = 9'b111110010;
assign micromatrizz[52][561] = 9'b111110010;
assign micromatrizz[52][562] = 9'b111110011;
assign micromatrizz[52][563] = 9'b111110011;
assign micromatrizz[52][564] = 9'b111110011;
assign micromatrizz[52][565] = 9'b111111111;
assign micromatrizz[52][566] = 9'b111111111;
assign micromatrizz[52][567] = 9'b111111111;
assign micromatrizz[52][568] = 9'b111111111;
assign micromatrizz[52][569] = 9'b111111111;
assign micromatrizz[52][570] = 9'b111111111;
assign micromatrizz[52][571] = 9'b111111111;
assign micromatrizz[52][572] = 9'b111111111;
assign micromatrizz[52][573] = 9'b111110111;
assign micromatrizz[52][574] = 9'b111110010;
assign micromatrizz[52][575] = 9'b111110011;
assign micromatrizz[52][576] = 9'b111110010;
assign micromatrizz[52][577] = 9'b111110111;
assign micromatrizz[52][578] = 9'b111111111;
assign micromatrizz[52][579] = 9'b111111111;
assign micromatrizz[52][580] = 9'b111111111;
assign micromatrizz[52][581] = 9'b111110010;
assign micromatrizz[52][582] = 9'b111110011;
assign micromatrizz[52][583] = 9'b111110011;
assign micromatrizz[52][584] = 9'b111110010;
assign micromatrizz[52][585] = 9'b111110010;
assign micromatrizz[52][586] = 9'b111110011;
assign micromatrizz[52][587] = 9'b111110011;
assign micromatrizz[52][588] = 9'b111111111;
assign micromatrizz[52][589] = 9'b111111111;
assign micromatrizz[52][590] = 9'b111111111;
assign micromatrizz[52][591] = 9'b111111111;
assign micromatrizz[52][592] = 9'b111111111;
assign micromatrizz[52][593] = 9'b111111111;
assign micromatrizz[52][594] = 9'b111111111;
assign micromatrizz[52][595] = 9'b111111111;
assign micromatrizz[52][596] = 9'b111111111;
assign micromatrizz[52][597] = 9'b111110111;
assign micromatrizz[52][598] = 9'b111110111;
assign micromatrizz[52][599] = 9'b111110111;
assign micromatrizz[52][600] = 9'b111110111;
assign micromatrizz[52][601] = 9'b111110111;
assign micromatrizz[52][602] = 9'b111111111;
assign micromatrizz[52][603] = 9'b111111111;
assign micromatrizz[52][604] = 9'b111111111;
assign micromatrizz[52][605] = 9'b111111111;
assign micromatrizz[52][606] = 9'b111111111;
assign micromatrizz[52][607] = 9'b111111111;
assign micromatrizz[52][608] = 9'b111111111;
assign micromatrizz[52][609] = 9'b111111111;
assign micromatrizz[52][610] = 9'b111111111;
assign micromatrizz[52][611] = 9'b111111111;
assign micromatrizz[52][612] = 9'b111111111;
assign micromatrizz[52][613] = 9'b111111111;
assign micromatrizz[52][614] = 9'b111110111;
assign micromatrizz[52][615] = 9'b111110011;
assign micromatrizz[52][616] = 9'b111110111;
assign micromatrizz[52][617] = 9'b111110111;
assign micromatrizz[52][618] = 9'b111110111;
assign micromatrizz[52][619] = 9'b111110111;
assign micromatrizz[52][620] = 9'b111111111;
assign micromatrizz[52][621] = 9'b111111111;
assign micromatrizz[52][622] = 9'b111111111;
assign micromatrizz[52][623] = 9'b111111111;
assign micromatrizz[52][624] = 9'b111111111;
assign micromatrizz[52][625] = 9'b111111111;
assign micromatrizz[52][626] = 9'b111111111;
assign micromatrizz[52][627] = 9'b111111111;
assign micromatrizz[52][628] = 9'b111111111;
assign micromatrizz[52][629] = 9'b111111111;
assign micromatrizz[52][630] = 9'b111111111;
assign micromatrizz[52][631] = 9'b111111111;
assign micromatrizz[52][632] = 9'b111111111;
assign micromatrizz[52][633] = 9'b111111111;
assign micromatrizz[52][634] = 9'b111111111;
assign micromatrizz[52][635] = 9'b111111111;
assign micromatrizz[52][636] = 9'b111111111;
assign micromatrizz[52][637] = 9'b111111111;
assign micromatrizz[52][638] = 9'b111111111;
assign micromatrizz[52][639] = 9'b111111111;
assign micromatrizz[53][0] = 9'b111111111;
assign micromatrizz[53][1] = 9'b111111111;
assign micromatrizz[53][2] = 9'b111111111;
assign micromatrizz[53][3] = 9'b111111111;
assign micromatrizz[53][4] = 9'b111111111;
assign micromatrizz[53][5] = 9'b111111111;
assign micromatrizz[53][6] = 9'b111111111;
assign micromatrizz[53][7] = 9'b111111111;
assign micromatrizz[53][8] = 9'b111111111;
assign micromatrizz[53][9] = 9'b111111111;
assign micromatrizz[53][10] = 9'b111110010;
assign micromatrizz[53][11] = 9'b111110010;
assign micromatrizz[53][12] = 9'b111110010;
assign micromatrizz[53][13] = 9'b111110111;
assign micromatrizz[53][14] = 9'b111111111;
assign micromatrizz[53][15] = 9'b111111111;
assign micromatrizz[53][16] = 9'b111111111;
assign micromatrizz[53][17] = 9'b111110111;
assign micromatrizz[53][18] = 9'b111110010;
assign micromatrizz[53][19] = 9'b111110111;
assign micromatrizz[53][20] = 9'b111111111;
assign micromatrizz[53][21] = 9'b111111111;
assign micromatrizz[53][22] = 9'b111111111;
assign micromatrizz[53][23] = 9'b111110111;
assign micromatrizz[53][24] = 9'b111110010;
assign micromatrizz[53][25] = 9'b111110010;
assign micromatrizz[53][26] = 9'b111110010;
assign micromatrizz[53][27] = 9'b111110011;
assign micromatrizz[53][28] = 9'b111110011;
assign micromatrizz[53][29] = 9'b111110011;
assign micromatrizz[53][30] = 9'b111110011;
assign micromatrizz[53][31] = 9'b111111111;
assign micromatrizz[53][32] = 9'b111111111;
assign micromatrizz[53][33] = 9'b111111111;
assign micromatrizz[53][34] = 9'b111111111;
assign micromatrizz[53][35] = 9'b111110111;
assign micromatrizz[53][36] = 9'b111110010;
assign micromatrizz[53][37] = 9'b111110010;
assign micromatrizz[53][38] = 9'b111110010;
assign micromatrizz[53][39] = 9'b111110010;
assign micromatrizz[53][40] = 9'b111110011;
assign micromatrizz[53][41] = 9'b111110011;
assign micromatrizz[53][42] = 9'b111110011;
assign micromatrizz[53][43] = 9'b111111111;
assign micromatrizz[53][44] = 9'b111111111;
assign micromatrizz[53][45] = 9'b111111111;
assign micromatrizz[53][46] = 9'b111111111;
assign micromatrizz[53][47] = 9'b111110010;
assign micromatrizz[53][48] = 9'b111110010;
assign micromatrizz[53][49] = 9'b111110010;
assign micromatrizz[53][50] = 9'b111110010;
assign micromatrizz[53][51] = 9'b111110010;
assign micromatrizz[53][52] = 9'b111110011;
assign micromatrizz[53][53] = 9'b111110010;
assign micromatrizz[53][54] = 9'b111110111;
assign micromatrizz[53][55] = 9'b111111111;
assign micromatrizz[53][56] = 9'b111110111;
assign micromatrizz[53][57] = 9'b111110111;
assign micromatrizz[53][58] = 9'b111110011;
assign micromatrizz[53][59] = 9'b111110010;
assign micromatrizz[53][60] = 9'b111110011;
assign micromatrizz[53][61] = 9'b111110010;
assign micromatrizz[53][62] = 9'b111110010;
assign micromatrizz[53][63] = 9'b111110111;
assign micromatrizz[53][64] = 9'b111111111;
assign micromatrizz[53][65] = 9'b111111111;
assign micromatrizz[53][66] = 9'b111111111;
assign micromatrizz[53][67] = 9'b111111111;
assign micromatrizz[53][68] = 9'b111111111;
assign micromatrizz[53][69] = 9'b111111111;
assign micromatrizz[53][70] = 9'b111111111;
assign micromatrizz[53][71] = 9'b111111111;
assign micromatrizz[53][72] = 9'b111110111;
assign micromatrizz[53][73] = 9'b111110010;
assign micromatrizz[53][74] = 9'b111110010;
assign micromatrizz[53][75] = 9'b111110111;
assign micromatrizz[53][76] = 9'b111111111;
assign micromatrizz[53][77] = 9'b111111111;
assign micromatrizz[53][78] = 9'b111111111;
assign micromatrizz[53][79] = 9'b111110010;
assign micromatrizz[53][80] = 9'b111110010;
assign micromatrizz[53][81] = 9'b111111111;
assign micromatrizz[53][82] = 9'b111111111;
assign micromatrizz[53][83] = 9'b111111111;
assign micromatrizz[53][84] = 9'b111111111;
assign micromatrizz[53][85] = 9'b111111111;
assign micromatrizz[53][86] = 9'b111111111;
assign micromatrizz[53][87] = 9'b111111111;
assign micromatrizz[53][88] = 9'b111110010;
assign micromatrizz[53][89] = 9'b111110010;
assign micromatrizz[53][90] = 9'b111110010;
assign micromatrizz[53][91] = 9'b111110011;
assign micromatrizz[53][92] = 9'b111110010;
assign micromatrizz[53][93] = 9'b111110010;
assign micromatrizz[53][94] = 9'b111110011;
assign micromatrizz[53][95] = 9'b111110111;
assign micromatrizz[53][96] = 9'b111111111;
assign micromatrizz[53][97] = 9'b111110111;
assign micromatrizz[53][98] = 9'b111110111;
assign micromatrizz[53][99] = 9'b111110111;
assign micromatrizz[53][100] = 9'b111110111;
assign micromatrizz[53][101] = 9'b111110010;
assign micromatrizz[53][102] = 9'b111110110;
assign micromatrizz[53][103] = 9'b111111111;
assign micromatrizz[53][104] = 9'b111111111;
assign micromatrizz[53][105] = 9'b111111111;
assign micromatrizz[53][106] = 9'b111110111;
assign micromatrizz[53][107] = 9'b111110010;
assign micromatrizz[53][108] = 9'b111110010;
assign micromatrizz[53][109] = 9'b111110111;
assign micromatrizz[53][110] = 9'b111111111;
assign micromatrizz[53][111] = 9'b111111111;
assign micromatrizz[53][112] = 9'b111111111;
assign micromatrizz[53][113] = 9'b111111111;
assign micromatrizz[53][114] = 9'b111110111;
assign micromatrizz[53][115] = 9'b111110110;
assign micromatrizz[53][116] = 9'b111111111;
assign micromatrizz[53][117] = 9'b111111111;
assign micromatrizz[53][118] = 9'b111111111;
assign micromatrizz[53][119] = 9'b111111111;
assign micromatrizz[53][120] = 9'b111111111;
assign micromatrizz[53][121] = 9'b111111111;
assign micromatrizz[53][122] = 9'b111111111;
assign micromatrizz[53][123] = 9'b111110010;
assign micromatrizz[53][124] = 9'b111110010;
assign micromatrizz[53][125] = 9'b111110011;
assign micromatrizz[53][126] = 9'b111110011;
assign micromatrizz[53][127] = 9'b111111111;
assign micromatrizz[53][128] = 9'b111111111;
assign micromatrizz[53][129] = 9'b111111111;
assign micromatrizz[53][130] = 9'b111110111;
assign micromatrizz[53][131] = 9'b111110111;
assign micromatrizz[53][132] = 9'b111111111;
assign micromatrizz[53][133] = 9'b111111111;
assign micromatrizz[53][134] = 9'b111111111;
assign micromatrizz[53][135] = 9'b111111111;
assign micromatrizz[53][136] = 9'b111111111;
assign micromatrizz[53][137] = 9'b111111111;
assign micromatrizz[53][138] = 9'b111110111;
assign micromatrizz[53][139] = 9'b111110010;
assign micromatrizz[53][140] = 9'b111110010;
assign micromatrizz[53][141] = 9'b111110010;
assign micromatrizz[53][142] = 9'b111110011;
assign micromatrizz[53][143] = 9'b111110011;
assign micromatrizz[53][144] = 9'b111110011;
assign micromatrizz[53][145] = 9'b111110011;
assign micromatrizz[53][146] = 9'b111110111;
assign micromatrizz[53][147] = 9'b111110110;
assign micromatrizz[53][148] = 9'b111110111;
assign micromatrizz[53][149] = 9'b111110111;
assign micromatrizz[53][150] = 9'b111110010;
assign micromatrizz[53][151] = 9'b111110010;
assign micromatrizz[53][152] = 9'b111110010;
assign micromatrizz[53][153] = 9'b111110011;
assign micromatrizz[53][154] = 9'b111110011;
assign micromatrizz[53][155] = 9'b111110010;
assign micromatrizz[53][156] = 9'b111110111;
assign micromatrizz[53][157] = 9'b111111111;
assign micromatrizz[53][158] = 9'b111111111;
assign micromatrizz[53][159] = 9'b111111111;
assign micromatrizz[53][160] = 9'b111111111;
assign micromatrizz[53][161] = 9'b111111111;
assign micromatrizz[53][162] = 9'b111111111;
assign micromatrizz[53][163] = 9'b111111111;
assign micromatrizz[53][164] = 9'b111110111;
assign micromatrizz[53][165] = 9'b111110110;
assign micromatrizz[53][166] = 9'b111111111;
assign micromatrizz[53][167] = 9'b111111111;
assign micromatrizz[53][168] = 9'b111111111;
assign micromatrizz[53][169] = 9'b111111111;
assign micromatrizz[53][170] = 9'b111111111;
assign micromatrizz[53][171] = 9'b111110111;
assign micromatrizz[53][172] = 9'b111110010;
assign micromatrizz[53][173] = 9'b111110010;
assign micromatrizz[53][174] = 9'b111110011;
assign micromatrizz[53][175] = 9'b111110010;
assign micromatrizz[53][176] = 9'b111110010;
assign micromatrizz[53][177] = 9'b111110111;
assign micromatrizz[53][178] = 9'b111111111;
assign micromatrizz[53][179] = 9'b111111111;
assign micromatrizz[53][180] = 9'b111111111;
assign micromatrizz[53][181] = 9'b111111111;
assign micromatrizz[53][182] = 9'b111111111;
assign micromatrizz[53][183] = 9'b111111111;
assign micromatrizz[53][184] = 9'b111111111;
assign micromatrizz[53][185] = 9'b111111111;
assign micromatrizz[53][186] = 9'b111110110;
assign micromatrizz[53][187] = 9'b111110010;
assign micromatrizz[53][188] = 9'b111110010;
assign micromatrizz[53][189] = 9'b111110011;
assign micromatrizz[53][190] = 9'b111110011;
assign micromatrizz[53][191] = 9'b111110111;
assign micromatrizz[53][192] = 9'b111110111;
assign micromatrizz[53][193] = 9'b111110111;
assign micromatrizz[53][194] = 9'b111111111;
assign micromatrizz[53][195] = 9'b111110010;
assign micromatrizz[53][196] = 9'b111110010;
assign micromatrizz[53][197] = 9'b111110011;
assign micromatrizz[53][198] = 9'b111110011;
assign micromatrizz[53][199] = 9'b111110010;
assign micromatrizz[53][200] = 9'b111110010;
assign micromatrizz[53][201] = 9'b111110011;
assign micromatrizz[53][202] = 9'b111110111;
assign micromatrizz[53][203] = 9'b111111111;
assign micromatrizz[53][204] = 9'b111111111;
assign micromatrizz[53][205] = 9'b111111111;
assign micromatrizz[53][206] = 9'b111111111;
assign micromatrizz[53][207] = 9'b111111111;
assign micromatrizz[53][208] = 9'b111111111;
assign micromatrizz[53][209] = 9'b111110111;
assign micromatrizz[53][210] = 9'b111110011;
assign micromatrizz[53][211] = 9'b111110011;
assign micromatrizz[53][212] = 9'b111110011;
assign micromatrizz[53][213] = 9'b111110111;
assign micromatrizz[53][214] = 9'b111111111;
assign micromatrizz[53][215] = 9'b111111111;
assign micromatrizz[53][216] = 9'b111111111;
assign micromatrizz[53][217] = 9'b111110111;
assign micromatrizz[53][218] = 9'b111110111;
assign micromatrizz[53][219] = 9'b111111111;
assign micromatrizz[53][220] = 9'b111111111;
assign micromatrizz[53][221] = 9'b111111111;
assign micromatrizz[53][222] = 9'b111111111;
assign micromatrizz[53][223] = 9'b111111111;
assign micromatrizz[53][224] = 9'b111111111;
assign micromatrizz[53][225] = 9'b111110111;
assign micromatrizz[53][226] = 9'b111110010;
assign micromatrizz[53][227] = 9'b111110010;
assign micromatrizz[53][228] = 9'b111110010;
assign micromatrizz[53][229] = 9'b111110010;
assign micromatrizz[53][230] = 9'b111110011;
assign micromatrizz[53][231] = 9'b111110010;
assign micromatrizz[53][232] = 9'b111110111;
assign micromatrizz[53][233] = 9'b111111111;
assign micromatrizz[53][234] = 9'b111111111;
assign micromatrizz[53][235] = 9'b111110111;
assign micromatrizz[53][236] = 9'b111110111;
assign micromatrizz[53][237] = 9'b111110111;
assign micromatrizz[53][238] = 9'b111110010;
assign micromatrizz[53][239] = 9'b111110010;
assign micromatrizz[53][240] = 9'b111111111;
assign micromatrizz[53][241] = 9'b111111111;
assign micromatrizz[53][242] = 9'b111111111;
assign micromatrizz[53][243] = 9'b111111111;
assign micromatrizz[53][244] = 9'b111111111;
assign micromatrizz[53][245] = 9'b111110011;
assign micromatrizz[53][246] = 9'b111110010;
assign micromatrizz[53][247] = 9'b111110011;
assign micromatrizz[53][248] = 9'b111111111;
assign micromatrizz[53][249] = 9'b111111111;
assign micromatrizz[53][250] = 9'b111111111;
assign micromatrizz[53][251] = 9'b111110010;
assign micromatrizz[53][252] = 9'b111110010;
assign micromatrizz[53][253] = 9'b111110111;
assign micromatrizz[53][254] = 9'b111111111;
assign micromatrizz[53][255] = 9'b111111111;
assign micromatrizz[53][256] = 9'b111111111;
assign micromatrizz[53][257] = 9'b111111111;
assign micromatrizz[53][258] = 9'b111111111;
assign micromatrizz[53][259] = 9'b111111111;
assign micromatrizz[53][260] = 9'b111111111;
assign micromatrizz[53][261] = 9'b111110111;
assign micromatrizz[53][262] = 9'b111110010;
assign micromatrizz[53][263] = 9'b111110010;
assign micromatrizz[53][264] = 9'b111110010;
assign micromatrizz[53][265] = 9'b111111111;
assign micromatrizz[53][266] = 9'b111111111;
assign micromatrizz[53][267] = 9'b111111111;
assign micromatrizz[53][268] = 9'b111111111;
assign micromatrizz[53][269] = 9'b111110111;
assign micromatrizz[53][270] = 9'b111110110;
assign micromatrizz[53][271] = 9'b111111111;
assign micromatrizz[53][272] = 9'b111111111;
assign micromatrizz[53][273] = 9'b111111111;
assign micromatrizz[53][274] = 9'b111111111;
assign micromatrizz[53][275] = 9'b111111111;
assign micromatrizz[53][276] = 9'b111111111;
assign micromatrizz[53][277] = 9'b111111111;
assign micromatrizz[53][278] = 9'b111110111;
assign micromatrizz[53][279] = 9'b111110110;
assign micromatrizz[53][280] = 9'b111111111;
assign micromatrizz[53][281] = 9'b111111111;
assign micromatrizz[53][282] = 9'b111111111;
assign micromatrizz[53][283] = 9'b111111111;
assign micromatrizz[53][284] = 9'b111111111;
assign micromatrizz[53][285] = 9'b111110111;
assign micromatrizz[53][286] = 9'b111110010;
assign micromatrizz[53][287] = 9'b111110010;
assign micromatrizz[53][288] = 9'b111110011;
assign micromatrizz[53][289] = 9'b111110010;
assign micromatrizz[53][290] = 9'b111110010;
assign micromatrizz[53][291] = 9'b111110111;
assign micromatrizz[53][292] = 9'b111111111;
assign micromatrizz[53][293] = 9'b111111111;
assign micromatrizz[53][294] = 9'b111111111;
assign micromatrizz[53][295] = 9'b111111111;
assign micromatrizz[53][296] = 9'b111110010;
assign micromatrizz[53][297] = 9'b111110010;
assign micromatrizz[53][298] = 9'b111110010;
assign micromatrizz[53][299] = 9'b111110010;
assign micromatrizz[53][300] = 9'b111110010;
assign micromatrizz[53][301] = 9'b111110010;
assign micromatrizz[53][302] = 9'b111110011;
assign micromatrizz[53][303] = 9'b111110010;
assign micromatrizz[53][304] = 9'b111110111;
assign micromatrizz[53][305] = 9'b111111111;
assign micromatrizz[53][306] = 9'b111111111;
assign micromatrizz[53][307] = 9'b111111111;
assign micromatrizz[53][308] = 9'b111111111;
assign micromatrizz[53][309] = 9'b111111111;
assign micromatrizz[53][310] = 9'b111111111;
assign micromatrizz[53][311] = 9'b111111111;
assign micromatrizz[53][312] = 9'b111111111;
assign micromatrizz[53][313] = 9'b111110010;
assign micromatrizz[53][314] = 9'b111111111;
assign micromatrizz[53][315] = 9'b111111111;
assign micromatrizz[53][316] = 9'b111111111;
assign micromatrizz[53][317] = 9'b111111111;
assign micromatrizz[53][318] = 9'b111111111;
assign micromatrizz[53][319] = 9'b111110111;
assign micromatrizz[53][320] = 9'b111110010;
assign micromatrizz[53][321] = 9'b111110011;
assign micromatrizz[53][322] = 9'b111110111;
assign micromatrizz[53][323] = 9'b111111111;
assign micromatrizz[53][324] = 9'b111111111;
assign micromatrizz[53][325] = 9'b111111111;
assign micromatrizz[53][326] = 9'b111110010;
assign micromatrizz[53][327] = 9'b111110010;
assign micromatrizz[53][328] = 9'b111111111;
assign micromatrizz[53][329] = 9'b111111111;
assign micromatrizz[53][330] = 9'b111111111;
assign micromatrizz[53][331] = 9'b111111111;
assign micromatrizz[53][332] = 9'b111111111;
assign micromatrizz[53][333] = 9'b111111111;
assign micromatrizz[53][334] = 9'b111111111;
assign micromatrizz[53][335] = 9'b111110010;
assign micromatrizz[53][336] = 9'b111110010;
assign micromatrizz[53][337] = 9'b111110011;
assign micromatrizz[53][338] = 9'b111110011;
assign micromatrizz[53][339] = 9'b111110011;
assign micromatrizz[53][340] = 9'b111110011;
assign micromatrizz[53][341] = 9'b111110010;
assign micromatrizz[53][342] = 9'b111110011;
assign micromatrizz[53][343] = 9'b111110111;
assign micromatrizz[53][344] = 9'b111110111;
assign micromatrizz[53][345] = 9'b111110111;
assign micromatrizz[53][346] = 9'b111110111;
assign micromatrizz[53][347] = 9'b111110010;
assign micromatrizz[53][348] = 9'b111110010;
assign micromatrizz[53][349] = 9'b111110011;
assign micromatrizz[53][350] = 9'b111110011;
assign micromatrizz[53][351] = 9'b111110011;
assign micromatrizz[53][352] = 9'b111110111;
assign micromatrizz[53][353] = 9'b111111111;
assign micromatrizz[53][354] = 9'b111111111;
assign micromatrizz[53][355] = 9'b111111111;
assign micromatrizz[53][356] = 9'b111111111;
assign micromatrizz[53][357] = 9'b111111111;
assign micromatrizz[53][358] = 9'b111111111;
assign micromatrizz[53][359] = 9'b111110010;
assign micromatrizz[53][360] = 9'b111110011;
assign micromatrizz[53][361] = 9'b111110010;
assign micromatrizz[53][362] = 9'b111110010;
assign micromatrizz[53][363] = 9'b111110010;
assign micromatrizz[53][364] = 9'b111110011;
assign micromatrizz[53][365] = 9'b111110011;
assign micromatrizz[53][366] = 9'b111111111;
assign micromatrizz[53][367] = 9'b111111111;
assign micromatrizz[53][368] = 9'b111111111;
assign micromatrizz[53][369] = 9'b111111111;
assign micromatrizz[53][370] = 9'b111111111;
assign micromatrizz[53][371] = 9'b111111111;
assign micromatrizz[53][372] = 9'b111110010;
assign micromatrizz[53][373] = 9'b111110010;
assign micromatrizz[53][374] = 9'b111110010;
assign micromatrizz[53][375] = 9'b111110011;
assign micromatrizz[53][376] = 9'b111110011;
assign micromatrizz[53][377] = 9'b111110011;
assign micromatrizz[53][378] = 9'b111110010;
assign micromatrizz[53][379] = 9'b111111111;
assign micromatrizz[53][380] = 9'b111111111;
assign micromatrizz[53][381] = 9'b111111111;
assign micromatrizz[53][382] = 9'b111111111;
assign micromatrizz[53][383] = 9'b111110111;
assign micromatrizz[53][384] = 9'b111110010;
assign micromatrizz[53][385] = 9'b111110011;
assign micromatrizz[53][386] = 9'b111110010;
assign micromatrizz[53][387] = 9'b111110011;
assign micromatrizz[53][388] = 9'b111110011;
assign micromatrizz[53][389] = 9'b111110011;
assign micromatrizz[53][390] = 9'b111110010;
assign micromatrizz[53][391] = 9'b111111111;
assign micromatrizz[53][392] = 9'b111111111;
assign micromatrizz[53][393] = 9'b111111111;
assign micromatrizz[53][394] = 9'b111111111;
assign micromatrizz[53][395] = 9'b111110111;
assign micromatrizz[53][396] = 9'b111110010;
assign micromatrizz[53][397] = 9'b111110010;
assign micromatrizz[53][398] = 9'b111110010;
assign micromatrizz[53][399] = 9'b111110011;
assign micromatrizz[53][400] = 9'b111110011;
assign micromatrizz[53][401] = 9'b111110010;
assign micromatrizz[53][402] = 9'b111110111;
assign micromatrizz[53][403] = 9'b111111111;
assign micromatrizz[53][404] = 9'b111110111;
assign micromatrizz[53][405] = 9'b111110111;
assign micromatrizz[53][406] = 9'b111110111;
assign micromatrizz[53][407] = 9'b111110111;
assign micromatrizz[53][408] = 9'b111110010;
assign micromatrizz[53][409] = 9'b111110010;
assign micromatrizz[53][410] = 9'b111111111;
assign micromatrizz[53][411] = 9'b111111111;
assign micromatrizz[53][412] = 9'b111111111;
assign micromatrizz[53][413] = 9'b111111111;
assign micromatrizz[53][414] = 9'b111111111;
assign micromatrizz[53][415] = 9'b111110010;
assign micromatrizz[53][416] = 9'b111110010;
assign micromatrizz[53][417] = 9'b111110010;
assign micromatrizz[53][418] = 9'b111111111;
assign micromatrizz[53][419] = 9'b111111111;
assign micromatrizz[53][420] = 9'b111111111;
assign micromatrizz[53][421] = 9'b111110010;
assign micromatrizz[53][422] = 9'b111110010;
assign micromatrizz[53][423] = 9'b111110111;
assign micromatrizz[53][424] = 9'b111111111;
assign micromatrizz[53][425] = 9'b111111111;
assign micromatrizz[53][426] = 9'b111111111;
assign micromatrizz[53][427] = 9'b111111111;
assign micromatrizz[53][428] = 9'b111111111;
assign micromatrizz[53][429] = 9'b111111111;
assign micromatrizz[53][430] = 9'b111110111;
assign micromatrizz[53][431] = 9'b111110010;
assign micromatrizz[53][432] = 9'b111110010;
assign micromatrizz[53][433] = 9'b111110010;
assign micromatrizz[53][434] = 9'b111110010;
assign micromatrizz[53][435] = 9'b111110010;
assign micromatrizz[53][436] = 9'b111110011;
assign micromatrizz[53][437] = 9'b111110011;
assign micromatrizz[53][438] = 9'b111111111;
assign micromatrizz[53][439] = 9'b111111111;
assign micromatrizz[53][440] = 9'b111110111;
assign micromatrizz[53][441] = 9'b111110111;
assign micromatrizz[53][442] = 9'b111110111;
assign micromatrizz[53][443] = 9'b111110011;
assign micromatrizz[53][444] = 9'b111110010;
assign micromatrizz[53][445] = 9'b111111111;
assign micromatrizz[53][446] = 9'b111111111;
assign micromatrizz[53][447] = 9'b111111111;
assign micromatrizz[53][448] = 9'b111111111;
assign micromatrizz[53][449] = 9'b111111111;
assign micromatrizz[53][450] = 9'b111110111;
assign micromatrizz[53][451] = 9'b111110010;
assign micromatrizz[53][452] = 9'b111110011;
assign micromatrizz[53][453] = 9'b111110011;
assign micromatrizz[53][454] = 9'b111111111;
assign micromatrizz[53][455] = 9'b111111111;
assign micromatrizz[53][456] = 9'b111111111;
assign micromatrizz[53][457] = 9'b111110111;
assign micromatrizz[53][458] = 9'b111110111;
assign micromatrizz[53][459] = 9'b111111111;
assign micromatrizz[53][460] = 9'b111111111;
assign micromatrizz[53][461] = 9'b111111111;
assign micromatrizz[53][462] = 9'b111111111;
assign micromatrizz[53][463] = 9'b111111111;
assign micromatrizz[53][464] = 9'b111111111;
assign micromatrizz[53][465] = 9'b111111111;
assign micromatrizz[53][466] = 9'b111111111;
assign micromatrizz[53][467] = 9'b111110011;
assign micromatrizz[53][468] = 9'b111110010;
assign micromatrizz[53][469] = 9'b111110010;
assign micromatrizz[53][470] = 9'b111110111;
assign micromatrizz[53][471] = 9'b111111111;
assign micromatrizz[53][472] = 9'b111111111;
assign micromatrizz[53][473] = 9'b111111111;
assign micromatrizz[53][474] = 9'b111111111;
assign micromatrizz[53][475] = 9'b111110110;
assign micromatrizz[53][476] = 9'b111110111;
assign micromatrizz[53][477] = 9'b111111111;
assign micromatrizz[53][478] = 9'b111111111;
assign micromatrizz[53][479] = 9'b111111111;
assign micromatrizz[53][480] = 9'b111111111;
assign micromatrizz[53][481] = 9'b111110010;
assign micromatrizz[53][482] = 9'b111110010;
assign micromatrizz[53][483] = 9'b111110010;
assign micromatrizz[53][484] = 9'b111110010;
assign micromatrizz[53][485] = 9'b111110010;
assign micromatrizz[53][486] = 9'b111110010;
assign micromatrizz[53][487] = 9'b111110010;
assign micromatrizz[53][488] = 9'b111110111;
assign micromatrizz[53][489] = 9'b111111111;
assign micromatrizz[53][490] = 9'b111110111;
assign micromatrizz[53][491] = 9'b111110111;
assign micromatrizz[53][492] = 9'b111110111;
assign micromatrizz[53][493] = 9'b111110111;
assign micromatrizz[53][494] = 9'b111110010;
assign micromatrizz[53][495] = 9'b111110110;
assign micromatrizz[53][496] = 9'b111111111;
assign micromatrizz[53][497] = 9'b111111111;
assign micromatrizz[53][498] = 9'b111111111;
assign micromatrizz[53][499] = 9'b111111111;
assign micromatrizz[53][500] = 9'b111110111;
assign micromatrizz[53][501] = 9'b111110011;
assign micromatrizz[53][502] = 9'b111110010;
assign micromatrizz[53][503] = 9'b111110010;
assign micromatrizz[53][504] = 9'b111111111;
assign micromatrizz[53][505] = 9'b111111111;
assign micromatrizz[53][506] = 9'b111111111;
assign micromatrizz[53][507] = 9'b111110010;
assign micromatrizz[53][508] = 9'b111110010;
assign micromatrizz[53][509] = 9'b111110111;
assign micromatrizz[53][510] = 9'b111111111;
assign micromatrizz[53][511] = 9'b111111111;
assign micromatrizz[53][512] = 9'b111111111;
assign micromatrizz[53][513] = 9'b111111111;
assign micromatrizz[53][514] = 9'b111111111;
assign micromatrizz[53][515] = 9'b111111111;
assign micromatrizz[53][516] = 9'b111110111;
assign micromatrizz[53][517] = 9'b111110011;
assign micromatrizz[53][518] = 9'b111110011;
assign micromatrizz[53][519] = 9'b111110011;
assign micromatrizz[53][520] = 9'b111110010;
assign micromatrizz[53][521] = 9'b111110011;
assign micromatrizz[53][522] = 9'b111110011;
assign micromatrizz[53][523] = 9'b111110111;
assign micromatrizz[53][524] = 9'b111111111;
assign micromatrizz[53][525] = 9'b111110111;
assign micromatrizz[53][526] = 9'b111110110;
assign micromatrizz[53][527] = 9'b111110111;
assign micromatrizz[53][528] = 9'b111110011;
assign micromatrizz[53][529] = 9'b111110011;
assign micromatrizz[53][530] = 9'b111110010;
assign micromatrizz[53][531] = 9'b111110010;
assign micromatrizz[53][532] = 9'b111110111;
assign micromatrizz[53][533] = 9'b111111111;
assign micromatrizz[53][534] = 9'b111111111;
assign micromatrizz[53][535] = 9'b111111111;
assign micromatrizz[53][536] = 9'b111111111;
assign micromatrizz[53][537] = 9'b111111111;
assign micromatrizz[53][538] = 9'b111111111;
assign micromatrizz[53][539] = 9'b111111111;
assign micromatrizz[53][540] = 9'b111111111;
assign micromatrizz[53][541] = 9'b111111111;
assign micromatrizz[53][542] = 9'b111110111;
assign micromatrizz[53][543] = 9'b111110011;
assign micromatrizz[53][544] = 9'b111110010;
assign micromatrizz[53][545] = 9'b111110111;
assign micromatrizz[53][546] = 9'b111111111;
assign micromatrizz[53][547] = 9'b111111111;
assign micromatrizz[53][548] = 9'b111111111;
assign micromatrizz[53][549] = 9'b111110010;
assign micromatrizz[53][550] = 9'b111110010;
assign micromatrizz[53][551] = 9'b111111111;
assign micromatrizz[53][552] = 9'b111111111;
assign micromatrizz[53][553] = 9'b111111111;
assign micromatrizz[53][554] = 9'b111111111;
assign micromatrizz[53][555] = 9'b111111111;
assign micromatrizz[53][556] = 9'b111111111;
assign micromatrizz[53][557] = 9'b111111111;
assign micromatrizz[53][558] = 9'b111110010;
assign micromatrizz[53][559] = 9'b111110010;
assign micromatrizz[53][560] = 9'b111110010;
assign micromatrizz[53][561] = 9'b111110010;
assign micromatrizz[53][562] = 9'b111110011;
assign micromatrizz[53][563] = 9'b111110011;
assign micromatrizz[53][564] = 9'b111110010;
assign micromatrizz[53][565] = 9'b111111111;
assign micromatrizz[53][566] = 9'b111111111;
assign micromatrizz[53][567] = 9'b111111111;
assign micromatrizz[53][568] = 9'b111111111;
assign micromatrizz[53][569] = 9'b111111111;
assign micromatrizz[53][570] = 9'b111111111;
assign micromatrizz[53][571] = 9'b111111111;
assign micromatrizz[53][572] = 9'b111110010;
assign micromatrizz[53][573] = 9'b111110010;
assign micromatrizz[53][574] = 9'b111110010;
assign micromatrizz[53][575] = 9'b111110010;
assign micromatrizz[53][576] = 9'b111110011;
assign micromatrizz[53][577] = 9'b111110111;
assign micromatrizz[53][578] = 9'b111110110;
assign micromatrizz[53][579] = 9'b111111111;
assign micromatrizz[53][580] = 9'b111111111;
assign micromatrizz[53][581] = 9'b111110010;
assign micromatrizz[53][582] = 9'b111110011;
assign micromatrizz[53][583] = 9'b111110011;
assign micromatrizz[53][584] = 9'b111110010;
assign micromatrizz[53][585] = 9'b111110010;
assign micromatrizz[53][586] = 9'b111110011;
assign micromatrizz[53][587] = 9'b111110011;
assign micromatrizz[53][588] = 9'b111111111;
assign micromatrizz[53][589] = 9'b111111111;
assign micromatrizz[53][590] = 9'b111111111;
assign micromatrizz[53][591] = 9'b111111111;
assign micromatrizz[53][592] = 9'b111111111;
assign micromatrizz[53][593] = 9'b111111111;
assign micromatrizz[53][594] = 9'b111111111;
assign micromatrizz[53][595] = 9'b111110111;
assign micromatrizz[53][596] = 9'b111110010;
assign micromatrizz[53][597] = 9'b111110010;
assign micromatrizz[53][598] = 9'b111110111;
assign micromatrizz[53][599] = 9'b111111111;
assign micromatrizz[53][600] = 9'b111111111;
assign micromatrizz[53][601] = 9'b111110111;
assign micromatrizz[53][602] = 9'b111110010;
assign micromatrizz[53][603] = 9'b111110010;
assign micromatrizz[53][604] = 9'b111111111;
assign micromatrizz[53][605] = 9'b111111111;
assign micromatrizz[53][606] = 9'b111111111;
assign micromatrizz[53][607] = 9'b111111111;
assign micromatrizz[53][608] = 9'b111111111;
assign micromatrizz[53][609] = 9'b111111111;
assign micromatrizz[53][610] = 9'b111111111;
assign micromatrizz[53][611] = 9'b111111111;
assign micromatrizz[53][612] = 9'b111110111;
assign micromatrizz[53][613] = 9'b111110010;
assign micromatrizz[53][614] = 9'b111110010;
assign micromatrizz[53][615] = 9'b111110011;
assign micromatrizz[53][616] = 9'b111111111;
assign micromatrizz[53][617] = 9'b111111111;
assign micromatrizz[53][618] = 9'b111111111;
assign micromatrizz[53][619] = 9'b111111111;
assign micromatrizz[53][620] = 9'b111110111;
assign micromatrizz[53][621] = 9'b111110110;
assign micromatrizz[53][622] = 9'b111111111;
assign micromatrizz[53][623] = 9'b111111111;
assign micromatrizz[53][624] = 9'b111111111;
assign micromatrizz[53][625] = 9'b111111111;
assign micromatrizz[53][626] = 9'b111111111;
assign micromatrizz[53][627] = 9'b111111111;
assign micromatrizz[53][628] = 9'b111111111;
assign micromatrizz[53][629] = 9'b111111111;
assign micromatrizz[53][630] = 9'b111111111;
assign micromatrizz[53][631] = 9'b111111111;
assign micromatrizz[53][632] = 9'b111111111;
assign micromatrizz[53][633] = 9'b111111111;
assign micromatrizz[53][634] = 9'b111111111;
assign micromatrizz[53][635] = 9'b111111111;
assign micromatrizz[53][636] = 9'b111111111;
assign micromatrizz[53][637] = 9'b111111111;
assign micromatrizz[53][638] = 9'b111111111;
assign micromatrizz[53][639] = 9'b111111111;
assign micromatrizz[54][0] = 9'b111111111;
assign micromatrizz[54][1] = 9'b111111111;
assign micromatrizz[54][2] = 9'b111111111;
assign micromatrizz[54][3] = 9'b111111111;
assign micromatrizz[54][4] = 9'b111111111;
assign micromatrizz[54][5] = 9'b111111111;
assign micromatrizz[54][6] = 9'b111111111;
assign micromatrizz[54][7] = 9'b111111111;
assign micromatrizz[54][8] = 9'b111111111;
assign micromatrizz[54][9] = 9'b111110010;
assign micromatrizz[54][10] = 9'b111110010;
assign micromatrizz[54][11] = 9'b111110010;
assign micromatrizz[54][12] = 9'b111110010;
assign micromatrizz[54][13] = 9'b111110111;
assign micromatrizz[54][14] = 9'b111111111;
assign micromatrizz[54][15] = 9'b111111111;
assign micromatrizz[54][16] = 9'b111111111;
assign micromatrizz[54][17] = 9'b111111111;
assign micromatrizz[54][18] = 9'b111111111;
assign micromatrizz[54][19] = 9'b111111111;
assign micromatrizz[54][20] = 9'b111111111;
assign micromatrizz[54][21] = 9'b111111111;
assign micromatrizz[54][22] = 9'b111111111;
assign micromatrizz[54][23] = 9'b111110111;
assign micromatrizz[54][24] = 9'b111110010;
assign micromatrizz[54][25] = 9'b111110010;
assign micromatrizz[54][26] = 9'b111110010;
assign micromatrizz[54][27] = 9'b111110011;
assign micromatrizz[54][28] = 9'b111110011;
assign micromatrizz[54][29] = 9'b111110011;
assign micromatrizz[54][30] = 9'b111110011;
assign micromatrizz[54][31] = 9'b111111111;
assign micromatrizz[54][32] = 9'b111111111;
assign micromatrizz[54][33] = 9'b111111111;
assign micromatrizz[54][34] = 9'b111111111;
assign micromatrizz[54][35] = 9'b111110111;
assign micromatrizz[54][36] = 9'b111110010;
assign micromatrizz[54][37] = 9'b111110011;
assign micromatrizz[54][38] = 9'b111110011;
assign micromatrizz[54][39] = 9'b111110011;
assign micromatrizz[54][40] = 9'b111110011;
assign micromatrizz[54][41] = 9'b111110011;
assign micromatrizz[54][42] = 9'b111110011;
assign micromatrizz[54][43] = 9'b111111111;
assign micromatrizz[54][44] = 9'b111111111;
assign micromatrizz[54][45] = 9'b111111111;
assign micromatrizz[54][46] = 9'b111111111;
assign micromatrizz[54][47] = 9'b111110010;
assign micromatrizz[54][48] = 9'b111110010;
assign micromatrizz[54][49] = 9'b111110010;
assign micromatrizz[54][50] = 9'b111110011;
assign micromatrizz[54][51] = 9'b111110011;
assign micromatrizz[54][52] = 9'b111110010;
assign micromatrizz[54][53] = 9'b111110011;
assign micromatrizz[54][54] = 9'b111110010;
assign micromatrizz[54][55] = 9'b111110010;
assign micromatrizz[54][56] = 9'b111111111;
assign micromatrizz[54][57] = 9'b111111111;
assign micromatrizz[54][58] = 9'b111110111;
assign micromatrizz[54][59] = 9'b111110010;
assign micromatrizz[54][60] = 9'b111110010;
assign micromatrizz[54][61] = 9'b111110011;
assign micromatrizz[54][62] = 9'b111110010;
assign micromatrizz[54][63] = 9'b111110010;
assign micromatrizz[54][64] = 9'b111110111;
assign micromatrizz[54][65] = 9'b111111111;
assign micromatrizz[54][66] = 9'b111111111;
assign micromatrizz[54][67] = 9'b111111111;
assign micromatrizz[54][68] = 9'b111111111;
assign micromatrizz[54][69] = 9'b111111111;
assign micromatrizz[54][70] = 9'b111111111;
assign micromatrizz[54][71] = 9'b111110111;
assign micromatrizz[54][72] = 9'b111110010;
assign micromatrizz[54][73] = 9'b111110010;
assign micromatrizz[54][74] = 9'b111110011;
assign micromatrizz[54][75] = 9'b111111111;
assign micromatrizz[54][76] = 9'b111111111;
assign micromatrizz[54][77] = 9'b111111111;
assign micromatrizz[54][78] = 9'b111111111;
assign micromatrizz[54][79] = 9'b111110010;
assign micromatrizz[54][80] = 9'b111110011;
assign micromatrizz[54][81] = 9'b111110011;
assign micromatrizz[54][82] = 9'b111111111;
assign micromatrizz[54][83] = 9'b111111111;
assign micromatrizz[54][84] = 9'b111111111;
assign micromatrizz[54][85] = 9'b111111111;
assign micromatrizz[54][86] = 9'b111111111;
assign micromatrizz[54][87] = 9'b111111111;
assign micromatrizz[54][88] = 9'b111110010;
assign micromatrizz[54][89] = 9'b111110010;
assign micromatrizz[54][90] = 9'b111110010;
assign micromatrizz[54][91] = 9'b111110011;
assign micromatrizz[54][92] = 9'b111110011;
assign micromatrizz[54][93] = 9'b111110010;
assign micromatrizz[54][94] = 9'b111110011;
assign micromatrizz[54][95] = 9'b111110011;
assign micromatrizz[54][96] = 9'b111110011;
assign micromatrizz[54][97] = 9'b111110111;
assign micromatrizz[54][98] = 9'b111111111;
assign micromatrizz[54][99] = 9'b111111111;
assign micromatrizz[54][100] = 9'b111111111;
assign micromatrizz[54][101] = 9'b111111111;
assign micromatrizz[54][102] = 9'b111111111;
assign micromatrizz[54][103] = 9'b111111111;
assign micromatrizz[54][104] = 9'b111111111;
assign micromatrizz[54][105] = 9'b111110010;
assign micromatrizz[54][106] = 9'b111110010;
assign micromatrizz[54][107] = 9'b111110011;
assign micromatrizz[54][108] = 9'b111110010;
assign micromatrizz[54][109] = 9'b111110011;
assign micromatrizz[54][110] = 9'b111111111;
assign micromatrizz[54][111] = 9'b111111111;
assign micromatrizz[54][112] = 9'b111111111;
assign micromatrizz[54][113] = 9'b111111111;
assign micromatrizz[54][114] = 9'b111111111;
assign micromatrizz[54][115] = 9'b111111111;
assign micromatrizz[54][116] = 9'b111111111;
assign micromatrizz[54][117] = 9'b111111111;
assign micromatrizz[54][118] = 9'b111111111;
assign micromatrizz[54][119] = 9'b111111111;
assign micromatrizz[54][120] = 9'b111111111;
assign micromatrizz[54][121] = 9'b111110111;
assign micromatrizz[54][122] = 9'b111110010;
assign micromatrizz[54][123] = 9'b111110010;
assign micromatrizz[54][124] = 9'b111110011;
assign micromatrizz[54][125] = 9'b111110011;
assign micromatrizz[54][126] = 9'b111110111;
assign micromatrizz[54][127] = 9'b111111111;
assign micromatrizz[54][128] = 9'b111111111;
assign micromatrizz[54][129] = 9'b111111111;
assign micromatrizz[54][130] = 9'b111111111;
assign micromatrizz[54][131] = 9'b111111111;
assign micromatrizz[54][132] = 9'b111110111;
assign micromatrizz[54][133] = 9'b111111111;
assign micromatrizz[54][134] = 9'b111111111;
assign micromatrizz[54][135] = 9'b111111111;
assign micromatrizz[54][136] = 9'b111111111;
assign micromatrizz[54][137] = 9'b111111111;
assign micromatrizz[54][138] = 9'b111110111;
assign micromatrizz[54][139] = 9'b111110010;
assign micromatrizz[54][140] = 9'b111110010;
assign micromatrizz[54][141] = 9'b111110010;
assign micromatrizz[54][142] = 9'b111110010;
assign micromatrizz[54][143] = 9'b111110011;
assign micromatrizz[54][144] = 9'b111110011;
assign micromatrizz[54][145] = 9'b111110010;
assign micromatrizz[54][146] = 9'b111110111;
assign micromatrizz[54][147] = 9'b111111111;
assign micromatrizz[54][148] = 9'b111111111;
assign micromatrizz[54][149] = 9'b111111111;
assign micromatrizz[54][150] = 9'b111110111;
assign micromatrizz[54][151] = 9'b111110010;
assign micromatrizz[54][152] = 9'b111110010;
assign micromatrizz[54][153] = 9'b111110011;
assign micromatrizz[54][154] = 9'b111110011;
assign micromatrizz[54][155] = 9'b111110011;
assign micromatrizz[54][156] = 9'b111110010;
assign micromatrizz[54][157] = 9'b111111111;
assign micromatrizz[54][158] = 9'b111111111;
assign micromatrizz[54][159] = 9'b111111111;
assign micromatrizz[54][160] = 9'b111111111;
assign micromatrizz[54][161] = 9'b111111111;
assign micromatrizz[54][162] = 9'b111111111;
assign micromatrizz[54][163] = 9'b111110010;
assign micromatrizz[54][164] = 9'b111110010;
assign micromatrizz[54][165] = 9'b111111111;
assign micromatrizz[54][166] = 9'b111111111;
assign micromatrizz[54][167] = 9'b111111111;
assign micromatrizz[54][168] = 9'b111111111;
assign micromatrizz[54][169] = 9'b111111111;
assign micromatrizz[54][170] = 9'b111111111;
assign micromatrizz[54][171] = 9'b111111111;
assign micromatrizz[54][172] = 9'b111110010;
assign micromatrizz[54][173] = 9'b111110010;
assign micromatrizz[54][174] = 9'b111110010;
assign micromatrizz[54][175] = 9'b111110010;
assign micromatrizz[54][176] = 9'b111110011;
assign micromatrizz[54][177] = 9'b111110010;
assign micromatrizz[54][178] = 9'b111110111;
assign micromatrizz[54][179] = 9'b111111111;
assign micromatrizz[54][180] = 9'b111111111;
assign micromatrizz[54][181] = 9'b111111111;
assign micromatrizz[54][182] = 9'b111111111;
assign micromatrizz[54][183] = 9'b111111111;
assign micromatrizz[54][184] = 9'b111111111;
assign micromatrizz[54][185] = 9'b111110010;
assign micromatrizz[54][186] = 9'b111110010;
assign micromatrizz[54][187] = 9'b111110011;
assign micromatrizz[54][188] = 9'b111110010;
assign micromatrizz[54][189] = 9'b111110010;
assign micromatrizz[54][190] = 9'b111110111;
assign micromatrizz[54][191] = 9'b111111111;
assign micromatrizz[54][192] = 9'b111111111;
assign micromatrizz[54][193] = 9'b111110111;
assign micromatrizz[54][194] = 9'b111110010;
assign micromatrizz[54][195] = 9'b111110010;
assign micromatrizz[54][196] = 9'b111110010;
assign micromatrizz[54][197] = 9'b111110011;
assign micromatrizz[54][198] = 9'b111110011;
assign micromatrizz[54][199] = 9'b111110010;
assign micromatrizz[54][200] = 9'b111110010;
assign micromatrizz[54][201] = 9'b111110011;
assign micromatrizz[54][202] = 9'b111110111;
assign micromatrizz[54][203] = 9'b111111111;
assign micromatrizz[54][204] = 9'b111111111;
assign micromatrizz[54][205] = 9'b111111111;
assign micromatrizz[54][206] = 9'b111111111;
assign micromatrizz[54][207] = 9'b111111111;
assign micromatrizz[54][208] = 9'b111110111;
assign micromatrizz[54][209] = 9'b111110010;
assign micromatrizz[54][210] = 9'b111110011;
assign micromatrizz[54][211] = 9'b111110011;
assign micromatrizz[54][212] = 9'b111110010;
assign micromatrizz[54][213] = 9'b111110111;
assign micromatrizz[54][214] = 9'b111111111;
assign micromatrizz[54][215] = 9'b111111111;
assign micromatrizz[54][216] = 9'b111111111;
assign micromatrizz[54][217] = 9'b111111111;
assign micromatrizz[54][218] = 9'b111110111;
assign micromatrizz[54][219] = 9'b111110111;
assign micromatrizz[54][220] = 9'b111111111;
assign micromatrizz[54][221] = 9'b111111111;
assign micromatrizz[54][222] = 9'b111111111;
assign micromatrizz[54][223] = 9'b111111111;
assign micromatrizz[54][224] = 9'b111111111;
assign micromatrizz[54][225] = 9'b111110111;
assign micromatrizz[54][226] = 9'b111110010;
assign micromatrizz[54][227] = 9'b111110010;
assign micromatrizz[54][228] = 9'b111110010;
assign micromatrizz[54][229] = 9'b111110011;
assign micromatrizz[54][230] = 9'b111110011;
assign micromatrizz[54][231] = 9'b111110011;
assign micromatrizz[54][232] = 9'b111110011;
assign micromatrizz[54][233] = 9'b111110111;
assign micromatrizz[54][234] = 9'b111110111;
assign micromatrizz[54][235] = 9'b111111111;
assign micromatrizz[54][236] = 9'b111111111;
assign micromatrizz[54][237] = 9'b111111111;
assign micromatrizz[54][238] = 9'b111111111;
assign micromatrizz[54][239] = 9'b111111111;
assign micromatrizz[54][240] = 9'b111111111;
assign micromatrizz[54][241] = 9'b111111111;
assign micromatrizz[54][242] = 9'b111111111;
assign micromatrizz[54][243] = 9'b111110111;
assign micromatrizz[54][244] = 9'b111110010;
assign micromatrizz[54][245] = 9'b111110010;
assign micromatrizz[54][246] = 9'b111110010;
assign micromatrizz[54][247] = 9'b111110111;
assign micromatrizz[54][248] = 9'b111111111;
assign micromatrizz[54][249] = 9'b111111111;
assign micromatrizz[54][250] = 9'b111111111;
assign micromatrizz[54][251] = 9'b111110111;
assign micromatrizz[54][252] = 9'b111110010;
assign micromatrizz[54][253] = 9'b111110010;
assign micromatrizz[54][254] = 9'b111110111;
assign micromatrizz[54][255] = 9'b111111111;
assign micromatrizz[54][256] = 9'b111111111;
assign micromatrizz[54][257] = 9'b111111111;
assign micromatrizz[54][258] = 9'b111111111;
assign micromatrizz[54][259] = 9'b111111111;
assign micromatrizz[54][260] = 9'b111111111;
assign micromatrizz[54][261] = 9'b111110010;
assign micromatrizz[54][262] = 9'b111110011;
assign micromatrizz[54][263] = 9'b111110011;
assign micromatrizz[54][264] = 9'b111110010;
assign micromatrizz[54][265] = 9'b111110111;
assign micromatrizz[54][266] = 9'b111111111;
assign micromatrizz[54][267] = 9'b111111111;
assign micromatrizz[54][268] = 9'b111111111;
assign micromatrizz[54][269] = 9'b111111111;
assign micromatrizz[54][270] = 9'b111111111;
assign micromatrizz[54][271] = 9'b111111111;
assign micromatrizz[54][272] = 9'b111111111;
assign micromatrizz[54][273] = 9'b111111111;
assign micromatrizz[54][274] = 9'b111111111;
assign micromatrizz[54][275] = 9'b111111111;
assign micromatrizz[54][276] = 9'b111111111;
assign micromatrizz[54][277] = 9'b111110010;
assign micromatrizz[54][278] = 9'b111110111;
assign micromatrizz[54][279] = 9'b111111111;
assign micromatrizz[54][280] = 9'b111111111;
assign micromatrizz[54][281] = 9'b111111111;
assign micromatrizz[54][282] = 9'b111111111;
assign micromatrizz[54][283] = 9'b111111111;
assign micromatrizz[54][284] = 9'b111111111;
assign micromatrizz[54][285] = 9'b111111111;
assign micromatrizz[54][286] = 9'b111110010;
assign micromatrizz[54][287] = 9'b111110010;
assign micromatrizz[54][288] = 9'b111110010;
assign micromatrizz[54][289] = 9'b111110010;
assign micromatrizz[54][290] = 9'b111110011;
assign micromatrizz[54][291] = 9'b111110010;
assign micromatrizz[54][292] = 9'b111110111;
assign micromatrizz[54][293] = 9'b111111111;
assign micromatrizz[54][294] = 9'b111111111;
assign micromatrizz[54][295] = 9'b111111111;
assign micromatrizz[54][296] = 9'b111110111;
assign micromatrizz[54][297] = 9'b111110010;
assign micromatrizz[54][298] = 9'b111110010;
assign micromatrizz[54][299] = 9'b111110010;
assign micromatrizz[54][300] = 9'b111110010;
assign micromatrizz[54][301] = 9'b111110010;
assign micromatrizz[54][302] = 9'b111110011;
assign micromatrizz[54][303] = 9'b111110010;
assign micromatrizz[54][304] = 9'b111110010;
assign micromatrizz[54][305] = 9'b111110111;
assign micromatrizz[54][306] = 9'b111111111;
assign micromatrizz[54][307] = 9'b111111111;
assign micromatrizz[54][308] = 9'b111111111;
assign micromatrizz[54][309] = 9'b111111111;
assign micromatrizz[54][310] = 9'b111111111;
assign micromatrizz[54][311] = 9'b111111111;
assign micromatrizz[54][312] = 9'b111110111;
assign micromatrizz[54][313] = 9'b111110010;
assign micromatrizz[54][314] = 9'b111111111;
assign micromatrizz[54][315] = 9'b111111111;
assign micromatrizz[54][316] = 9'b111111111;
assign micromatrizz[54][317] = 9'b111111111;
assign micromatrizz[54][318] = 9'b111110111;
assign micromatrizz[54][319] = 9'b111110010;
assign micromatrizz[54][320] = 9'b111110011;
assign micromatrizz[54][321] = 9'b111110011;
assign micromatrizz[54][322] = 9'b111111111;
assign micromatrizz[54][323] = 9'b111111111;
assign micromatrizz[54][324] = 9'b111111111;
assign micromatrizz[54][325] = 9'b111111111;
assign micromatrizz[54][326] = 9'b111110010;
assign micromatrizz[54][327] = 9'b111110010;
assign micromatrizz[54][328] = 9'b111110010;
assign micromatrizz[54][329] = 9'b111110111;
assign micromatrizz[54][330] = 9'b111111111;
assign micromatrizz[54][331] = 9'b111111111;
assign micromatrizz[54][332] = 9'b111111111;
assign micromatrizz[54][333] = 9'b111111111;
assign micromatrizz[54][334] = 9'b111111111;
assign micromatrizz[54][335] = 9'b111110010;
assign micromatrizz[54][336] = 9'b111110010;
assign micromatrizz[54][337] = 9'b111110011;
assign micromatrizz[54][338] = 9'b111110011;
assign micromatrizz[54][339] = 9'b111110011;
assign micromatrizz[54][340] = 9'b111110011;
assign micromatrizz[54][341] = 9'b111110011;
assign micromatrizz[54][342] = 9'b111110011;
assign micromatrizz[54][343] = 9'b111110111;
assign micromatrizz[54][344] = 9'b111111111;
assign micromatrizz[54][345] = 9'b111111111;
assign micromatrizz[54][346] = 9'b111111111;
assign micromatrizz[54][347] = 9'b111110010;
assign micromatrizz[54][348] = 9'b111110010;
assign micromatrizz[54][349] = 9'b111110011;
assign micromatrizz[54][350] = 9'b111110011;
assign micromatrizz[54][351] = 9'b111110011;
assign micromatrizz[54][352] = 9'b111110011;
assign micromatrizz[54][353] = 9'b111110111;
assign micromatrizz[54][354] = 9'b111111111;
assign micromatrizz[54][355] = 9'b111111111;
assign micromatrizz[54][356] = 9'b111111111;
assign micromatrizz[54][357] = 9'b111111111;
assign micromatrizz[54][358] = 9'b111111111;
assign micromatrizz[54][359] = 9'b111110010;
assign micromatrizz[54][360] = 9'b111110011;
assign micromatrizz[54][361] = 9'b111110010;
assign micromatrizz[54][362] = 9'b111110010;
assign micromatrizz[54][363] = 9'b111110011;
assign micromatrizz[54][364] = 9'b111110011;
assign micromatrizz[54][365] = 9'b111110010;
assign micromatrizz[54][366] = 9'b111111111;
assign micromatrizz[54][367] = 9'b111111111;
assign micromatrizz[54][368] = 9'b111111111;
assign micromatrizz[54][369] = 9'b111111111;
assign micromatrizz[54][370] = 9'b111111111;
assign micromatrizz[54][371] = 9'b111111111;
assign micromatrizz[54][372] = 9'b111110010;
assign micromatrizz[54][373] = 9'b111110011;
assign micromatrizz[54][374] = 9'b111110011;
assign micromatrizz[54][375] = 9'b111110011;
assign micromatrizz[54][376] = 9'b111110011;
assign micromatrizz[54][377] = 9'b111110011;
assign micromatrizz[54][378] = 9'b111110011;
assign micromatrizz[54][379] = 9'b111111111;
assign micromatrizz[54][380] = 9'b111111111;
assign micromatrizz[54][381] = 9'b111111111;
assign micromatrizz[54][382] = 9'b111111111;
assign micromatrizz[54][383] = 9'b111110111;
assign micromatrizz[54][384] = 9'b111110010;
assign micromatrizz[54][385] = 9'b111110010;
assign micromatrizz[54][386] = 9'b111110011;
assign micromatrizz[54][387] = 9'b111110011;
assign micromatrizz[54][388] = 9'b111110011;
assign micromatrizz[54][389] = 9'b111110011;
assign micromatrizz[54][390] = 9'b111110010;
assign micromatrizz[54][391] = 9'b111111111;
assign micromatrizz[54][392] = 9'b111111111;
assign micromatrizz[54][393] = 9'b111111111;
assign micromatrizz[54][394] = 9'b111111111;
assign micromatrizz[54][395] = 9'b111110111;
assign micromatrizz[54][396] = 9'b111110010;
assign micromatrizz[54][397] = 9'b111110010;
assign micromatrizz[54][398] = 9'b111110010;
assign micromatrizz[54][399] = 9'b111110011;
assign micromatrizz[54][400] = 9'b111110011;
assign micromatrizz[54][401] = 9'b111110011;
assign micromatrizz[54][402] = 9'b111110011;
assign micromatrizz[54][403] = 9'b111110111;
assign micromatrizz[54][404] = 9'b111110111;
assign micromatrizz[54][405] = 9'b111111111;
assign micromatrizz[54][406] = 9'b111111111;
assign micromatrizz[54][407] = 9'b111111111;
assign micromatrizz[54][408] = 9'b111111111;
assign micromatrizz[54][409] = 9'b111111111;
assign micromatrizz[54][410] = 9'b111111111;
assign micromatrizz[54][411] = 9'b111111111;
assign micromatrizz[54][412] = 9'b111111111;
assign micromatrizz[54][413] = 9'b111110111;
assign micromatrizz[54][414] = 9'b111110011;
assign micromatrizz[54][415] = 9'b111110010;
assign micromatrizz[54][416] = 9'b111110010;
assign micromatrizz[54][417] = 9'b111110111;
assign micromatrizz[54][418] = 9'b111111111;
assign micromatrizz[54][419] = 9'b111111111;
assign micromatrizz[54][420] = 9'b111111111;
assign micromatrizz[54][421] = 9'b111110111;
assign micromatrizz[54][422] = 9'b111110010;
assign micromatrizz[54][423] = 9'b111110010;
assign micromatrizz[54][424] = 9'b111110111;
assign micromatrizz[54][425] = 9'b111111111;
assign micromatrizz[54][426] = 9'b111111111;
assign micromatrizz[54][427] = 9'b111111111;
assign micromatrizz[54][428] = 9'b111111111;
assign micromatrizz[54][429] = 9'b111111111;
assign micromatrizz[54][430] = 9'b111110111;
assign micromatrizz[54][431] = 9'b111110010;
assign micromatrizz[54][432] = 9'b111110010;
assign micromatrizz[54][433] = 9'b111110010;
assign micromatrizz[54][434] = 9'b111110011;
assign micromatrizz[54][435] = 9'b111110011;
assign micromatrizz[54][436] = 9'b111110011;
assign micromatrizz[54][437] = 9'b111110011;
assign micromatrizz[54][438] = 9'b111110111;
assign micromatrizz[54][439] = 9'b111110111;
assign micromatrizz[54][440] = 9'b111111111;
assign micromatrizz[54][441] = 9'b111111111;
assign micromatrizz[54][442] = 9'b111111111;
assign micromatrizz[54][443] = 9'b111111111;
assign micromatrizz[54][444] = 9'b111111111;
assign micromatrizz[54][445] = 9'b111111111;
assign micromatrizz[54][446] = 9'b111111111;
assign micromatrizz[54][447] = 9'b111111111;
assign micromatrizz[54][448] = 9'b111111111;
assign micromatrizz[54][449] = 9'b111110010;
assign micromatrizz[54][450] = 9'b111110010;
assign micromatrizz[54][451] = 9'b111110011;
assign micromatrizz[54][452] = 9'b111110011;
assign micromatrizz[54][453] = 9'b111110011;
assign micromatrizz[54][454] = 9'b111111111;
assign micromatrizz[54][455] = 9'b111111111;
assign micromatrizz[54][456] = 9'b111111111;
assign micromatrizz[54][457] = 9'b111111111;
assign micromatrizz[54][458] = 9'b111111111;
assign micromatrizz[54][459] = 9'b111110111;
assign micromatrizz[54][460] = 9'b111111111;
assign micromatrizz[54][461] = 9'b111111111;
assign micromatrizz[54][462] = 9'b111111111;
assign micromatrizz[54][463] = 9'b111111111;
assign micromatrizz[54][464] = 9'b111111111;
assign micromatrizz[54][465] = 9'b111111111;
assign micromatrizz[54][466] = 9'b111110010;
assign micromatrizz[54][467] = 9'b111110010;
assign micromatrizz[54][468] = 9'b111110011;
assign micromatrizz[54][469] = 9'b111110010;
assign micromatrizz[54][470] = 9'b111110111;
assign micromatrizz[54][471] = 9'b111111111;
assign micromatrizz[54][472] = 9'b111111111;
assign micromatrizz[54][473] = 9'b111111111;
assign micromatrizz[54][474] = 9'b111111111;
assign micromatrizz[54][475] = 9'b111111111;
assign micromatrizz[54][476] = 9'b111111111;
assign micromatrizz[54][477] = 9'b111111111;
assign micromatrizz[54][478] = 9'b111111111;
assign micromatrizz[54][479] = 9'b111111111;
assign micromatrizz[54][480] = 9'b111111111;
assign micromatrizz[54][481] = 9'b111110010;
assign micromatrizz[54][482] = 9'b111110010;
assign micromatrizz[54][483] = 9'b111110010;
assign micromatrizz[54][484] = 9'b111110010;
assign micromatrizz[54][485] = 9'b111110011;
assign micromatrizz[54][486] = 9'b111110011;
assign micromatrizz[54][487] = 9'b111110010;
assign micromatrizz[54][488] = 9'b111110111;
assign micromatrizz[54][489] = 9'b111110011;
assign micromatrizz[54][490] = 9'b111110111;
assign micromatrizz[54][491] = 9'b111111111;
assign micromatrizz[54][492] = 9'b111111111;
assign micromatrizz[54][493] = 9'b111111111;
assign micromatrizz[54][494] = 9'b111111111;
assign micromatrizz[54][495] = 9'b111111111;
assign micromatrizz[54][496] = 9'b111111111;
assign micromatrizz[54][497] = 9'b111111111;
assign micromatrizz[54][498] = 9'b111111111;
assign micromatrizz[54][499] = 9'b111110111;
assign micromatrizz[54][500] = 9'b111110010;
assign micromatrizz[54][501] = 9'b111110011;
assign micromatrizz[54][502] = 9'b111110010;
assign micromatrizz[54][503] = 9'b111110111;
assign micromatrizz[54][504] = 9'b111111111;
assign micromatrizz[54][505] = 9'b111111111;
assign micromatrizz[54][506] = 9'b111111111;
assign micromatrizz[54][507] = 9'b111110010;
assign micromatrizz[54][508] = 9'b111110010;
assign micromatrizz[54][509] = 9'b111110010;
assign micromatrizz[54][510] = 9'b111110111;
assign micromatrizz[54][511] = 9'b111111111;
assign micromatrizz[54][512] = 9'b111111111;
assign micromatrizz[54][513] = 9'b111111111;
assign micromatrizz[54][514] = 9'b111111111;
assign micromatrizz[54][515] = 9'b111111111;
assign micromatrizz[54][516] = 9'b111110111;
assign micromatrizz[54][517] = 9'b111110010;
assign micromatrizz[54][518] = 9'b111110011;
assign micromatrizz[54][519] = 9'b111110011;
assign micromatrizz[54][520] = 9'b111110010;
assign micromatrizz[54][521] = 9'b111110010;
assign micromatrizz[54][522] = 9'b111110011;
assign micromatrizz[54][523] = 9'b111110011;
assign micromatrizz[54][524] = 9'b111110010;
assign micromatrizz[54][525] = 9'b111110111;
assign micromatrizz[54][526] = 9'b111111111;
assign micromatrizz[54][527] = 9'b111111111;
assign micromatrizz[54][528] = 9'b111110111;
assign micromatrizz[54][529] = 9'b111110010;
assign micromatrizz[54][530] = 9'b111110011;
assign micromatrizz[54][531] = 9'b111110011;
assign micromatrizz[54][532] = 9'b111110011;
assign micromatrizz[54][533] = 9'b111110010;
assign micromatrizz[54][534] = 9'b111111111;
assign micromatrizz[54][535] = 9'b111111111;
assign micromatrizz[54][536] = 9'b111111111;
assign micromatrizz[54][537] = 9'b111111111;
assign micromatrizz[54][538] = 9'b111111111;
assign micromatrizz[54][539] = 9'b111111111;
assign micromatrizz[54][540] = 9'b111111111;
assign micromatrizz[54][541] = 9'b111110111;
assign micromatrizz[54][542] = 9'b111110010;
assign micromatrizz[54][543] = 9'b111110011;
assign micromatrizz[54][544] = 9'b111110010;
assign micromatrizz[54][545] = 9'b111111111;
assign micromatrizz[54][546] = 9'b111111111;
assign micromatrizz[54][547] = 9'b111111111;
assign micromatrizz[54][548] = 9'b111111111;
assign micromatrizz[54][549] = 9'b111110010;
assign micromatrizz[54][550] = 9'b111110010;
assign micromatrizz[54][551] = 9'b111110010;
assign micromatrizz[54][552] = 9'b111111111;
assign micromatrizz[54][553] = 9'b111111111;
assign micromatrizz[54][554] = 9'b111111111;
assign micromatrizz[54][555] = 9'b111111111;
assign micromatrizz[54][556] = 9'b111111111;
assign micromatrizz[54][557] = 9'b111111111;
assign micromatrizz[54][558] = 9'b111110010;
assign micromatrizz[54][559] = 9'b111110010;
assign micromatrizz[54][560] = 9'b111110010;
assign micromatrizz[54][561] = 9'b111110010;
assign micromatrizz[54][562] = 9'b111110011;
assign micromatrizz[54][563] = 9'b111110011;
assign micromatrizz[54][564] = 9'b111110010;
assign micromatrizz[54][565] = 9'b111111111;
assign micromatrizz[54][566] = 9'b111111111;
assign micromatrizz[54][567] = 9'b111111111;
assign micromatrizz[54][568] = 9'b111111111;
assign micromatrizz[54][569] = 9'b111111111;
assign micromatrizz[54][570] = 9'b111110111;
assign micromatrizz[54][571] = 9'b111110010;
assign micromatrizz[54][572] = 9'b111110010;
assign micromatrizz[54][573] = 9'b111110011;
assign micromatrizz[54][574] = 9'b111110011;
assign micromatrizz[54][575] = 9'b111110010;
assign micromatrizz[54][576] = 9'b111111111;
assign micromatrizz[54][577] = 9'b111111111;
assign micromatrizz[54][578] = 9'b111111111;
assign micromatrizz[54][579] = 9'b111110010;
assign micromatrizz[54][580] = 9'b111110010;
assign micromatrizz[54][581] = 9'b111110010;
assign micromatrizz[54][582] = 9'b111110011;
assign micromatrizz[54][583] = 9'b111110011;
assign micromatrizz[54][584] = 9'b111110010;
assign micromatrizz[54][585] = 9'b111110010;
assign micromatrizz[54][586] = 9'b111110011;
assign micromatrizz[54][587] = 9'b111110011;
assign micromatrizz[54][588] = 9'b111111111;
assign micromatrizz[54][589] = 9'b111111111;
assign micromatrizz[54][590] = 9'b111111111;
assign micromatrizz[54][591] = 9'b111111111;
assign micromatrizz[54][592] = 9'b111111111;
assign micromatrizz[54][593] = 9'b111111111;
assign micromatrizz[54][594] = 9'b111110111;
assign micromatrizz[54][595] = 9'b111110010;
assign micromatrizz[54][596] = 9'b111110010;
assign micromatrizz[54][597] = 9'b111110010;
assign micromatrizz[54][598] = 9'b111111111;
assign micromatrizz[54][599] = 9'b111111111;
assign micromatrizz[54][600] = 9'b111111111;
assign micromatrizz[54][601] = 9'b111111111;
assign micromatrizz[54][602] = 9'b111110010;
assign micromatrizz[54][603] = 9'b111110010;
assign micromatrizz[54][604] = 9'b111110010;
assign micromatrizz[54][605] = 9'b111111111;
assign micromatrizz[54][606] = 9'b111111111;
assign micromatrizz[54][607] = 9'b111111111;
assign micromatrizz[54][608] = 9'b111111111;
assign micromatrizz[54][609] = 9'b111111111;
assign micromatrizz[54][610] = 9'b111111111;
assign micromatrizz[54][611] = 9'b111110010;
assign micromatrizz[54][612] = 9'b111110010;
assign micromatrizz[54][613] = 9'b111110010;
assign micromatrizz[54][614] = 9'b111110010;
assign micromatrizz[54][615] = 9'b111110011;
assign micromatrizz[54][616] = 9'b111111111;
assign micromatrizz[54][617] = 9'b111111111;
assign micromatrizz[54][618] = 9'b111111111;
assign micromatrizz[54][619] = 9'b111111111;
assign micromatrizz[54][620] = 9'b111111111;
assign micromatrizz[54][621] = 9'b111111111;
assign micromatrizz[54][622] = 9'b111111111;
assign micromatrizz[54][623] = 9'b111111111;
assign micromatrizz[54][624] = 9'b111111111;
assign micromatrizz[54][625] = 9'b111111111;
assign micromatrizz[54][626] = 9'b111111111;
assign micromatrizz[54][627] = 9'b111111111;
assign micromatrizz[54][628] = 9'b111111111;
assign micromatrizz[54][629] = 9'b111111111;
assign micromatrizz[54][630] = 9'b111111111;
assign micromatrizz[54][631] = 9'b111111111;
assign micromatrizz[54][632] = 9'b111111111;
assign micromatrizz[54][633] = 9'b111111111;
assign micromatrizz[54][634] = 9'b111111111;
assign micromatrizz[54][635] = 9'b111111111;
assign micromatrizz[54][636] = 9'b111111111;
assign micromatrizz[54][637] = 9'b111111111;
assign micromatrizz[54][638] = 9'b111111111;
assign micromatrizz[54][639] = 9'b111111111;
assign micromatrizz[55][0] = 9'b111111111;
assign micromatrizz[55][1] = 9'b111111111;
assign micromatrizz[55][2] = 9'b111111111;
assign micromatrizz[55][3] = 9'b111111111;
assign micromatrizz[55][4] = 9'b111111111;
assign micromatrizz[55][5] = 9'b111111111;
assign micromatrizz[55][6] = 9'b111111111;
assign micromatrizz[55][7] = 9'b111111111;
assign micromatrizz[55][8] = 9'b111110110;
assign micromatrizz[55][9] = 9'b111110010;
assign micromatrizz[55][10] = 9'b111110010;
assign micromatrizz[55][11] = 9'b111110010;
assign micromatrizz[55][12] = 9'b111110011;
assign micromatrizz[55][13] = 9'b111110011;
assign micromatrizz[55][14] = 9'b111111111;
assign micromatrizz[55][15] = 9'b111111111;
assign micromatrizz[55][16] = 9'b111111111;
assign micromatrizz[55][17] = 9'b111111111;
assign micromatrizz[55][18] = 9'b111111111;
assign micromatrizz[55][19] = 9'b111111111;
assign micromatrizz[55][20] = 9'b111111111;
assign micromatrizz[55][21] = 9'b111111111;
assign micromatrizz[55][22] = 9'b111111111;
assign micromatrizz[55][23] = 9'b111110111;
assign micromatrizz[55][24] = 9'b111110010;
assign micromatrizz[55][25] = 9'b111110010;
assign micromatrizz[55][26] = 9'b111110010;
assign micromatrizz[55][27] = 9'b111110011;
assign micromatrizz[55][28] = 9'b111110011;
assign micromatrizz[55][29] = 9'b111110011;
assign micromatrizz[55][30] = 9'b111110011;
assign micromatrizz[55][31] = 9'b111111111;
assign micromatrizz[55][32] = 9'b111111111;
assign micromatrizz[55][33] = 9'b111111111;
assign micromatrizz[55][34] = 9'b111111111;
assign micromatrizz[55][35] = 9'b111110111;
assign micromatrizz[55][36] = 9'b111110010;
assign micromatrizz[55][37] = 9'b111110010;
assign micromatrizz[55][38] = 9'b111110010;
assign micromatrizz[55][39] = 9'b111110011;
assign micromatrizz[55][40] = 9'b111110011;
assign micromatrizz[55][41] = 9'b111110011;
assign micromatrizz[55][42] = 9'b111110011;
assign micromatrizz[55][43] = 9'b111111111;
assign micromatrizz[55][44] = 9'b111111111;
assign micromatrizz[55][45] = 9'b111111111;
assign micromatrizz[55][46] = 9'b111111111;
assign micromatrizz[55][47] = 9'b111110010;
assign micromatrizz[55][48] = 9'b111110010;
assign micromatrizz[55][49] = 9'b111110010;
assign micromatrizz[55][50] = 9'b111110011;
assign micromatrizz[55][51] = 9'b111110011;
assign micromatrizz[55][52] = 9'b111110010;
assign micromatrizz[55][53] = 9'b111110010;
assign micromatrizz[55][54] = 9'b111110011;
assign micromatrizz[55][55] = 9'b111111111;
assign micromatrizz[55][56] = 9'b111111111;
assign micromatrizz[55][57] = 9'b111111111;
assign micromatrizz[55][58] = 9'b111111111;
assign micromatrizz[55][59] = 9'b111110010;
assign micromatrizz[55][60] = 9'b111110010;
assign micromatrizz[55][61] = 9'b111110011;
assign micromatrizz[55][62] = 9'b111110010;
assign micromatrizz[55][63] = 9'b111110011;
assign micromatrizz[55][64] = 9'b111110010;
assign micromatrizz[55][65] = 9'b111110111;
assign micromatrizz[55][66] = 9'b111111111;
assign micromatrizz[55][67] = 9'b111111111;
assign micromatrizz[55][68] = 9'b111111111;
assign micromatrizz[55][69] = 9'b111111111;
assign micromatrizz[55][70] = 9'b111110111;
assign micromatrizz[55][71] = 9'b111110010;
assign micromatrizz[55][72] = 9'b111110011;
assign micromatrizz[55][73] = 9'b111110011;
assign micromatrizz[55][74] = 9'b111110011;
assign micromatrizz[55][75] = 9'b111111111;
assign micromatrizz[55][76] = 9'b111111111;
assign micromatrizz[55][77] = 9'b111111111;
assign micromatrizz[55][78] = 9'b111111111;
assign micromatrizz[55][79] = 9'b111110010;
assign micromatrizz[55][80] = 9'b111110011;
assign micromatrizz[55][81] = 9'b111110011;
assign micromatrizz[55][82] = 9'b111110010;
assign micromatrizz[55][83] = 9'b111111111;
assign micromatrizz[55][84] = 9'b111111111;
assign micromatrizz[55][85] = 9'b111111111;
assign micromatrizz[55][86] = 9'b111111111;
assign micromatrizz[55][87] = 9'b111111111;
assign micromatrizz[55][88] = 9'b111110010;
assign micromatrizz[55][89] = 9'b111110010;
assign micromatrizz[55][90] = 9'b111110010;
assign micromatrizz[55][91] = 9'b111110010;
assign micromatrizz[55][92] = 9'b111110010;
assign micromatrizz[55][93] = 9'b111110011;
assign micromatrizz[55][94] = 9'b111110011;
assign micromatrizz[55][95] = 9'b111110011;
assign micromatrizz[55][96] = 9'b111110111;
assign micromatrizz[55][97] = 9'b111111111;
assign micromatrizz[55][98] = 9'b111111111;
assign micromatrizz[55][99] = 9'b111111111;
assign micromatrizz[55][100] = 9'b111111111;
assign micromatrizz[55][101] = 9'b111111111;
assign micromatrizz[55][102] = 9'b111111111;
assign micromatrizz[55][103] = 9'b111111111;
assign micromatrizz[55][104] = 9'b111110111;
assign micromatrizz[55][105] = 9'b111110010;
assign micromatrizz[55][106] = 9'b111110010;
assign micromatrizz[55][107] = 9'b111110011;
assign micromatrizz[55][108] = 9'b111110011;
assign micromatrizz[55][109] = 9'b111110011;
assign micromatrizz[55][110] = 9'b111110111;
assign micromatrizz[55][111] = 9'b111111111;
assign micromatrizz[55][112] = 9'b111111111;
assign micromatrizz[55][113] = 9'b111111111;
assign micromatrizz[55][114] = 9'b111111111;
assign micromatrizz[55][115] = 9'b111111111;
assign micromatrizz[55][116] = 9'b111111111;
assign micromatrizz[55][117] = 9'b111111111;
assign micromatrizz[55][118] = 9'b111111111;
assign micromatrizz[55][119] = 9'b111111111;
assign micromatrizz[55][120] = 9'b111111111;
assign micromatrizz[55][121] = 9'b111110010;
assign micromatrizz[55][122] = 9'b111110010;
assign micromatrizz[55][123] = 9'b111110011;
assign micromatrizz[55][124] = 9'b111110011;
assign micromatrizz[55][125] = 9'b111110010;
assign micromatrizz[55][126] = 9'b111110111;
assign micromatrizz[55][127] = 9'b111111111;
assign micromatrizz[55][128] = 9'b111111111;
assign micromatrizz[55][129] = 9'b111111111;
assign micromatrizz[55][130] = 9'b111111111;
assign micromatrizz[55][131] = 9'b111111111;
assign micromatrizz[55][132] = 9'b111111111;
assign micromatrizz[55][133] = 9'b111110110;
assign micromatrizz[55][134] = 9'b111111111;
assign micromatrizz[55][135] = 9'b111111111;
assign micromatrizz[55][136] = 9'b111111111;
assign micromatrizz[55][137] = 9'b111111111;
assign micromatrizz[55][138] = 9'b111110111;
assign micromatrizz[55][139] = 9'b111110010;
assign micromatrizz[55][140] = 9'b111110010;
assign micromatrizz[55][141] = 9'b111110010;
assign micromatrizz[55][142] = 9'b111110010;
assign micromatrizz[55][143] = 9'b111110011;
assign micromatrizz[55][144] = 9'b111110011;
assign micromatrizz[55][145] = 9'b111110011;
assign micromatrizz[55][146] = 9'b111111111;
assign micromatrizz[55][147] = 9'b111111111;
assign micromatrizz[55][148] = 9'b111111111;
assign micromatrizz[55][149] = 9'b111111111;
assign micromatrizz[55][150] = 9'b111110111;
assign micromatrizz[55][151] = 9'b111110010;
assign micromatrizz[55][152] = 9'b111110011;
assign micromatrizz[55][153] = 9'b111110011;
assign micromatrizz[55][154] = 9'b111110011;
assign micromatrizz[55][155] = 9'b111110011;
assign micromatrizz[55][156] = 9'b111110010;
assign micromatrizz[55][157] = 9'b111110111;
assign micromatrizz[55][158] = 9'b111111111;
assign micromatrizz[55][159] = 9'b111111111;
assign micromatrizz[55][160] = 9'b111111111;
assign micromatrizz[55][161] = 9'b111111111;
assign micromatrizz[55][162] = 9'b111111111;
assign micromatrizz[55][163] = 9'b111111111;
assign micromatrizz[55][164] = 9'b111111111;
assign micromatrizz[55][165] = 9'b111111111;
assign micromatrizz[55][166] = 9'b111111111;
assign micromatrizz[55][167] = 9'b111111111;
assign micromatrizz[55][168] = 9'b111111111;
assign micromatrizz[55][169] = 9'b111111111;
assign micromatrizz[55][170] = 9'b111111111;
assign micromatrizz[55][171] = 9'b111111111;
assign micromatrizz[55][172] = 9'b111110010;
assign micromatrizz[55][173] = 9'b111110010;
assign micromatrizz[55][174] = 9'b111110011;
assign micromatrizz[55][175] = 9'b111110010;
assign micromatrizz[55][176] = 9'b111110011;
assign micromatrizz[55][177] = 9'b111110011;
assign micromatrizz[55][178] = 9'b111110011;
assign micromatrizz[55][179] = 9'b111111111;
assign micromatrizz[55][180] = 9'b111111111;
assign micromatrizz[55][181] = 9'b111111111;
assign micromatrizz[55][182] = 9'b111111111;
assign micromatrizz[55][183] = 9'b111111111;
assign micromatrizz[55][184] = 9'b111110110;
assign micromatrizz[55][185] = 9'b111110010;
assign micromatrizz[55][186] = 9'b111110010;
assign micromatrizz[55][187] = 9'b111110011;
assign micromatrizz[55][188] = 9'b111110011;
assign micromatrizz[55][189] = 9'b111110011;
assign micromatrizz[55][190] = 9'b111110111;
assign micromatrizz[55][191] = 9'b111111111;
assign micromatrizz[55][192] = 9'b111111111;
assign micromatrizz[55][193] = 9'b111111111;
assign micromatrizz[55][194] = 9'b111110110;
assign micromatrizz[55][195] = 9'b111110010;
assign micromatrizz[55][196] = 9'b111110011;
assign micromatrizz[55][197] = 9'b111110011;
assign micromatrizz[55][198] = 9'b111110011;
assign micromatrizz[55][199] = 9'b111110010;
assign micromatrizz[55][200] = 9'b111110010;
assign micromatrizz[55][201] = 9'b111110011;
assign micromatrizz[55][202] = 9'b111110111;
assign micromatrizz[55][203] = 9'b111111111;
assign micromatrizz[55][204] = 9'b111111111;
assign micromatrizz[55][205] = 9'b111111111;
assign micromatrizz[55][206] = 9'b111111111;
assign micromatrizz[55][207] = 9'b111110111;
assign micromatrizz[55][208] = 9'b111110010;
assign micromatrizz[55][209] = 9'b111110011;
assign micromatrizz[55][210] = 9'b111110011;
assign micromatrizz[55][211] = 9'b111110011;
assign micromatrizz[55][212] = 9'b111110011;
assign micromatrizz[55][213] = 9'b111110111;
assign micromatrizz[55][214] = 9'b111111111;
assign micromatrizz[55][215] = 9'b111111111;
assign micromatrizz[55][216] = 9'b111111111;
assign micromatrizz[55][217] = 9'b111111111;
assign micromatrizz[55][218] = 9'b111111111;
assign micromatrizz[55][219] = 9'b111110111;
assign micromatrizz[55][220] = 9'b111111111;
assign micromatrizz[55][221] = 9'b111111111;
assign micromatrizz[55][222] = 9'b111111111;
assign micromatrizz[55][223] = 9'b111111111;
assign micromatrizz[55][224] = 9'b111111111;
assign micromatrizz[55][225] = 9'b111110111;
assign micromatrizz[55][226] = 9'b111110010;
assign micromatrizz[55][227] = 9'b111110010;
assign micromatrizz[55][228] = 9'b111110010;
assign micromatrizz[55][229] = 9'b111110011;
assign micromatrizz[55][230] = 9'b111110011;
assign micromatrizz[55][231] = 9'b111110011;
assign micromatrizz[55][232] = 9'b111110011;
assign micromatrizz[55][233] = 9'b111110011;
assign micromatrizz[55][234] = 9'b111111111;
assign micromatrizz[55][235] = 9'b111111111;
assign micromatrizz[55][236] = 9'b111111111;
assign micromatrizz[55][237] = 9'b111111111;
assign micromatrizz[55][238] = 9'b111111111;
assign micromatrizz[55][239] = 9'b111111111;
assign micromatrizz[55][240] = 9'b111111111;
assign micromatrizz[55][241] = 9'b111111111;
assign micromatrizz[55][242] = 9'b111110111;
assign micromatrizz[55][243] = 9'b111110010;
assign micromatrizz[55][244] = 9'b111110011;
assign micromatrizz[55][245] = 9'b111110011;
assign micromatrizz[55][246] = 9'b111110010;
assign micromatrizz[55][247] = 9'b111110111;
assign micromatrizz[55][248] = 9'b111111111;
assign micromatrizz[55][249] = 9'b111111111;
assign micromatrizz[55][250] = 9'b111111111;
assign micromatrizz[55][251] = 9'b111110111;
assign micromatrizz[55][252] = 9'b111110010;
assign micromatrizz[55][253] = 9'b111110010;
assign micromatrizz[55][254] = 9'b111110011;
assign micromatrizz[55][255] = 9'b111110111;
assign micromatrizz[55][256] = 9'b111111111;
assign micromatrizz[55][257] = 9'b111111111;
assign micromatrizz[55][258] = 9'b111111111;
assign micromatrizz[55][259] = 9'b111111111;
assign micromatrizz[55][260] = 9'b111110010;
assign micromatrizz[55][261] = 9'b111110010;
assign micromatrizz[55][262] = 9'b111110011;
assign micromatrizz[55][263] = 9'b111110011;
assign micromatrizz[55][264] = 9'b111110011;
assign micromatrizz[55][265] = 9'b111110011;
assign micromatrizz[55][266] = 9'b111111111;
assign micromatrizz[55][267] = 9'b111111111;
assign micromatrizz[55][268] = 9'b111111111;
assign micromatrizz[55][269] = 9'b111111111;
assign micromatrizz[55][270] = 9'b111111111;
assign micromatrizz[55][271] = 9'b111111111;
assign micromatrizz[55][272] = 9'b111111111;
assign micromatrizz[55][273] = 9'b111111111;
assign micromatrizz[55][274] = 9'b111111111;
assign micromatrizz[55][275] = 9'b111111111;
assign micromatrizz[55][276] = 9'b111111111;
assign micromatrizz[55][277] = 9'b111111111;
assign micromatrizz[55][278] = 9'b111111111;
assign micromatrizz[55][279] = 9'b111111111;
assign micromatrizz[55][280] = 9'b111111111;
assign micromatrizz[55][281] = 9'b111111111;
assign micromatrizz[55][282] = 9'b111111111;
assign micromatrizz[55][283] = 9'b111111111;
assign micromatrizz[55][284] = 9'b111111111;
assign micromatrizz[55][285] = 9'b111111111;
assign micromatrizz[55][286] = 9'b111110010;
assign micromatrizz[55][287] = 9'b111110010;
assign micromatrizz[55][288] = 9'b111110011;
assign micromatrizz[55][289] = 9'b111110011;
assign micromatrizz[55][290] = 9'b111110011;
assign micromatrizz[55][291] = 9'b111110011;
assign micromatrizz[55][292] = 9'b111110010;
assign micromatrizz[55][293] = 9'b111111111;
assign micromatrizz[55][294] = 9'b111111111;
assign micromatrizz[55][295] = 9'b111111111;
assign micromatrizz[55][296] = 9'b111111111;
assign micromatrizz[55][297] = 9'b111110010;
assign micromatrizz[55][298] = 9'b111110010;
assign micromatrizz[55][299] = 9'b111110011;
assign micromatrizz[55][300] = 9'b111110011;
assign micromatrizz[55][301] = 9'b111110011;
assign micromatrizz[55][302] = 9'b111110010;
assign micromatrizz[55][303] = 9'b111110011;
assign micromatrizz[55][304] = 9'b111110011;
assign micromatrizz[55][305] = 9'b111110011;
assign micromatrizz[55][306] = 9'b111111111;
assign micromatrizz[55][307] = 9'b111111111;
assign micromatrizz[55][308] = 9'b111111111;
assign micromatrizz[55][309] = 9'b111111111;
assign micromatrizz[55][310] = 9'b111111111;
assign micromatrizz[55][311] = 9'b111111111;
assign micromatrizz[55][312] = 9'b111110010;
assign micromatrizz[55][313] = 9'b111111111;
assign micromatrizz[55][314] = 9'b111111111;
assign micromatrizz[55][315] = 9'b111111111;
assign micromatrizz[55][316] = 9'b111111111;
assign micromatrizz[55][317] = 9'b111110110;
assign micromatrizz[55][318] = 9'b111110010;
assign micromatrizz[55][319] = 9'b111110010;
assign micromatrizz[55][320] = 9'b111110010;
assign micromatrizz[55][321] = 9'b111110010;
assign micromatrizz[55][322] = 9'b111111111;
assign micromatrizz[55][323] = 9'b111111111;
assign micromatrizz[55][324] = 9'b111111111;
assign micromatrizz[55][325] = 9'b111111111;
assign micromatrizz[55][326] = 9'b111110010;
assign micromatrizz[55][327] = 9'b111110010;
assign micromatrizz[55][328] = 9'b111110010;
assign micromatrizz[55][329] = 9'b111110010;
assign micromatrizz[55][330] = 9'b111111111;
assign micromatrizz[55][331] = 9'b111111111;
assign micromatrizz[55][332] = 9'b111111111;
assign micromatrizz[55][333] = 9'b111111111;
assign micromatrizz[55][334] = 9'b111111111;
assign micromatrizz[55][335] = 9'b111110010;
assign micromatrizz[55][336] = 9'b111110010;
assign micromatrizz[55][337] = 9'b111110010;
assign micromatrizz[55][338] = 9'b111110011;
assign micromatrizz[55][339] = 9'b111110011;
assign micromatrizz[55][340] = 9'b111110011;
assign micromatrizz[55][341] = 9'b111110011;
assign micromatrizz[55][342] = 9'b111110111;
assign micromatrizz[55][343] = 9'b111111111;
assign micromatrizz[55][344] = 9'b111111111;
assign micromatrizz[55][345] = 9'b111111111;
assign micromatrizz[55][346] = 9'b111111111;
assign micromatrizz[55][347] = 9'b111110010;
assign micromatrizz[55][348] = 9'b111110010;
assign micromatrizz[55][349] = 9'b111110011;
assign micromatrizz[55][350] = 9'b111110011;
assign micromatrizz[55][351] = 9'b111110011;
assign micromatrizz[55][352] = 9'b111110011;
assign micromatrizz[55][353] = 9'b111110011;
assign micromatrizz[55][354] = 9'b111111111;
assign micromatrizz[55][355] = 9'b111111111;
assign micromatrizz[55][356] = 9'b111111111;
assign micromatrizz[55][357] = 9'b111111111;
assign micromatrizz[55][358] = 9'b111111111;
assign micromatrizz[55][359] = 9'b111110010;
assign micromatrizz[55][360] = 9'b111110011;
assign micromatrizz[55][361] = 9'b111110010;
assign micromatrizz[55][362] = 9'b111110010;
assign micromatrizz[55][363] = 9'b111110011;
assign micromatrizz[55][364] = 9'b111110011;
assign micromatrizz[55][365] = 9'b111110011;
assign micromatrizz[55][366] = 9'b111111111;
assign micromatrizz[55][367] = 9'b111111111;
assign micromatrizz[55][368] = 9'b111111111;
assign micromatrizz[55][369] = 9'b111111111;
assign micromatrizz[55][370] = 9'b111111111;
assign micromatrizz[55][371] = 9'b111111111;
assign micromatrizz[55][372] = 9'b111110010;
assign micromatrizz[55][373] = 9'b111110011;
assign micromatrizz[55][374] = 9'b111110011;
assign micromatrizz[55][375] = 9'b111110011;
assign micromatrizz[55][376] = 9'b111110011;
assign micromatrizz[55][377] = 9'b111110011;
assign micromatrizz[55][378] = 9'b111110010;
assign micromatrizz[55][379] = 9'b111111111;
assign micromatrizz[55][380] = 9'b111111111;
assign micromatrizz[55][381] = 9'b111111111;
assign micromatrizz[55][382] = 9'b111111111;
assign micromatrizz[55][383] = 9'b111110111;
assign micromatrizz[55][384] = 9'b111110010;
assign micromatrizz[55][385] = 9'b111110010;
assign micromatrizz[55][386] = 9'b111110011;
assign micromatrizz[55][387] = 9'b111110011;
assign micromatrizz[55][388] = 9'b111110011;
assign micromatrizz[55][389] = 9'b111110011;
assign micromatrizz[55][390] = 9'b111110011;
assign micromatrizz[55][391] = 9'b111111111;
assign micromatrizz[55][392] = 9'b111111111;
assign micromatrizz[55][393] = 9'b111111111;
assign micromatrizz[55][394] = 9'b111111111;
assign micromatrizz[55][395] = 9'b111110010;
assign micromatrizz[55][396] = 9'b111110010;
assign micromatrizz[55][397] = 9'b111110010;
assign micromatrizz[55][398] = 9'b111110011;
assign micromatrizz[55][399] = 9'b111110011;
assign micromatrizz[55][400] = 9'b111110011;
assign micromatrizz[55][401] = 9'b111110011;
assign micromatrizz[55][402] = 9'b111110011;
assign micromatrizz[55][403] = 9'b111110111;
assign micromatrizz[55][404] = 9'b111111111;
assign micromatrizz[55][405] = 9'b111111111;
assign micromatrizz[55][406] = 9'b111111111;
assign micromatrizz[55][407] = 9'b111111111;
assign micromatrizz[55][408] = 9'b111111111;
assign micromatrizz[55][409] = 9'b111111111;
assign micromatrizz[55][410] = 9'b111111111;
assign micromatrizz[55][411] = 9'b111111111;
assign micromatrizz[55][412] = 9'b111111111;
assign micromatrizz[55][413] = 9'b111110010;
assign micromatrizz[55][414] = 9'b111110011;
assign micromatrizz[55][415] = 9'b111110011;
assign micromatrizz[55][416] = 9'b111110010;
assign micromatrizz[55][417] = 9'b111110111;
assign micromatrizz[55][418] = 9'b111111111;
assign micromatrizz[55][419] = 9'b111111111;
assign micromatrizz[55][420] = 9'b111111111;
assign micromatrizz[55][421] = 9'b111110111;
assign micromatrizz[55][422] = 9'b111110010;
assign micromatrizz[55][423] = 9'b111110010;
assign micromatrizz[55][424] = 9'b111110011;
assign micromatrizz[55][425] = 9'b111110111;
assign micromatrizz[55][426] = 9'b111111111;
assign micromatrizz[55][427] = 9'b111111111;
assign micromatrizz[55][428] = 9'b111111111;
assign micromatrizz[55][429] = 9'b111111111;
assign micromatrizz[55][430] = 9'b111110111;
assign micromatrizz[55][431] = 9'b111110010;
assign micromatrizz[55][432] = 9'b111110010;
assign micromatrizz[55][433] = 9'b111110010;
assign micromatrizz[55][434] = 9'b111110011;
assign micromatrizz[55][435] = 9'b111110011;
assign micromatrizz[55][436] = 9'b111110011;
assign micromatrizz[55][437] = 9'b111110011;
assign micromatrizz[55][438] = 9'b111110011;
assign micromatrizz[55][439] = 9'b111111111;
assign micromatrizz[55][440] = 9'b111111111;
assign micromatrizz[55][441] = 9'b111111111;
assign micromatrizz[55][442] = 9'b111111111;
assign micromatrizz[55][443] = 9'b111111111;
assign micromatrizz[55][444] = 9'b111111111;
assign micromatrizz[55][445] = 9'b111111111;
assign micromatrizz[55][446] = 9'b111111111;
assign micromatrizz[55][447] = 9'b111111111;
assign micromatrizz[55][448] = 9'b111110010;
assign micromatrizz[55][449] = 9'b111110010;
assign micromatrizz[55][450] = 9'b111110011;
assign micromatrizz[55][451] = 9'b111110011;
assign micromatrizz[55][452] = 9'b111110010;
assign micromatrizz[55][453] = 9'b111110011;
assign micromatrizz[55][454] = 9'b111111111;
assign micromatrizz[55][455] = 9'b111111111;
assign micromatrizz[55][456] = 9'b111111111;
assign micromatrizz[55][457] = 9'b111111111;
assign micromatrizz[55][458] = 9'b111111111;
assign micromatrizz[55][459] = 9'b111111111;
assign micromatrizz[55][460] = 9'b111110110;
assign micromatrizz[55][461] = 9'b111111111;
assign micromatrizz[55][462] = 9'b111111111;
assign micromatrizz[55][463] = 9'b111111111;
assign micromatrizz[55][464] = 9'b111111111;
assign micromatrizz[55][465] = 9'b111110111;
assign micromatrizz[55][466] = 9'b111110010;
assign micromatrizz[55][467] = 9'b111110011;
assign micromatrizz[55][468] = 9'b111110011;
assign micromatrizz[55][469] = 9'b111110011;
assign micromatrizz[55][470] = 9'b111110010;
assign micromatrizz[55][471] = 9'b111111111;
assign micromatrizz[55][472] = 9'b111111111;
assign micromatrizz[55][473] = 9'b111111111;
assign micromatrizz[55][474] = 9'b111111111;
assign micromatrizz[55][475] = 9'b111111111;
assign micromatrizz[55][476] = 9'b111111111;
assign micromatrizz[55][477] = 9'b111111111;
assign micromatrizz[55][478] = 9'b111111111;
assign micromatrizz[55][479] = 9'b111111111;
assign micromatrizz[55][480] = 9'b111111111;
assign micromatrizz[55][481] = 9'b111110010;
assign micromatrizz[55][482] = 9'b111110010;
assign micromatrizz[55][483] = 9'b111110010;
assign micromatrizz[55][484] = 9'b111110010;
assign micromatrizz[55][485] = 9'b111110011;
assign micromatrizz[55][486] = 9'b111110011;
assign micromatrizz[55][487] = 9'b111110011;
assign micromatrizz[55][488] = 9'b111110010;
assign micromatrizz[55][489] = 9'b111110111;
assign micromatrizz[55][490] = 9'b111111111;
assign micromatrizz[55][491] = 9'b111111111;
assign micromatrizz[55][492] = 9'b111111111;
assign micromatrizz[55][493] = 9'b111111111;
assign micromatrizz[55][494] = 9'b111111111;
assign micromatrizz[55][495] = 9'b111111111;
assign micromatrizz[55][496] = 9'b111111111;
assign micromatrizz[55][497] = 9'b111111111;
assign micromatrizz[55][498] = 9'b111110111;
assign micromatrizz[55][499] = 9'b111110010;
assign micromatrizz[55][500] = 9'b111110011;
assign micromatrizz[55][501] = 9'b111110011;
assign micromatrizz[55][502] = 9'b111110010;
assign micromatrizz[55][503] = 9'b111110111;
assign micromatrizz[55][504] = 9'b111111111;
assign micromatrizz[55][505] = 9'b111111111;
assign micromatrizz[55][506] = 9'b111111111;
assign micromatrizz[55][507] = 9'b111110010;
assign micromatrizz[55][508] = 9'b111110010;
assign micromatrizz[55][509] = 9'b111110011;
assign micromatrizz[55][510] = 9'b111110011;
assign micromatrizz[55][511] = 9'b111110111;
assign micromatrizz[55][512] = 9'b111111111;
assign micromatrizz[55][513] = 9'b111111111;
assign micromatrizz[55][514] = 9'b111111111;
assign micromatrizz[55][515] = 9'b111111111;
assign micromatrizz[55][516] = 9'b111110111;
assign micromatrizz[55][517] = 9'b111110010;
assign micromatrizz[55][518] = 9'b111110011;
assign micromatrizz[55][519] = 9'b111110011;
assign micromatrizz[55][520] = 9'b111110010;
assign micromatrizz[55][521] = 9'b111110010;
assign micromatrizz[55][522] = 9'b111110011;
assign micromatrizz[55][523] = 9'b111110011;
assign micromatrizz[55][524] = 9'b111110111;
assign micromatrizz[55][525] = 9'b111111111;
assign micromatrizz[55][526] = 9'b111111111;
assign micromatrizz[55][527] = 9'b111111111;
assign micromatrizz[55][528] = 9'b111110111;
assign micromatrizz[55][529] = 9'b111110010;
assign micromatrizz[55][530] = 9'b111110011;
assign micromatrizz[55][531] = 9'b111110011;
assign micromatrizz[55][532] = 9'b111110011;
assign micromatrizz[55][533] = 9'b111110010;
assign micromatrizz[55][534] = 9'b111110011;
assign micromatrizz[55][535] = 9'b111111111;
assign micromatrizz[55][536] = 9'b111111111;
assign micromatrizz[55][537] = 9'b111111111;
assign micromatrizz[55][538] = 9'b111111111;
assign micromatrizz[55][539] = 9'b111111111;
assign micromatrizz[55][540] = 9'b111110111;
assign micromatrizz[55][541] = 9'b111110010;
assign micromatrizz[55][542] = 9'b111110010;
assign micromatrizz[55][543] = 9'b111110011;
assign micromatrizz[55][544] = 9'b111110010;
assign micromatrizz[55][545] = 9'b111111111;
assign micromatrizz[55][546] = 9'b111111111;
assign micromatrizz[55][547] = 9'b111111111;
assign micromatrizz[55][548] = 9'b111111111;
assign micromatrizz[55][549] = 9'b111110010;
assign micromatrizz[55][550] = 9'b111110011;
assign micromatrizz[55][551] = 9'b111110011;
assign micromatrizz[55][552] = 9'b111110010;
assign micromatrizz[55][553] = 9'b111111111;
assign micromatrizz[55][554] = 9'b111111111;
assign micromatrizz[55][555] = 9'b111111111;
assign micromatrizz[55][556] = 9'b111111111;
assign micromatrizz[55][557] = 9'b111111111;
assign micromatrizz[55][558] = 9'b111110010;
assign micromatrizz[55][559] = 9'b111110010;
assign micromatrizz[55][560] = 9'b111110010;
assign micromatrizz[55][561] = 9'b111110010;
assign micromatrizz[55][562] = 9'b111110011;
assign micromatrizz[55][563] = 9'b111110011;
assign micromatrizz[55][564] = 9'b111110011;
assign micromatrizz[55][565] = 9'b111111111;
assign micromatrizz[55][566] = 9'b111111111;
assign micromatrizz[55][567] = 9'b111111111;
assign micromatrizz[55][568] = 9'b111111111;
assign micromatrizz[55][569] = 9'b111111111;
assign micromatrizz[55][570] = 9'b111110010;
assign micromatrizz[55][571] = 9'b111110010;
assign micromatrizz[55][572] = 9'b111110011;
assign micromatrizz[55][573] = 9'b111110010;
assign micromatrizz[55][574] = 9'b111110010;
assign micromatrizz[55][575] = 9'b111110011;
assign micromatrizz[55][576] = 9'b111111111;
assign micromatrizz[55][577] = 9'b111111111;
assign micromatrizz[55][578] = 9'b111111111;
assign micromatrizz[55][579] = 9'b111111111;
assign micromatrizz[55][580] = 9'b111110110;
assign micromatrizz[55][581] = 9'b111110010;
assign micromatrizz[55][582] = 9'b111110010;
assign micromatrizz[55][583] = 9'b111110011;
assign micromatrizz[55][584] = 9'b111110010;
assign micromatrizz[55][585] = 9'b111110010;
assign micromatrizz[55][586] = 9'b111110011;
assign micromatrizz[55][587] = 9'b111110011;
assign micromatrizz[55][588] = 9'b111111111;
assign micromatrizz[55][589] = 9'b111111111;
assign micromatrizz[55][590] = 9'b111111111;
assign micromatrizz[55][591] = 9'b111111111;
assign micromatrizz[55][592] = 9'b111111111;
assign micromatrizz[55][593] = 9'b111110010;
assign micromatrizz[55][594] = 9'b111110010;
assign micromatrizz[55][595] = 9'b111110011;
assign micromatrizz[55][596] = 9'b111110011;
assign micromatrizz[55][597] = 9'b111110010;
assign micromatrizz[55][598] = 9'b111111111;
assign micromatrizz[55][599] = 9'b111111111;
assign micromatrizz[55][600] = 9'b111111111;
assign micromatrizz[55][601] = 9'b111111111;
assign micromatrizz[55][602] = 9'b111110010;
assign micromatrizz[55][603] = 9'b111110011;
assign micromatrizz[55][604] = 9'b111110011;
assign micromatrizz[55][605] = 9'b111110010;
assign micromatrizz[55][606] = 9'b111111111;
assign micromatrizz[55][607] = 9'b111111111;
assign micromatrizz[55][608] = 9'b111111111;
assign micromatrizz[55][609] = 9'b111111111;
assign micromatrizz[55][610] = 9'b111110111;
assign micromatrizz[55][611] = 9'b111110010;
assign micromatrizz[55][612] = 9'b111110011;
assign micromatrizz[55][613] = 9'b111110010;
assign micromatrizz[55][614] = 9'b111110011;
assign micromatrizz[55][615] = 9'b111110010;
assign micromatrizz[55][616] = 9'b111110111;
assign micromatrizz[55][617] = 9'b111111111;
assign micromatrizz[55][618] = 9'b111111111;
assign micromatrizz[55][619] = 9'b111111111;
assign micromatrizz[55][620] = 9'b111111111;
assign micromatrizz[55][621] = 9'b111111111;
assign micromatrizz[55][622] = 9'b111111111;
assign micromatrizz[55][623] = 9'b111111111;
assign micromatrizz[55][624] = 9'b111111111;
assign micromatrizz[55][625] = 9'b111111111;
assign micromatrizz[55][626] = 9'b111111111;
assign micromatrizz[55][627] = 9'b111111111;
assign micromatrizz[55][628] = 9'b111111111;
assign micromatrizz[55][629] = 9'b111111111;
assign micromatrizz[55][630] = 9'b111111111;
assign micromatrizz[55][631] = 9'b111111111;
assign micromatrizz[55][632] = 9'b111111111;
assign micromatrizz[55][633] = 9'b111111111;
assign micromatrizz[55][634] = 9'b111111111;
assign micromatrizz[55][635] = 9'b111111111;
assign micromatrizz[55][636] = 9'b111111111;
assign micromatrizz[55][637] = 9'b111111111;
assign micromatrizz[55][638] = 9'b111111111;
assign micromatrizz[55][639] = 9'b111111111;
assign micromatrizz[56][0] = 9'b111111111;
assign micromatrizz[56][1] = 9'b111111111;
assign micromatrizz[56][2] = 9'b111111111;
assign micromatrizz[56][3] = 9'b111111111;
assign micromatrizz[56][4] = 9'b111111111;
assign micromatrizz[56][5] = 9'b111111111;
assign micromatrizz[56][6] = 9'b111111111;
assign micromatrizz[56][7] = 9'b111111111;
assign micromatrizz[56][8] = 9'b111110010;
assign micromatrizz[56][9] = 9'b111110011;
assign micromatrizz[56][10] = 9'b111110010;
assign micromatrizz[56][11] = 9'b111110010;
assign micromatrizz[56][12] = 9'b111110011;
assign micromatrizz[56][13] = 9'b111110011;
assign micromatrizz[56][14] = 9'b111110011;
assign micromatrizz[56][15] = 9'b111111111;
assign micromatrizz[56][16] = 9'b111111111;
assign micromatrizz[56][17] = 9'b111111111;
assign micromatrizz[56][18] = 9'b111111111;
assign micromatrizz[56][19] = 9'b111111111;
assign micromatrizz[56][20] = 9'b111111111;
assign micromatrizz[56][21] = 9'b111111111;
assign micromatrizz[56][22] = 9'b111111111;
assign micromatrizz[56][23] = 9'b111111111;
assign micromatrizz[56][24] = 9'b111110010;
assign micromatrizz[56][25] = 9'b111110010;
assign micromatrizz[56][26] = 9'b111110010;
assign micromatrizz[56][27] = 9'b111110011;
assign micromatrizz[56][28] = 9'b111110011;
assign micromatrizz[56][29] = 9'b111110011;
assign micromatrizz[56][30] = 9'b111110011;
assign micromatrizz[56][31] = 9'b111111111;
assign micromatrizz[56][32] = 9'b111111111;
assign micromatrizz[56][33] = 9'b111111111;
assign micromatrizz[56][34] = 9'b111111111;
assign micromatrizz[56][35] = 9'b111110111;
assign micromatrizz[56][36] = 9'b111110010;
assign micromatrizz[56][37] = 9'b111110010;
assign micromatrizz[56][38] = 9'b111110010;
assign micromatrizz[56][39] = 9'b111110011;
assign micromatrizz[56][40] = 9'b111110011;
assign micromatrizz[56][41] = 9'b111110011;
assign micromatrizz[56][42] = 9'b111110011;
assign micromatrizz[56][43] = 9'b111111111;
assign micromatrizz[56][44] = 9'b111111111;
assign micromatrizz[56][45] = 9'b111111111;
assign micromatrizz[56][46] = 9'b111111111;
assign micromatrizz[56][47] = 9'b111110010;
assign micromatrizz[56][48] = 9'b111110010;
assign micromatrizz[56][49] = 9'b111110010;
assign micromatrizz[56][50] = 9'b111110011;
assign micromatrizz[56][51] = 9'b111110011;
assign micromatrizz[56][52] = 9'b111110011;
assign micromatrizz[56][53] = 9'b111110010;
assign micromatrizz[56][54] = 9'b111110111;
assign micromatrizz[56][55] = 9'b111111111;
assign micromatrizz[56][56] = 9'b111111111;
assign micromatrizz[56][57] = 9'b111111111;
assign micromatrizz[56][58] = 9'b111111111;
assign micromatrizz[56][59] = 9'b111110010;
assign micromatrizz[56][60] = 9'b111110010;
assign micromatrizz[56][61] = 9'b111110010;
assign micromatrizz[56][62] = 9'b111110010;
assign micromatrizz[56][63] = 9'b111110011;
assign micromatrizz[56][64] = 9'b111110011;
assign micromatrizz[56][65] = 9'b111110011;
assign micromatrizz[56][66] = 9'b111111111;
assign micromatrizz[56][67] = 9'b111111111;
assign micromatrizz[56][68] = 9'b111111111;
assign micromatrizz[56][69] = 9'b111110111;
assign micromatrizz[56][70] = 9'b111110010;
assign micromatrizz[56][71] = 9'b111110010;
assign micromatrizz[56][72] = 9'b111110011;
assign micromatrizz[56][73] = 9'b111110011;
assign micromatrizz[56][74] = 9'b111110010;
assign micromatrizz[56][75] = 9'b111111111;
assign micromatrizz[56][76] = 9'b111111111;
assign micromatrizz[56][77] = 9'b111111111;
assign micromatrizz[56][78] = 9'b111111111;
assign micromatrizz[56][79] = 9'b111110010;
assign micromatrizz[56][80] = 9'b111110010;
assign micromatrizz[56][81] = 9'b111110011;
assign micromatrizz[56][82] = 9'b111110011;
assign micromatrizz[56][83] = 9'b111110011;
assign micromatrizz[56][84] = 9'b111111111;
assign micromatrizz[56][85] = 9'b111111111;
assign micromatrizz[56][86] = 9'b111111111;
assign micromatrizz[56][87] = 9'b111111111;
assign micromatrizz[56][88] = 9'b111110110;
assign micromatrizz[56][89] = 9'b111110010;
assign micromatrizz[56][90] = 9'b111110010;
assign micromatrizz[56][91] = 9'b111110010;
assign micromatrizz[56][92] = 9'b111110011;
assign micromatrizz[56][93] = 9'b111110011;
assign micromatrizz[56][94] = 9'b111110011;
assign micromatrizz[56][95] = 9'b111110011;
assign micromatrizz[56][96] = 9'b111111111;
assign micromatrizz[56][97] = 9'b111111111;
assign micromatrizz[56][98] = 9'b111111111;
assign micromatrizz[56][99] = 9'b111111111;
assign micromatrizz[56][100] = 9'b111111111;
assign micromatrizz[56][101] = 9'b111111111;
assign micromatrizz[56][102] = 9'b111111111;
assign micromatrizz[56][103] = 9'b111111111;
assign micromatrizz[56][104] = 9'b111110010;
assign micromatrizz[56][105] = 9'b111110010;
assign micromatrizz[56][106] = 9'b111110010;
assign micromatrizz[56][107] = 9'b111110010;
assign micromatrizz[56][108] = 9'b111110011;
assign micromatrizz[56][109] = 9'b111110011;
assign micromatrizz[56][110] = 9'b111110010;
assign micromatrizz[56][111] = 9'b111111111;
assign micromatrizz[56][112] = 9'b111111111;
assign micromatrizz[56][113] = 9'b111111111;
assign micromatrizz[56][114] = 9'b111111111;
assign micromatrizz[56][115] = 9'b111111111;
assign micromatrizz[56][116] = 9'b111111111;
assign micromatrizz[56][117] = 9'b111111111;
assign micromatrizz[56][118] = 9'b111111111;
assign micromatrizz[56][119] = 9'b111111111;
assign micromatrizz[56][120] = 9'b111110010;
assign micromatrizz[56][121] = 9'b111110010;
assign micromatrizz[56][122] = 9'b111110010;
assign micromatrizz[56][123] = 9'b111110010;
assign micromatrizz[56][124] = 9'b111110011;
assign micromatrizz[56][125] = 9'b111110011;
assign micromatrizz[56][126] = 9'b111110111;
assign micromatrizz[56][127] = 9'b111111111;
assign micromatrizz[56][128] = 9'b111111111;
assign micromatrizz[56][129] = 9'b111111111;
assign micromatrizz[56][130] = 9'b111111111;
assign micromatrizz[56][131] = 9'b111111111;
assign micromatrizz[56][132] = 9'b111111111;
assign micromatrizz[56][133] = 9'b111110111;
assign micromatrizz[56][134] = 9'b111110111;
assign micromatrizz[56][135] = 9'b111111111;
assign micromatrizz[56][136] = 9'b111111111;
assign micromatrizz[56][137] = 9'b111111111;
assign micromatrizz[56][138] = 9'b111110111;
assign micromatrizz[56][139] = 9'b111110010;
assign micromatrizz[56][140] = 9'b111110010;
assign micromatrizz[56][141] = 9'b111110010;
assign micromatrizz[56][142] = 9'b111110011;
assign micromatrizz[56][143] = 9'b111110011;
assign micromatrizz[56][144] = 9'b111110011;
assign micromatrizz[56][145] = 9'b111110011;
assign micromatrizz[56][146] = 9'b111111111;
assign micromatrizz[56][147] = 9'b111111111;
assign micromatrizz[56][148] = 9'b111111111;
assign micromatrizz[56][149] = 9'b111111111;
assign micromatrizz[56][150] = 9'b111110111;
assign micromatrizz[56][151] = 9'b111110010;
assign micromatrizz[56][152] = 9'b111110011;
assign micromatrizz[56][153] = 9'b111110011;
assign micromatrizz[56][154] = 9'b111110011;
assign micromatrizz[56][155] = 9'b111110010;
assign micromatrizz[56][156] = 9'b111110011;
assign micromatrizz[56][157] = 9'b111110111;
assign micromatrizz[56][158] = 9'b111111111;
assign micromatrizz[56][159] = 9'b111111111;
assign micromatrizz[56][160] = 9'b111111111;
assign micromatrizz[56][161] = 9'b111111111;
assign micromatrizz[56][162] = 9'b111111111;
assign micromatrizz[56][163] = 9'b111111111;
assign micromatrizz[56][164] = 9'b111111111;
assign micromatrizz[56][165] = 9'b111111111;
assign micromatrizz[56][166] = 9'b111111111;
assign micromatrizz[56][167] = 9'b111111111;
assign micromatrizz[56][168] = 9'b111111111;
assign micromatrizz[56][169] = 9'b111111111;
assign micromatrizz[56][170] = 9'b111111111;
assign micromatrizz[56][171] = 9'b111111111;
assign micromatrizz[56][172] = 9'b111110010;
assign micromatrizz[56][173] = 9'b111110010;
assign micromatrizz[56][174] = 9'b111110011;
assign micromatrizz[56][175] = 9'b111110010;
assign micromatrizz[56][176] = 9'b111110011;
assign micromatrizz[56][177] = 9'b111110011;
assign micromatrizz[56][178] = 9'b111110011;
assign micromatrizz[56][179] = 9'b111110111;
assign micromatrizz[56][180] = 9'b111111111;
assign micromatrizz[56][181] = 9'b111111111;
assign micromatrizz[56][182] = 9'b111111111;
assign micromatrizz[56][183] = 9'b111110111;
assign micromatrizz[56][184] = 9'b111110010;
assign micromatrizz[56][185] = 9'b111110010;
assign micromatrizz[56][186] = 9'b111110010;
assign micromatrizz[56][187] = 9'b111110010;
assign micromatrizz[56][188] = 9'b111110011;
assign micromatrizz[56][189] = 9'b111110011;
assign micromatrizz[56][190] = 9'b111110111;
assign micromatrizz[56][191] = 9'b111111111;
assign micromatrizz[56][192] = 9'b111111111;
assign micromatrizz[56][193] = 9'b111111111;
assign micromatrizz[56][194] = 9'b111111111;
assign micromatrizz[56][195] = 9'b111110010;
assign micromatrizz[56][196] = 9'b111110011;
assign micromatrizz[56][197] = 9'b111110011;
assign micromatrizz[56][198] = 9'b111110011;
assign micromatrizz[56][199] = 9'b111110010;
assign micromatrizz[56][200] = 9'b111110010;
assign micromatrizz[56][201] = 9'b111110011;
assign micromatrizz[56][202] = 9'b111110111;
assign micromatrizz[56][203] = 9'b111111111;
assign micromatrizz[56][204] = 9'b111111111;
assign micromatrizz[56][205] = 9'b111111111;
assign micromatrizz[56][206] = 9'b111111111;
assign micromatrizz[56][207] = 9'b111110010;
assign micromatrizz[56][208] = 9'b111110011;
assign micromatrizz[56][209] = 9'b111110011;
assign micromatrizz[56][210] = 9'b111110011;
assign micromatrizz[56][211] = 9'b111110011;
assign micromatrizz[56][212] = 9'b111110011;
assign micromatrizz[56][213] = 9'b111110111;
assign micromatrizz[56][214] = 9'b111111111;
assign micromatrizz[56][215] = 9'b111111111;
assign micromatrizz[56][216] = 9'b111111111;
assign micromatrizz[56][217] = 9'b111111111;
assign micromatrizz[56][218] = 9'b111111111;
assign micromatrizz[56][219] = 9'b111111111;
assign micromatrizz[56][220] = 9'b111110010;
assign micromatrizz[56][221] = 9'b111111111;
assign micromatrizz[56][222] = 9'b111111111;
assign micromatrizz[56][223] = 9'b111111111;
assign micromatrizz[56][224] = 9'b111111111;
assign micromatrizz[56][225] = 9'b111110111;
assign micromatrizz[56][226] = 9'b111110010;
assign micromatrizz[56][227] = 9'b111110010;
assign micromatrizz[56][228] = 9'b111110010;
assign micromatrizz[56][229] = 9'b111110010;
assign micromatrizz[56][230] = 9'b111110011;
assign micromatrizz[56][231] = 9'b111110011;
assign micromatrizz[56][232] = 9'b111110011;
assign micromatrizz[56][233] = 9'b111111111;
assign micromatrizz[56][234] = 9'b111111111;
assign micromatrizz[56][235] = 9'b111111111;
assign micromatrizz[56][236] = 9'b111111111;
assign micromatrizz[56][237] = 9'b111111111;
assign micromatrizz[56][238] = 9'b111111111;
assign micromatrizz[56][239] = 9'b111111111;
assign micromatrizz[56][240] = 9'b111111111;
assign micromatrizz[56][241] = 9'b111111111;
assign micromatrizz[56][242] = 9'b111110010;
assign micromatrizz[56][243] = 9'b111110010;
assign micromatrizz[56][244] = 9'b111110011;
assign micromatrizz[56][245] = 9'b111110011;
assign micromatrizz[56][246] = 9'b111110011;
assign micromatrizz[56][247] = 9'b111110111;
assign micromatrizz[56][248] = 9'b111111111;
assign micromatrizz[56][249] = 9'b111111111;
assign micromatrizz[56][250] = 9'b111111111;
assign micromatrizz[56][251] = 9'b111110110;
assign micromatrizz[56][252] = 9'b111110010;
assign micromatrizz[56][253] = 9'b111110010;
assign micromatrizz[56][254] = 9'b111110011;
assign micromatrizz[56][255] = 9'b111110011;
assign micromatrizz[56][256] = 9'b111111111;
assign micromatrizz[56][257] = 9'b111111111;
assign micromatrizz[56][258] = 9'b111111111;
assign micromatrizz[56][259] = 9'b111110111;
assign micromatrizz[56][260] = 9'b111110010;
assign micromatrizz[56][261] = 9'b111110010;
assign micromatrizz[56][262] = 9'b111110010;
assign micromatrizz[56][263] = 9'b111110010;
assign micromatrizz[56][264] = 9'b111110010;
assign micromatrizz[56][265] = 9'b111110011;
assign micromatrizz[56][266] = 9'b111110111;
assign micromatrizz[56][267] = 9'b111111111;
assign micromatrizz[56][268] = 9'b111111111;
assign micromatrizz[56][269] = 9'b111111111;
assign micromatrizz[56][270] = 9'b111111111;
assign micromatrizz[56][271] = 9'b111111111;
assign micromatrizz[56][272] = 9'b111111111;
assign micromatrizz[56][273] = 9'b111111111;
assign micromatrizz[56][274] = 9'b111111111;
assign micromatrizz[56][275] = 9'b111111111;
assign micromatrizz[56][276] = 9'b111111111;
assign micromatrizz[56][277] = 9'b111111111;
assign micromatrizz[56][278] = 9'b111111111;
assign micromatrizz[56][279] = 9'b111111111;
assign micromatrizz[56][280] = 9'b111111111;
assign micromatrizz[56][281] = 9'b111111111;
assign micromatrizz[56][282] = 9'b111111111;
assign micromatrizz[56][283] = 9'b111111111;
assign micromatrizz[56][284] = 9'b111111111;
assign micromatrizz[56][285] = 9'b111111111;
assign micromatrizz[56][286] = 9'b111110010;
assign micromatrizz[56][287] = 9'b111110010;
assign micromatrizz[56][288] = 9'b111110010;
assign micromatrizz[56][289] = 9'b111110011;
assign micromatrizz[56][290] = 9'b111110011;
assign micromatrizz[56][291] = 9'b111110011;
assign micromatrizz[56][292] = 9'b111110010;
assign micromatrizz[56][293] = 9'b111111111;
assign micromatrizz[56][294] = 9'b111111111;
assign micromatrizz[56][295] = 9'b111111111;
assign micromatrizz[56][296] = 9'b111111111;
assign micromatrizz[56][297] = 9'b111110111;
assign micromatrizz[56][298] = 9'b111110010;
assign micromatrizz[56][299] = 9'b111110010;
assign micromatrizz[56][300] = 9'b111110011;
assign micromatrizz[56][301] = 9'b111110011;
assign micromatrizz[56][302] = 9'b111110011;
assign micromatrizz[56][303] = 9'b111110011;
assign micromatrizz[56][304] = 9'b111110011;
assign micromatrizz[56][305] = 9'b111110011;
assign micromatrizz[56][306] = 9'b111110111;
assign micromatrizz[56][307] = 9'b111111111;
assign micromatrizz[56][308] = 9'b111111111;
assign micromatrizz[56][309] = 9'b111111111;
assign micromatrizz[56][310] = 9'b111111111;
assign micromatrizz[56][311] = 9'b111110111;
assign micromatrizz[56][312] = 9'b111110010;
assign micromatrizz[56][313] = 9'b111111111;
assign micromatrizz[56][314] = 9'b111111111;
assign micromatrizz[56][315] = 9'b111111111;
assign micromatrizz[56][316] = 9'b111110111;
assign micromatrizz[56][317] = 9'b111110010;
assign micromatrizz[56][318] = 9'b111110010;
assign micromatrizz[56][319] = 9'b111110010;
assign micromatrizz[56][320] = 9'b111110010;
assign micromatrizz[56][321] = 9'b111110011;
assign micromatrizz[56][322] = 9'b111111111;
assign micromatrizz[56][323] = 9'b111111111;
assign micromatrizz[56][324] = 9'b111111111;
assign micromatrizz[56][325] = 9'b111111111;
assign micromatrizz[56][326] = 9'b111110010;
assign micromatrizz[56][327] = 9'b111110010;
assign micromatrizz[56][328] = 9'b111110010;
assign micromatrizz[56][329] = 9'b111110010;
assign micromatrizz[56][330] = 9'b111110111;
assign micromatrizz[56][331] = 9'b111111111;
assign micromatrizz[56][332] = 9'b111111111;
assign micromatrizz[56][333] = 9'b111111111;
assign micromatrizz[56][334] = 9'b111111111;
assign micromatrizz[56][335] = 9'b111110010;
assign micromatrizz[56][336] = 9'b111110010;
assign micromatrizz[56][337] = 9'b111110010;
assign micromatrizz[56][338] = 9'b111110011;
assign micromatrizz[56][339] = 9'b111110011;
assign micromatrizz[56][340] = 9'b111110011;
assign micromatrizz[56][341] = 9'b111110010;
assign micromatrizz[56][342] = 9'b111110111;
assign micromatrizz[56][343] = 9'b111111111;
assign micromatrizz[56][344] = 9'b111111111;
assign micromatrizz[56][345] = 9'b111111111;
assign micromatrizz[56][346] = 9'b111111111;
assign micromatrizz[56][347] = 9'b111110010;
assign micromatrizz[56][348] = 9'b111110010;
assign micromatrizz[56][349] = 9'b111110011;
assign micromatrizz[56][350] = 9'b111110011;
assign micromatrizz[56][351] = 9'b111110011;
assign micromatrizz[56][352] = 9'b111110011;
assign micromatrizz[56][353] = 9'b111110011;
assign micromatrizz[56][354] = 9'b111111111;
assign micromatrizz[56][355] = 9'b111111111;
assign micromatrizz[56][356] = 9'b111111111;
assign micromatrizz[56][357] = 9'b111111111;
assign micromatrizz[56][358] = 9'b111111111;
assign micromatrizz[56][359] = 9'b111110010;
assign micromatrizz[56][360] = 9'b111110011;
assign micromatrizz[56][361] = 9'b111110010;
assign micromatrizz[56][362] = 9'b111110010;
assign micromatrizz[56][363] = 9'b111110011;
assign micromatrizz[56][364] = 9'b111110011;
assign micromatrizz[56][365] = 9'b111110011;
assign micromatrizz[56][366] = 9'b111111111;
assign micromatrizz[56][367] = 9'b111111111;
assign micromatrizz[56][368] = 9'b111111111;
assign micromatrizz[56][369] = 9'b111111111;
assign micromatrizz[56][370] = 9'b111111111;
assign micromatrizz[56][371] = 9'b111111111;
assign micromatrizz[56][372] = 9'b111110010;
assign micromatrizz[56][373] = 9'b111110011;
assign micromatrizz[56][374] = 9'b111110011;
assign micromatrizz[56][375] = 9'b111110011;
assign micromatrizz[56][376] = 9'b111110011;
assign micromatrizz[56][377] = 9'b111110011;
assign micromatrizz[56][378] = 9'b111110011;
assign micromatrizz[56][379] = 9'b111111111;
assign micromatrizz[56][380] = 9'b111111111;
assign micromatrizz[56][381] = 9'b111111111;
assign micromatrizz[56][382] = 9'b111111111;
assign micromatrizz[56][383] = 9'b111110111;
assign micromatrizz[56][384] = 9'b111110010;
assign micromatrizz[56][385] = 9'b111110010;
assign micromatrizz[56][386] = 9'b111110011;
assign micromatrizz[56][387] = 9'b111110011;
assign micromatrizz[56][388] = 9'b111110011;
assign micromatrizz[56][389] = 9'b111110011;
assign micromatrizz[56][390] = 9'b111110011;
assign micromatrizz[56][391] = 9'b111111111;
assign micromatrizz[56][392] = 9'b111111111;
assign micromatrizz[56][393] = 9'b111111111;
assign micromatrizz[56][394] = 9'b111111111;
assign micromatrizz[56][395] = 9'b111110010;
assign micromatrizz[56][396] = 9'b111110010;
assign micromatrizz[56][397] = 9'b111110010;
assign micromatrizz[56][398] = 9'b111110010;
assign micromatrizz[56][399] = 9'b111110011;
assign micromatrizz[56][400] = 9'b111110011;
assign micromatrizz[56][401] = 9'b111110011;
assign micromatrizz[56][402] = 9'b111110011;
assign micromatrizz[56][403] = 9'b111111111;
assign micromatrizz[56][404] = 9'b111111111;
assign micromatrizz[56][405] = 9'b111111111;
assign micromatrizz[56][406] = 9'b111111111;
assign micromatrizz[56][407] = 9'b111111111;
assign micromatrizz[56][408] = 9'b111111111;
assign micromatrizz[56][409] = 9'b111111111;
assign micromatrizz[56][410] = 9'b111111111;
assign micromatrizz[56][411] = 9'b111111111;
assign micromatrizz[56][412] = 9'b111110110;
assign micromatrizz[56][413] = 9'b111110011;
assign micromatrizz[56][414] = 9'b111110010;
assign micromatrizz[56][415] = 9'b111110011;
assign micromatrizz[56][416] = 9'b111110010;
assign micromatrizz[56][417] = 9'b111110111;
assign micromatrizz[56][418] = 9'b111111111;
assign micromatrizz[56][419] = 9'b111111111;
assign micromatrizz[56][420] = 9'b111111111;
assign micromatrizz[56][421] = 9'b111110111;
assign micromatrizz[56][422] = 9'b111110010;
assign micromatrizz[56][423] = 9'b111110011;
assign micromatrizz[56][424] = 9'b111110011;
assign micromatrizz[56][425] = 9'b111110010;
assign micromatrizz[56][426] = 9'b111111111;
assign micromatrizz[56][427] = 9'b111111111;
assign micromatrizz[56][428] = 9'b111111111;
assign micromatrizz[56][429] = 9'b111111111;
assign micromatrizz[56][430] = 9'b111110111;
assign micromatrizz[56][431] = 9'b111110010;
assign micromatrizz[56][432] = 9'b111110010;
assign micromatrizz[56][433] = 9'b111110010;
assign micromatrizz[56][434] = 9'b111110011;
assign micromatrizz[56][435] = 9'b111110011;
assign micromatrizz[56][436] = 9'b111110011;
assign micromatrizz[56][437] = 9'b111110011;
assign micromatrizz[56][438] = 9'b111110111;
assign micromatrizz[56][439] = 9'b111111111;
assign micromatrizz[56][440] = 9'b111111111;
assign micromatrizz[56][441] = 9'b111111111;
assign micromatrizz[56][442] = 9'b111111111;
assign micromatrizz[56][443] = 9'b111111111;
assign micromatrizz[56][444] = 9'b111111111;
assign micromatrizz[56][445] = 9'b111111111;
assign micromatrizz[56][446] = 9'b111111111;
assign micromatrizz[56][447] = 9'b111110110;
assign micromatrizz[56][448] = 9'b111110010;
assign micromatrizz[56][449] = 9'b111110011;
assign micromatrizz[56][450] = 9'b111110010;
assign micromatrizz[56][451] = 9'b111110011;
assign micromatrizz[56][452] = 9'b111110011;
assign micromatrizz[56][453] = 9'b111110011;
assign micromatrizz[56][454] = 9'b111111111;
assign micromatrizz[56][455] = 9'b111111111;
assign micromatrizz[56][456] = 9'b111111111;
assign micromatrizz[56][457] = 9'b111111111;
assign micromatrizz[56][458] = 9'b111111111;
assign micromatrizz[56][459] = 9'b111111111;
assign micromatrizz[56][460] = 9'b111110111;
assign micromatrizz[56][461] = 9'b111110110;
assign micromatrizz[56][462] = 9'b111111111;
assign micromatrizz[56][463] = 9'b111111111;
assign micromatrizz[56][464] = 9'b111111111;
assign micromatrizz[56][465] = 9'b111110010;
assign micromatrizz[56][466] = 9'b111110010;
assign micromatrizz[56][467] = 9'b111110011;
assign micromatrizz[56][468] = 9'b111110010;
assign micromatrizz[56][469] = 9'b111110010;
assign micromatrizz[56][470] = 9'b111110011;
assign micromatrizz[56][471] = 9'b111110011;
assign micromatrizz[56][472] = 9'b111111111;
assign micromatrizz[56][473] = 9'b111111111;
assign micromatrizz[56][474] = 9'b111111111;
assign micromatrizz[56][475] = 9'b111111111;
assign micromatrizz[56][476] = 9'b111111111;
assign micromatrizz[56][477] = 9'b111111111;
assign micromatrizz[56][478] = 9'b111111111;
assign micromatrizz[56][479] = 9'b111111111;
assign micromatrizz[56][480] = 9'b111111111;
assign micromatrizz[56][481] = 9'b111110010;
assign micromatrizz[56][482] = 9'b111110010;
assign micromatrizz[56][483] = 9'b111110010;
assign micromatrizz[56][484] = 9'b111110010;
assign micromatrizz[56][485] = 9'b111110011;
assign micromatrizz[56][486] = 9'b111110011;
assign micromatrizz[56][487] = 9'b111110011;
assign micromatrizz[56][488] = 9'b111110011;
assign micromatrizz[56][489] = 9'b111111111;
assign micromatrizz[56][490] = 9'b111111111;
assign micromatrizz[56][491] = 9'b111111111;
assign micromatrizz[56][492] = 9'b111111111;
assign micromatrizz[56][493] = 9'b111111111;
assign micromatrizz[56][494] = 9'b111111111;
assign micromatrizz[56][495] = 9'b111111111;
assign micromatrizz[56][496] = 9'b111111111;
assign micromatrizz[56][497] = 9'b111111111;
assign micromatrizz[56][498] = 9'b111110010;
assign micromatrizz[56][499] = 9'b111110010;
assign micromatrizz[56][500] = 9'b111110010;
assign micromatrizz[56][501] = 9'b111110011;
assign micromatrizz[56][502] = 9'b111110010;
assign micromatrizz[56][503] = 9'b111110111;
assign micromatrizz[56][504] = 9'b111111111;
assign micromatrizz[56][505] = 9'b111111111;
assign micromatrizz[56][506] = 9'b111111111;
assign micromatrizz[56][507] = 9'b111110010;
assign micromatrizz[56][508] = 9'b111110010;
assign micromatrizz[56][509] = 9'b111110010;
assign micromatrizz[56][510] = 9'b111110011;
assign micromatrizz[56][511] = 9'b111110011;
assign micromatrizz[56][512] = 9'b111111111;
assign micromatrizz[56][513] = 9'b111111111;
assign micromatrizz[56][514] = 9'b111111111;
assign micromatrizz[56][515] = 9'b111111111;
assign micromatrizz[56][516] = 9'b111110111;
assign micromatrizz[56][517] = 9'b111110010;
assign micromatrizz[56][518] = 9'b111110011;
assign micromatrizz[56][519] = 9'b111110011;
assign micromatrizz[56][520] = 9'b111110010;
assign micromatrizz[56][521] = 9'b111110010;
assign micromatrizz[56][522] = 9'b111110011;
assign micromatrizz[56][523] = 9'b111110011;
assign micromatrizz[56][524] = 9'b111111111;
assign micromatrizz[56][525] = 9'b111111111;
assign micromatrizz[56][526] = 9'b111111111;
assign micromatrizz[56][527] = 9'b111111111;
assign micromatrizz[56][528] = 9'b111111111;
assign micromatrizz[56][529] = 9'b111110010;
assign micromatrizz[56][530] = 9'b111110011;
assign micromatrizz[56][531] = 9'b111110011;
assign micromatrizz[56][532] = 9'b111110011;
assign micromatrizz[56][533] = 9'b111110011;
assign micromatrizz[56][534] = 9'b111110011;
assign micromatrizz[56][535] = 9'b111110111;
assign micromatrizz[56][536] = 9'b111111111;
assign micromatrizz[56][537] = 9'b111111111;
assign micromatrizz[56][538] = 9'b111111111;
assign micromatrizz[56][539] = 9'b111110111;
assign micromatrizz[56][540] = 9'b111110010;
assign micromatrizz[56][541] = 9'b111110010;
assign micromatrizz[56][542] = 9'b111110011;
assign micromatrizz[56][543] = 9'b111110010;
assign micromatrizz[56][544] = 9'b111110010;
assign micromatrizz[56][545] = 9'b111111111;
assign micromatrizz[56][546] = 9'b111111111;
assign micromatrizz[56][547] = 9'b111111111;
assign micromatrizz[56][548] = 9'b111111111;
assign micromatrizz[56][549] = 9'b111110010;
assign micromatrizz[56][550] = 9'b111110011;
assign micromatrizz[56][551] = 9'b111110011;
assign micromatrizz[56][552] = 9'b111110011;
assign micromatrizz[56][553] = 9'b111110011;
assign micromatrizz[56][554] = 9'b111111111;
assign micromatrizz[56][555] = 9'b111111111;
assign micromatrizz[56][556] = 9'b111111111;
assign micromatrizz[56][557] = 9'b111111111;
assign micromatrizz[56][558] = 9'b111110010;
assign micromatrizz[56][559] = 9'b111110010;
assign micromatrizz[56][560] = 9'b111110010;
assign micromatrizz[56][561] = 9'b111110010;
assign micromatrizz[56][562] = 9'b111110011;
assign micromatrizz[56][563] = 9'b111110011;
assign micromatrizz[56][564] = 9'b111110010;
assign micromatrizz[56][565] = 9'b111111111;
assign micromatrizz[56][566] = 9'b111111111;
assign micromatrizz[56][567] = 9'b111111111;
assign micromatrizz[56][568] = 9'b111111111;
assign micromatrizz[56][569] = 9'b111110010;
assign micromatrizz[56][570] = 9'b111110010;
assign micromatrizz[56][571] = 9'b111110010;
assign micromatrizz[56][572] = 9'b111110010;
assign micromatrizz[56][573] = 9'b111110010;
assign micromatrizz[56][574] = 9'b111110011;
assign micromatrizz[56][575] = 9'b111110011;
assign micromatrizz[56][576] = 9'b111111111;
assign micromatrizz[56][577] = 9'b111111111;
assign micromatrizz[56][578] = 9'b111111111;
assign micromatrizz[56][579] = 9'b111111111;
assign micromatrizz[56][580] = 9'b111111111;
assign micromatrizz[56][581] = 9'b111110010;
assign micromatrizz[56][582] = 9'b111110011;
assign micromatrizz[56][583] = 9'b111110011;
assign micromatrizz[56][584] = 9'b111110010;
assign micromatrizz[56][585] = 9'b111110010;
assign micromatrizz[56][586] = 9'b111110011;
assign micromatrizz[56][587] = 9'b111110011;
assign micromatrizz[56][588] = 9'b111110111;
assign micromatrizz[56][589] = 9'b111111111;
assign micromatrizz[56][590] = 9'b111111111;
assign micromatrizz[56][591] = 9'b111111111;
assign micromatrizz[56][592] = 9'b111110111;
assign micromatrizz[56][593] = 9'b111110010;
assign micromatrizz[56][594] = 9'b111110011;
assign micromatrizz[56][595] = 9'b111110011;
assign micromatrizz[56][596] = 9'b111110011;
assign micromatrizz[56][597] = 9'b111110010;
assign micromatrizz[56][598] = 9'b111111111;
assign micromatrizz[56][599] = 9'b111111111;
assign micromatrizz[56][600] = 9'b111111111;
assign micromatrizz[56][601] = 9'b111111111;
assign micromatrizz[56][602] = 9'b111110010;
assign micromatrizz[56][603] = 9'b111110010;
assign micromatrizz[56][604] = 9'b111110011;
assign micromatrizz[56][605] = 9'b111110011;
assign micromatrizz[56][606] = 9'b111110011;
assign micromatrizz[56][607] = 9'b111111111;
assign micromatrizz[56][608] = 9'b111111111;
assign micromatrizz[56][609] = 9'b111111111;
assign micromatrizz[56][610] = 9'b111110010;
assign micromatrizz[56][611] = 9'b111110011;
assign micromatrizz[56][612] = 9'b111110010;
assign micromatrizz[56][613] = 9'b111110010;
assign micromatrizz[56][614] = 9'b111110011;
assign micromatrizz[56][615] = 9'b111110010;
assign micromatrizz[56][616] = 9'b111110011;
assign micromatrizz[56][617] = 9'b111110111;
assign micromatrizz[56][618] = 9'b111111111;
assign micromatrizz[56][619] = 9'b111111111;
assign micromatrizz[56][620] = 9'b111111111;
assign micromatrizz[56][621] = 9'b111111111;
assign micromatrizz[56][622] = 9'b111111111;
assign micromatrizz[56][623] = 9'b111111111;
assign micromatrizz[56][624] = 9'b111111111;
assign micromatrizz[56][625] = 9'b111111111;
assign micromatrizz[56][626] = 9'b111111111;
assign micromatrizz[56][627] = 9'b111111111;
assign micromatrizz[56][628] = 9'b111111111;
assign micromatrizz[56][629] = 9'b111111111;
assign micromatrizz[56][630] = 9'b111111111;
assign micromatrizz[56][631] = 9'b111111111;
assign micromatrizz[56][632] = 9'b111111111;
assign micromatrizz[56][633] = 9'b111111111;
assign micromatrizz[56][634] = 9'b111111111;
assign micromatrizz[56][635] = 9'b111111111;
assign micromatrizz[56][636] = 9'b111111111;
assign micromatrizz[56][637] = 9'b111111111;
assign micromatrizz[56][638] = 9'b111111111;
assign micromatrizz[56][639] = 9'b111111111;
assign micromatrizz[57][0] = 9'b111111111;
assign micromatrizz[57][1] = 9'b111111111;
assign micromatrizz[57][2] = 9'b111111111;
assign micromatrizz[57][3] = 9'b111111111;
assign micromatrizz[57][4] = 9'b111111111;
assign micromatrizz[57][5] = 9'b111111111;
assign micromatrizz[57][6] = 9'b111111111;
assign micromatrizz[57][7] = 9'b111110111;
assign micromatrizz[57][8] = 9'b111110010;
assign micromatrizz[57][9] = 9'b111110010;
assign micromatrizz[57][10] = 9'b111110010;
assign micromatrizz[57][11] = 9'b111110011;
assign micromatrizz[57][12] = 9'b111110011;
assign micromatrizz[57][13] = 9'b111110011;
assign micromatrizz[57][14] = 9'b111110011;
assign micromatrizz[57][15] = 9'b111110011;
assign micromatrizz[57][16] = 9'b111111111;
assign micromatrizz[57][17] = 9'b111111111;
assign micromatrizz[57][18] = 9'b111111111;
assign micromatrizz[57][19] = 9'b111111111;
assign micromatrizz[57][20] = 9'b111111111;
assign micromatrizz[57][21] = 9'b111111111;
assign micromatrizz[57][22] = 9'b111111111;
assign micromatrizz[57][23] = 9'b111111111;
assign micromatrizz[57][24] = 9'b111110010;
assign micromatrizz[57][25] = 9'b111110010;
assign micromatrizz[57][26] = 9'b111110010;
assign micromatrizz[57][27] = 9'b111110011;
assign micromatrizz[57][28] = 9'b111110011;
assign micromatrizz[57][29] = 9'b111110011;
assign micromatrizz[57][30] = 9'b111110011;
assign micromatrizz[57][31] = 9'b111111111;
assign micromatrizz[57][32] = 9'b111111111;
assign micromatrizz[57][33] = 9'b111111111;
assign micromatrizz[57][34] = 9'b111111111;
assign micromatrizz[57][35] = 9'b111110111;
assign micromatrizz[57][36] = 9'b111110010;
assign micromatrizz[57][37] = 9'b111110010;
assign micromatrizz[57][38] = 9'b111110011;
assign micromatrizz[57][39] = 9'b111110011;
assign micromatrizz[57][40] = 9'b111110011;
assign micromatrizz[57][41] = 9'b111110011;
assign micromatrizz[57][42] = 9'b111110011;
assign micromatrizz[57][43] = 9'b111111111;
assign micromatrizz[57][44] = 9'b111111111;
assign micromatrizz[57][45] = 9'b111111111;
assign micromatrizz[57][46] = 9'b111111111;
assign micromatrizz[57][47] = 9'b111110010;
assign micromatrizz[57][48] = 9'b111110010;
assign micromatrizz[57][49] = 9'b111110010;
assign micromatrizz[57][50] = 9'b111110011;
assign micromatrizz[57][51] = 9'b111110011;
assign micromatrizz[57][52] = 9'b111110011;
assign micromatrizz[57][53] = 9'b111110011;
assign micromatrizz[57][54] = 9'b111110111;
assign micromatrizz[57][55] = 9'b111111111;
assign micromatrizz[57][56] = 9'b111111111;
assign micromatrizz[57][57] = 9'b111111111;
assign micromatrizz[57][58] = 9'b111111111;
assign micromatrizz[57][59] = 9'b111110010;
assign micromatrizz[57][60] = 9'b111110011;
assign micromatrizz[57][61] = 9'b111110010;
assign micromatrizz[57][62] = 9'b111110010;
assign micromatrizz[57][63] = 9'b111110010;
assign micromatrizz[57][64] = 9'b111110011;
assign micromatrizz[57][65] = 9'b111110011;
assign micromatrizz[57][66] = 9'b111111111;
assign micromatrizz[57][67] = 9'b111111111;
assign micromatrizz[57][68] = 9'b111111111;
assign micromatrizz[57][69] = 9'b111110010;
assign micromatrizz[57][70] = 9'b111110010;
assign micromatrizz[57][71] = 9'b111110010;
assign micromatrizz[57][72] = 9'b111110010;
assign micromatrizz[57][73] = 9'b111110011;
assign micromatrizz[57][74] = 9'b111110011;
assign micromatrizz[57][75] = 9'b111111111;
assign micromatrizz[57][76] = 9'b111111111;
assign micromatrizz[57][77] = 9'b111111111;
assign micromatrizz[57][78] = 9'b111111111;
assign micromatrizz[57][79] = 9'b111110010;
assign micromatrizz[57][80] = 9'b111110011;
assign micromatrizz[57][81] = 9'b111110011;
assign micromatrizz[57][82] = 9'b111110011;
assign micromatrizz[57][83] = 9'b111110011;
assign micromatrizz[57][84] = 9'b111111111;
assign micromatrizz[57][85] = 9'b111111111;
assign micromatrizz[57][86] = 9'b111111111;
assign micromatrizz[57][87] = 9'b111111111;
assign micromatrizz[57][88] = 9'b111110010;
assign micromatrizz[57][89] = 9'b111110010;
assign micromatrizz[57][90] = 9'b111110010;
assign micromatrizz[57][91] = 9'b111110011;
assign micromatrizz[57][92] = 9'b111110011;
assign micromatrizz[57][93] = 9'b111110011;
assign micromatrizz[57][94] = 9'b111110011;
assign micromatrizz[57][95] = 9'b111110111;
assign micromatrizz[57][96] = 9'b111111111;
assign micromatrizz[57][97] = 9'b111111111;
assign micromatrizz[57][98] = 9'b111111111;
assign micromatrizz[57][99] = 9'b111111111;
assign micromatrizz[57][100] = 9'b111111111;
assign micromatrizz[57][101] = 9'b111111111;
assign micromatrizz[57][102] = 9'b111111111;
assign micromatrizz[57][103] = 9'b111111111;
assign micromatrizz[57][104] = 9'b111110010;
assign micromatrizz[57][105] = 9'b111110010;
assign micromatrizz[57][106] = 9'b111110010;
assign micromatrizz[57][107] = 9'b111110011;
assign micromatrizz[57][108] = 9'b111110011;
assign micromatrizz[57][109] = 9'b111110011;
assign micromatrizz[57][110] = 9'b111110011;
assign micromatrizz[57][111] = 9'b111110011;
assign micromatrizz[57][112] = 9'b111111111;
assign micromatrizz[57][113] = 9'b111111111;
assign micromatrizz[57][114] = 9'b111111111;
assign micromatrizz[57][115] = 9'b111111111;
assign micromatrizz[57][116] = 9'b111111111;
assign micromatrizz[57][117] = 9'b111111111;
assign micromatrizz[57][118] = 9'b111111111;
assign micromatrizz[57][119] = 9'b111111111;
assign micromatrizz[57][120] = 9'b111110010;
assign micromatrizz[57][121] = 9'b111110010;
assign micromatrizz[57][122] = 9'b111110010;
assign micromatrizz[57][123] = 9'b111110011;
assign micromatrizz[57][124] = 9'b111110011;
assign micromatrizz[57][125] = 9'b111110011;
assign micromatrizz[57][126] = 9'b111110111;
assign micromatrizz[57][127] = 9'b111111111;
assign micromatrizz[57][128] = 9'b111111111;
assign micromatrizz[57][129] = 9'b111111111;
assign micromatrizz[57][130] = 9'b111111111;
assign micromatrizz[57][131] = 9'b111111111;
assign micromatrizz[57][132] = 9'b111111111;
assign micromatrizz[57][133] = 9'b111111111;
assign micromatrizz[57][134] = 9'b111110111;
assign micromatrizz[57][135] = 9'b111111111;
assign micromatrizz[57][136] = 9'b111111111;
assign micromatrizz[57][137] = 9'b111111111;
assign micromatrizz[57][138] = 9'b111110111;
assign micromatrizz[57][139] = 9'b111110010;
assign micromatrizz[57][140] = 9'b111110010;
assign micromatrizz[57][141] = 9'b111110010;
assign micromatrizz[57][142] = 9'b111110010;
assign micromatrizz[57][143] = 9'b111110011;
assign micromatrizz[57][144] = 9'b111110011;
assign micromatrizz[57][145] = 9'b111110011;
assign micromatrizz[57][146] = 9'b111111111;
assign micromatrizz[57][147] = 9'b111111111;
assign micromatrizz[57][148] = 9'b111111111;
assign micromatrizz[57][149] = 9'b111111111;
assign micromatrizz[57][150] = 9'b111110111;
assign micromatrizz[57][151] = 9'b111110010;
assign micromatrizz[57][152] = 9'b111110011;
assign micromatrizz[57][153] = 9'b111110011;
assign micromatrizz[57][154] = 9'b111110011;
assign micromatrizz[57][155] = 9'b111110011;
assign micromatrizz[57][156] = 9'b111110011;
assign micromatrizz[57][157] = 9'b111110111;
assign micromatrizz[57][158] = 9'b111111111;
assign micromatrizz[57][159] = 9'b111111111;
assign micromatrizz[57][160] = 9'b111111111;
assign micromatrizz[57][161] = 9'b111111111;
assign micromatrizz[57][162] = 9'b111111111;
assign micromatrizz[57][163] = 9'b111111111;
assign micromatrizz[57][164] = 9'b111111111;
assign micromatrizz[57][165] = 9'b111111111;
assign micromatrizz[57][166] = 9'b111111111;
assign micromatrizz[57][167] = 9'b111111111;
assign micromatrizz[57][168] = 9'b111111111;
assign micromatrizz[57][169] = 9'b111111111;
assign micromatrizz[57][170] = 9'b111111111;
assign micromatrizz[57][171] = 9'b111111111;
assign micromatrizz[57][172] = 9'b111110010;
assign micromatrizz[57][173] = 9'b111110010;
assign micromatrizz[57][174] = 9'b111110010;
assign micromatrizz[57][175] = 9'b111110011;
assign micromatrizz[57][176] = 9'b111110011;
assign micromatrizz[57][177] = 9'b111110011;
assign micromatrizz[57][178] = 9'b111110011;
assign micromatrizz[57][179] = 9'b111110111;
assign micromatrizz[57][180] = 9'b111111111;
assign micromatrizz[57][181] = 9'b111111111;
assign micromatrizz[57][182] = 9'b111111111;
assign micromatrizz[57][183] = 9'b111110010;
assign micromatrizz[57][184] = 9'b111110010;
assign micromatrizz[57][185] = 9'b111110010;
assign micromatrizz[57][186] = 9'b111110010;
assign micromatrizz[57][187] = 9'b111110010;
assign micromatrizz[57][188] = 9'b111110010;
assign micromatrizz[57][189] = 9'b111110011;
assign micromatrizz[57][190] = 9'b111110111;
assign micromatrizz[57][191] = 9'b111111111;
assign micromatrizz[57][192] = 9'b111111111;
assign micromatrizz[57][193] = 9'b111111111;
assign micromatrizz[57][194] = 9'b111111111;
assign micromatrizz[57][195] = 9'b111110010;
assign micromatrizz[57][196] = 9'b111110010;
assign micromatrizz[57][197] = 9'b111110011;
assign micromatrizz[57][198] = 9'b111110011;
assign micromatrizz[57][199] = 9'b111110010;
assign micromatrizz[57][200] = 9'b111110010;
assign micromatrizz[57][201] = 9'b111110011;
assign micromatrizz[57][202] = 9'b111110111;
assign micromatrizz[57][203] = 9'b111111111;
assign micromatrizz[57][204] = 9'b111111111;
assign micromatrizz[57][205] = 9'b111111111;
assign micromatrizz[57][206] = 9'b111110110;
assign micromatrizz[57][207] = 9'b111110010;
assign micromatrizz[57][208] = 9'b111110010;
assign micromatrizz[57][209] = 9'b111110010;
assign micromatrizz[57][210] = 9'b111110011;
assign micromatrizz[57][211] = 9'b111110011;
assign micromatrizz[57][212] = 9'b111110011;
assign micromatrizz[57][213] = 9'b111110111;
assign micromatrizz[57][214] = 9'b111111111;
assign micromatrizz[57][215] = 9'b111111111;
assign micromatrizz[57][216] = 9'b111111111;
assign micromatrizz[57][217] = 9'b111111111;
assign micromatrizz[57][218] = 9'b111111111;
assign micromatrizz[57][219] = 9'b111111111;
assign micromatrizz[57][220] = 9'b111110111;
assign micromatrizz[57][221] = 9'b111110111;
assign micromatrizz[57][222] = 9'b111111111;
assign micromatrizz[57][223] = 9'b111111111;
assign micromatrizz[57][224] = 9'b111111111;
assign micromatrizz[57][225] = 9'b111110111;
assign micromatrizz[57][226] = 9'b111110010;
assign micromatrizz[57][227] = 9'b111110010;
assign micromatrizz[57][228] = 9'b111110010;
assign micromatrizz[57][229] = 9'b111110010;
assign micromatrizz[57][230] = 9'b111110011;
assign micromatrizz[57][231] = 9'b111110011;
assign micromatrizz[57][232] = 9'b111110111;
assign micromatrizz[57][233] = 9'b111111111;
assign micromatrizz[57][234] = 9'b111111111;
assign micromatrizz[57][235] = 9'b111111111;
assign micromatrizz[57][236] = 9'b111111111;
assign micromatrizz[57][237] = 9'b111111111;
assign micromatrizz[57][238] = 9'b111111111;
assign micromatrizz[57][239] = 9'b111111111;
assign micromatrizz[57][240] = 9'b111111111;
assign micromatrizz[57][241] = 9'b111111111;
assign micromatrizz[57][242] = 9'b111110010;
assign micromatrizz[57][243] = 9'b111110010;
assign micromatrizz[57][244] = 9'b111110010;
assign micromatrizz[57][245] = 9'b111110011;
assign micromatrizz[57][246] = 9'b111110011;
assign micromatrizz[57][247] = 9'b111110111;
assign micromatrizz[57][248] = 9'b111111111;
assign micromatrizz[57][249] = 9'b111111111;
assign micromatrizz[57][250] = 9'b111111111;
assign micromatrizz[57][251] = 9'b111110110;
assign micromatrizz[57][252] = 9'b111110010;
assign micromatrizz[57][253] = 9'b111110010;
assign micromatrizz[57][254] = 9'b111110011;
assign micromatrizz[57][255] = 9'b111110011;
assign micromatrizz[57][256] = 9'b111110111;
assign micromatrizz[57][257] = 9'b111111111;
assign micromatrizz[57][258] = 9'b111111111;
assign micromatrizz[57][259] = 9'b111110111;
assign micromatrizz[57][260] = 9'b111110010;
assign micromatrizz[57][261] = 9'b111110010;
assign micromatrizz[57][262] = 9'b111110011;
assign micromatrizz[57][263] = 9'b111110011;
assign micromatrizz[57][264] = 9'b111110011;
assign micromatrizz[57][265] = 9'b111110011;
assign micromatrizz[57][266] = 9'b111110010;
assign micromatrizz[57][267] = 9'b111110111;
assign micromatrizz[57][268] = 9'b111111111;
assign micromatrizz[57][269] = 9'b111111111;
assign micromatrizz[57][270] = 9'b111111111;
assign micromatrizz[57][271] = 9'b111111111;
assign micromatrizz[57][272] = 9'b111111111;
assign micromatrizz[57][273] = 9'b111111111;
assign micromatrizz[57][274] = 9'b111111111;
assign micromatrizz[57][275] = 9'b111111111;
assign micromatrizz[57][276] = 9'b111111111;
assign micromatrizz[57][277] = 9'b111111111;
assign micromatrizz[57][278] = 9'b111111111;
assign micromatrizz[57][279] = 9'b111111111;
assign micromatrizz[57][280] = 9'b111111111;
assign micromatrizz[57][281] = 9'b111111111;
assign micromatrizz[57][282] = 9'b111111111;
assign micromatrizz[57][283] = 9'b111111111;
assign micromatrizz[57][284] = 9'b111111111;
assign micromatrizz[57][285] = 9'b111111111;
assign micromatrizz[57][286] = 9'b111110010;
assign micromatrizz[57][287] = 9'b111110011;
assign micromatrizz[57][288] = 9'b111110010;
assign micromatrizz[57][289] = 9'b111110010;
assign micromatrizz[57][290] = 9'b111110011;
assign micromatrizz[57][291] = 9'b111110011;
assign micromatrizz[57][292] = 9'b111110011;
assign micromatrizz[57][293] = 9'b111110111;
assign micromatrizz[57][294] = 9'b111111111;
assign micromatrizz[57][295] = 9'b111111111;
assign micromatrizz[57][296] = 9'b111111111;
assign micromatrizz[57][297] = 9'b111111111;
assign micromatrizz[57][298] = 9'b111110111;
assign micromatrizz[57][299] = 9'b111110010;
assign micromatrizz[57][300] = 9'b111110011;
assign micromatrizz[57][301] = 9'b111110010;
assign micromatrizz[57][302] = 9'b111110011;
assign micromatrizz[57][303] = 9'b111110011;
assign micromatrizz[57][304] = 9'b111110011;
assign micromatrizz[57][305] = 9'b111110011;
assign micromatrizz[57][306] = 9'b111110011;
assign micromatrizz[57][307] = 9'b111111111;
assign micromatrizz[57][308] = 9'b111111111;
assign micromatrizz[57][309] = 9'b111111111;
assign micromatrizz[57][310] = 9'b111111111;
assign micromatrizz[57][311] = 9'b111110010;
assign micromatrizz[57][312] = 9'b111111111;
assign micromatrizz[57][313] = 9'b111111111;
assign micromatrizz[57][314] = 9'b111111111;
assign micromatrizz[57][315] = 9'b111111111;
assign micromatrizz[57][316] = 9'b111110010;
assign micromatrizz[57][317] = 9'b111110010;
assign micromatrizz[57][318] = 9'b111110010;
assign micromatrizz[57][319] = 9'b111110011;
assign micromatrizz[57][320] = 9'b111110011;
assign micromatrizz[57][321] = 9'b111110011;
assign micromatrizz[57][322] = 9'b111111111;
assign micromatrizz[57][323] = 9'b111111111;
assign micromatrizz[57][324] = 9'b111111111;
assign micromatrizz[57][325] = 9'b111111111;
assign micromatrizz[57][326] = 9'b111110010;
assign micromatrizz[57][327] = 9'b111110010;
assign micromatrizz[57][328] = 9'b111110010;
assign micromatrizz[57][329] = 9'b111110011;
assign micromatrizz[57][330] = 9'b111110010;
assign micromatrizz[57][331] = 9'b111111111;
assign micromatrizz[57][332] = 9'b111111111;
assign micromatrizz[57][333] = 9'b111111111;
assign micromatrizz[57][334] = 9'b111111111;
assign micromatrizz[57][335] = 9'b111110010;
assign micromatrizz[57][336] = 9'b111110010;
assign micromatrizz[57][337] = 9'b111110010;
assign micromatrizz[57][338] = 9'b111110011;
assign micromatrizz[57][339] = 9'b111110011;
assign micromatrizz[57][340] = 9'b111110011;
assign micromatrizz[57][341] = 9'b111110010;
assign micromatrizz[57][342] = 9'b111111111;
assign micromatrizz[57][343] = 9'b111111111;
assign micromatrizz[57][344] = 9'b111111111;
assign micromatrizz[57][345] = 9'b111111111;
assign micromatrizz[57][346] = 9'b111111111;
assign micromatrizz[57][347] = 9'b111110010;
assign micromatrizz[57][348] = 9'b111110010;
assign micromatrizz[57][349] = 9'b111110010;
assign micromatrizz[57][350] = 9'b111110011;
assign micromatrizz[57][351] = 9'b111110011;
assign micromatrizz[57][352] = 9'b111110011;
assign micromatrizz[57][353] = 9'b111110011;
assign micromatrizz[57][354] = 9'b111111111;
assign micromatrizz[57][355] = 9'b111111111;
assign micromatrizz[57][356] = 9'b111111111;
assign micromatrizz[57][357] = 9'b111111111;
assign micromatrizz[57][358] = 9'b111111111;
assign micromatrizz[57][359] = 9'b111110010;
assign micromatrizz[57][360] = 9'b111110011;
assign micromatrizz[57][361] = 9'b111110010;
assign micromatrizz[57][362] = 9'b111110010;
assign micromatrizz[57][363] = 9'b111110011;
assign micromatrizz[57][364] = 9'b111110011;
assign micromatrizz[57][365] = 9'b111110011;
assign micromatrizz[57][366] = 9'b111111111;
assign micromatrizz[57][367] = 9'b111111111;
assign micromatrizz[57][368] = 9'b111111111;
assign micromatrizz[57][369] = 9'b111111111;
assign micromatrizz[57][370] = 9'b111111111;
assign micromatrizz[57][371] = 9'b111111111;
assign micromatrizz[57][372] = 9'b111110010;
assign micromatrizz[57][373] = 9'b111110011;
assign micromatrizz[57][374] = 9'b111110011;
assign micromatrizz[57][375] = 9'b111110011;
assign micromatrizz[57][376] = 9'b111110011;
assign micromatrizz[57][377] = 9'b111110011;
assign micromatrizz[57][378] = 9'b111110011;
assign micromatrizz[57][379] = 9'b111111111;
assign micromatrizz[57][380] = 9'b111111111;
assign micromatrizz[57][381] = 9'b111111111;
assign micromatrizz[57][382] = 9'b111111111;
assign micromatrizz[57][383] = 9'b111110111;
assign micromatrizz[57][384] = 9'b111110010;
assign micromatrizz[57][385] = 9'b111110010;
assign micromatrizz[57][386] = 9'b111110011;
assign micromatrizz[57][387] = 9'b111110011;
assign micromatrizz[57][388] = 9'b111110011;
assign micromatrizz[57][389] = 9'b111110011;
assign micromatrizz[57][390] = 9'b111110011;
assign micromatrizz[57][391] = 9'b111111111;
assign micromatrizz[57][392] = 9'b111111111;
assign micromatrizz[57][393] = 9'b111111111;
assign micromatrizz[57][394] = 9'b111111111;
assign micromatrizz[57][395] = 9'b111110010;
assign micromatrizz[57][396] = 9'b111110010;
assign micromatrizz[57][397] = 9'b111110010;
assign micromatrizz[57][398] = 9'b111110010;
assign micromatrizz[57][399] = 9'b111110011;
assign micromatrizz[57][400] = 9'b111110011;
assign micromatrizz[57][401] = 9'b111110011;
assign micromatrizz[57][402] = 9'b111110111;
assign micromatrizz[57][403] = 9'b111111111;
assign micromatrizz[57][404] = 9'b111111111;
assign micromatrizz[57][405] = 9'b111111111;
assign micromatrizz[57][406] = 9'b111111111;
assign micromatrizz[57][407] = 9'b111111111;
assign micromatrizz[57][408] = 9'b111111111;
assign micromatrizz[57][409] = 9'b111111111;
assign micromatrizz[57][410] = 9'b111111111;
assign micromatrizz[57][411] = 9'b111110111;
assign micromatrizz[57][412] = 9'b111110010;
assign micromatrizz[57][413] = 9'b111110011;
assign micromatrizz[57][414] = 9'b111110010;
assign micromatrizz[57][415] = 9'b111110011;
assign micromatrizz[57][416] = 9'b111110011;
assign micromatrizz[57][417] = 9'b111110111;
assign micromatrizz[57][418] = 9'b111111111;
assign micromatrizz[57][419] = 9'b111111111;
assign micromatrizz[57][420] = 9'b111111111;
assign micromatrizz[57][421] = 9'b111110111;
assign micromatrizz[57][422] = 9'b111110010;
assign micromatrizz[57][423] = 9'b111110011;
assign micromatrizz[57][424] = 9'b111110011;
assign micromatrizz[57][425] = 9'b111110011;
assign micromatrizz[57][426] = 9'b111110111;
assign micromatrizz[57][427] = 9'b111111111;
assign micromatrizz[57][428] = 9'b111111111;
assign micromatrizz[57][429] = 9'b111111111;
assign micromatrizz[57][430] = 9'b111110111;
assign micromatrizz[57][431] = 9'b111110010;
assign micromatrizz[57][432] = 9'b111110010;
assign micromatrizz[57][433] = 9'b111110010;
assign micromatrizz[57][434] = 9'b111110011;
assign micromatrizz[57][435] = 9'b111110011;
assign micromatrizz[57][436] = 9'b111110011;
assign micromatrizz[57][437] = 9'b111110011;
assign micromatrizz[57][438] = 9'b111111111;
assign micromatrizz[57][439] = 9'b111111111;
assign micromatrizz[57][440] = 9'b111111111;
assign micromatrizz[57][441] = 9'b111111111;
assign micromatrizz[57][442] = 9'b111111111;
assign micromatrizz[57][443] = 9'b111111111;
assign micromatrizz[57][444] = 9'b111111111;
assign micromatrizz[57][445] = 9'b111111111;
assign micromatrizz[57][446] = 9'b111111111;
assign micromatrizz[57][447] = 9'b111110010;
assign micromatrizz[57][448] = 9'b111110010;
assign micromatrizz[57][449] = 9'b111110011;
assign micromatrizz[57][450] = 9'b111110011;
assign micromatrizz[57][451] = 9'b111110011;
assign micromatrizz[57][452] = 9'b111110011;
assign micromatrizz[57][453] = 9'b111110011;
assign micromatrizz[57][454] = 9'b111111111;
assign micromatrizz[57][455] = 9'b111111111;
assign micromatrizz[57][456] = 9'b111111111;
assign micromatrizz[57][457] = 9'b111111111;
assign micromatrizz[57][458] = 9'b111111111;
assign micromatrizz[57][459] = 9'b111111111;
assign micromatrizz[57][460] = 9'b111111111;
assign micromatrizz[57][461] = 9'b111110110;
assign micromatrizz[57][462] = 9'b111111111;
assign micromatrizz[57][463] = 9'b111111111;
assign micromatrizz[57][464] = 9'b111110111;
assign micromatrizz[57][465] = 9'b111110010;
assign micromatrizz[57][466] = 9'b111110010;
assign micromatrizz[57][467] = 9'b111110011;
assign micromatrizz[57][468] = 9'b111110011;
assign micromatrizz[57][469] = 9'b111110011;
assign micromatrizz[57][470] = 9'b111110011;
assign micromatrizz[57][471] = 9'b111110011;
assign micromatrizz[57][472] = 9'b111110011;
assign micromatrizz[57][473] = 9'b111111111;
assign micromatrizz[57][474] = 9'b111111111;
assign micromatrizz[57][475] = 9'b111111111;
assign micromatrizz[57][476] = 9'b111111111;
assign micromatrizz[57][477] = 9'b111111111;
assign micromatrizz[57][478] = 9'b111111111;
assign micromatrizz[57][479] = 9'b111111111;
assign micromatrizz[57][480] = 9'b111111111;
assign micromatrizz[57][481] = 9'b111110010;
assign micromatrizz[57][482] = 9'b111110010;
assign micromatrizz[57][483] = 9'b111110010;
assign micromatrizz[57][484] = 9'b111110010;
assign micromatrizz[57][485] = 9'b111110011;
assign micromatrizz[57][486] = 9'b111110011;
assign micromatrizz[57][487] = 9'b111110011;
assign micromatrizz[57][488] = 9'b111110111;
assign micromatrizz[57][489] = 9'b111111111;
assign micromatrizz[57][490] = 9'b111111111;
assign micromatrizz[57][491] = 9'b111111111;
assign micromatrizz[57][492] = 9'b111111111;
assign micromatrizz[57][493] = 9'b111111111;
assign micromatrizz[57][494] = 9'b111111111;
assign micromatrizz[57][495] = 9'b111111111;
assign micromatrizz[57][496] = 9'b111111111;
assign micromatrizz[57][497] = 9'b111110111;
assign micromatrizz[57][498] = 9'b111110010;
assign micromatrizz[57][499] = 9'b111110010;
assign micromatrizz[57][500] = 9'b111110011;
assign micromatrizz[57][501] = 9'b111110011;
assign micromatrizz[57][502] = 9'b111110010;
assign micromatrizz[57][503] = 9'b111110111;
assign micromatrizz[57][504] = 9'b111111111;
assign micromatrizz[57][505] = 9'b111111111;
assign micromatrizz[57][506] = 9'b111111111;
assign micromatrizz[57][507] = 9'b111110010;
assign micromatrizz[57][508] = 9'b111110010;
assign micromatrizz[57][509] = 9'b111110011;
assign micromatrizz[57][510] = 9'b111110011;
assign micromatrizz[57][511] = 9'b111110011;
assign micromatrizz[57][512] = 9'b111110111;
assign micromatrizz[57][513] = 9'b111111111;
assign micromatrizz[57][514] = 9'b111111111;
assign micromatrizz[57][515] = 9'b111111111;
assign micromatrizz[57][516] = 9'b111110111;
assign micromatrizz[57][517] = 9'b111110010;
assign micromatrizz[57][518] = 9'b111110011;
assign micromatrizz[57][519] = 9'b111110011;
assign micromatrizz[57][520] = 9'b111110010;
assign micromatrizz[57][521] = 9'b111110010;
assign micromatrizz[57][522] = 9'b111110010;
assign micromatrizz[57][523] = 9'b111110111;
assign micromatrizz[57][524] = 9'b111111111;
assign micromatrizz[57][525] = 9'b111111111;
assign micromatrizz[57][526] = 9'b111111111;
assign micromatrizz[57][527] = 9'b111111111;
assign micromatrizz[57][528] = 9'b111110111;
assign micromatrizz[57][529] = 9'b111110010;
assign micromatrizz[57][530] = 9'b111110011;
assign micromatrizz[57][531] = 9'b111110011;
assign micromatrizz[57][532] = 9'b111110011;
assign micromatrizz[57][533] = 9'b111110011;
assign micromatrizz[57][534] = 9'b111110011;
assign micromatrizz[57][535] = 9'b111110111;
assign micromatrizz[57][536] = 9'b111111111;
assign micromatrizz[57][537] = 9'b111111111;
assign micromatrizz[57][538] = 9'b111111111;
assign micromatrizz[57][539] = 9'b111110010;
assign micromatrizz[57][540] = 9'b111110010;
assign micromatrizz[57][541] = 9'b111110011;
assign micromatrizz[57][542] = 9'b111110010;
assign micromatrizz[57][543] = 9'b111110011;
assign micromatrizz[57][544] = 9'b111110010;
assign micromatrizz[57][545] = 9'b111111111;
assign micromatrizz[57][546] = 9'b111111111;
assign micromatrizz[57][547] = 9'b111111111;
assign micromatrizz[57][548] = 9'b111111111;
assign micromatrizz[57][549] = 9'b111110010;
assign micromatrizz[57][550] = 9'b111110011;
assign micromatrizz[57][551] = 9'b111110011;
assign micromatrizz[57][552] = 9'b111110011;
assign micromatrizz[57][553] = 9'b111110011;
assign micromatrizz[57][554] = 9'b111111111;
assign micromatrizz[57][555] = 9'b111111111;
assign micromatrizz[57][556] = 9'b111111111;
assign micromatrizz[57][557] = 9'b111111111;
assign micromatrizz[57][558] = 9'b111110010;
assign micromatrizz[57][559] = 9'b111110010;
assign micromatrizz[57][560] = 9'b111110010;
assign micromatrizz[57][561] = 9'b111110010;
assign micromatrizz[57][562] = 9'b111110011;
assign micromatrizz[57][563] = 9'b111110011;
assign micromatrizz[57][564] = 9'b111110010;
assign micromatrizz[57][565] = 9'b111111111;
assign micromatrizz[57][566] = 9'b111111111;
assign micromatrizz[57][567] = 9'b111111111;
assign micromatrizz[57][568] = 9'b111111111;
assign micromatrizz[57][569] = 9'b111110010;
assign micromatrizz[57][570] = 9'b111110010;
assign micromatrizz[57][571] = 9'b111110010;
assign micromatrizz[57][572] = 9'b111110010;
assign micromatrizz[57][573] = 9'b111110011;
assign micromatrizz[57][574] = 9'b111110011;
assign micromatrizz[57][575] = 9'b111110011;
assign micromatrizz[57][576] = 9'b111111111;
assign micromatrizz[57][577] = 9'b111111111;
assign micromatrizz[57][578] = 9'b111111111;
assign micromatrizz[57][579] = 9'b111111111;
assign micromatrizz[57][580] = 9'b111111111;
assign micromatrizz[57][581] = 9'b111110010;
assign micromatrizz[57][582] = 9'b111110011;
assign micromatrizz[57][583] = 9'b111110011;
assign micromatrizz[57][584] = 9'b111110010;
assign micromatrizz[57][585] = 9'b111110010;
assign micromatrizz[57][586] = 9'b111110011;
assign micromatrizz[57][587] = 9'b111110011;
assign micromatrizz[57][588] = 9'b111111111;
assign micromatrizz[57][589] = 9'b111111111;
assign micromatrizz[57][590] = 9'b111111111;
assign micromatrizz[57][591] = 9'b111111111;
assign micromatrizz[57][592] = 9'b111110010;
assign micromatrizz[57][593] = 9'b111110011;
assign micromatrizz[57][594] = 9'b111110010;
assign micromatrizz[57][595] = 9'b111110011;
assign micromatrizz[57][596] = 9'b111110011;
assign micromatrizz[57][597] = 9'b111110011;
assign micromatrizz[57][598] = 9'b111111111;
assign micromatrizz[57][599] = 9'b111111111;
assign micromatrizz[57][600] = 9'b111111111;
assign micromatrizz[57][601] = 9'b111111111;
assign micromatrizz[57][602] = 9'b111110010;
assign micromatrizz[57][603] = 9'b111110011;
assign micromatrizz[57][604] = 9'b111110011;
assign micromatrizz[57][605] = 9'b111110011;
assign micromatrizz[57][606] = 9'b111110010;
assign micromatrizz[57][607] = 9'b111111111;
assign micromatrizz[57][608] = 9'b111111111;
assign micromatrizz[57][609] = 9'b111111111;
assign micromatrizz[57][610] = 9'b111110010;
assign micromatrizz[57][611] = 9'b111110010;
assign micromatrizz[57][612] = 9'b111110010;
assign micromatrizz[57][613] = 9'b111110010;
assign micromatrizz[57][614] = 9'b111110010;
assign micromatrizz[57][615] = 9'b111110011;
assign micromatrizz[57][616] = 9'b111110011;
assign micromatrizz[57][617] = 9'b111110011;
assign micromatrizz[57][618] = 9'b111111111;
assign micromatrizz[57][619] = 9'b111111111;
assign micromatrizz[57][620] = 9'b111111111;
assign micromatrizz[57][621] = 9'b111111111;
assign micromatrizz[57][622] = 9'b111111111;
assign micromatrizz[57][623] = 9'b111111111;
assign micromatrizz[57][624] = 9'b111111111;
assign micromatrizz[57][625] = 9'b111111111;
assign micromatrizz[57][626] = 9'b111111111;
assign micromatrizz[57][627] = 9'b111111111;
assign micromatrizz[57][628] = 9'b111111111;
assign micromatrizz[57][629] = 9'b111111111;
assign micromatrizz[57][630] = 9'b111111111;
assign micromatrizz[57][631] = 9'b111111111;
assign micromatrizz[57][632] = 9'b111111111;
assign micromatrizz[57][633] = 9'b111111111;
assign micromatrizz[57][634] = 9'b111111111;
assign micromatrizz[57][635] = 9'b111111111;
assign micromatrizz[57][636] = 9'b111111111;
assign micromatrizz[57][637] = 9'b111111111;
assign micromatrizz[57][638] = 9'b111111111;
assign micromatrizz[57][639] = 9'b111111111;
assign micromatrizz[58][0] = 9'b111111111;
assign micromatrizz[58][1] = 9'b111111111;
assign micromatrizz[58][2] = 9'b111111111;
assign micromatrizz[58][3] = 9'b111111111;
assign micromatrizz[58][4] = 9'b111111111;
assign micromatrizz[58][5] = 9'b111111111;
assign micromatrizz[58][6] = 9'b111111111;
assign micromatrizz[58][7] = 9'b111111111;
assign micromatrizz[58][8] = 9'b111110010;
assign micromatrizz[58][9] = 9'b111110010;
assign micromatrizz[58][10] = 9'b111110011;
assign micromatrizz[58][11] = 9'b111110010;
assign micromatrizz[58][12] = 9'b111110011;
assign micromatrizz[58][13] = 9'b111110011;
assign micromatrizz[58][14] = 9'b111110011;
assign micromatrizz[58][15] = 9'b111110011;
assign micromatrizz[58][16] = 9'b111110011;
assign micromatrizz[58][17] = 9'b111111111;
assign micromatrizz[58][18] = 9'b111111111;
assign micromatrizz[58][19] = 9'b111111111;
assign micromatrizz[58][20] = 9'b111111111;
assign micromatrizz[58][21] = 9'b111111111;
assign micromatrizz[58][22] = 9'b111111111;
assign micromatrizz[58][23] = 9'b111110111;
assign micromatrizz[58][24] = 9'b111110010;
assign micromatrizz[58][25] = 9'b111110010;
assign micromatrizz[58][26] = 9'b111110010;
assign micromatrizz[58][27] = 9'b111110011;
assign micromatrizz[58][28] = 9'b111110011;
assign micromatrizz[58][29] = 9'b111110011;
assign micromatrizz[58][30] = 9'b111110011;
assign micromatrizz[58][31] = 9'b111111111;
assign micromatrizz[58][32] = 9'b111111111;
assign micromatrizz[58][33] = 9'b111111111;
assign micromatrizz[58][34] = 9'b111111111;
assign micromatrizz[58][35] = 9'b111110111;
assign micromatrizz[58][36] = 9'b111110010;
assign micromatrizz[58][37] = 9'b111110010;
assign micromatrizz[58][38] = 9'b111110011;
assign micromatrizz[58][39] = 9'b111110011;
assign micromatrizz[58][40] = 9'b111110011;
assign micromatrizz[58][41] = 9'b111110011;
assign micromatrizz[58][42] = 9'b111110011;
assign micromatrizz[58][43] = 9'b111111111;
assign micromatrizz[58][44] = 9'b111111111;
assign micromatrizz[58][45] = 9'b111111111;
assign micromatrizz[58][46] = 9'b111111111;
assign micromatrizz[58][47] = 9'b111110010;
assign micromatrizz[58][48] = 9'b111110010;
assign micromatrizz[58][49] = 9'b111110010;
assign micromatrizz[58][50] = 9'b111110011;
assign micromatrizz[58][51] = 9'b111110011;
assign micromatrizz[58][52] = 9'b111110011;
assign micromatrizz[58][53] = 9'b111110010;
assign micromatrizz[58][54] = 9'b111110111;
assign micromatrizz[58][55] = 9'b111111111;
assign micromatrizz[58][56] = 9'b111111111;
assign micromatrizz[58][57] = 9'b111111111;
assign micromatrizz[58][58] = 9'b111111111;
assign micromatrizz[58][59] = 9'b111110010;
assign micromatrizz[58][60] = 9'b111110010;
assign micromatrizz[58][61] = 9'b111110010;
assign micromatrizz[58][62] = 9'b111110010;
assign micromatrizz[58][63] = 9'b111110010;
assign micromatrizz[58][64] = 9'b111110011;
assign micromatrizz[58][65] = 9'b111110010;
assign micromatrizz[58][66] = 9'b111110111;
assign micromatrizz[58][67] = 9'b111111111;
assign micromatrizz[58][68] = 9'b111111111;
assign micromatrizz[58][69] = 9'b111110010;
assign micromatrizz[58][70] = 9'b111110010;
assign micromatrizz[58][71] = 9'b111110010;
assign micromatrizz[58][72] = 9'b111110010;
assign micromatrizz[58][73] = 9'b111110011;
assign micromatrizz[58][74] = 9'b111110010;
assign micromatrizz[58][75] = 9'b111111111;
assign micromatrizz[58][76] = 9'b111111111;
assign micromatrizz[58][77] = 9'b111111111;
assign micromatrizz[58][78] = 9'b111111111;
assign micromatrizz[58][79] = 9'b111110010;
assign micromatrizz[58][80] = 9'b111110010;
assign micromatrizz[58][81] = 9'b111110011;
assign micromatrizz[58][82] = 9'b111110011;
assign micromatrizz[58][83] = 9'b111110011;
assign micromatrizz[58][84] = 9'b111110111;
assign micromatrizz[58][85] = 9'b111111111;
assign micromatrizz[58][86] = 9'b111111111;
assign micromatrizz[58][87] = 9'b111111111;
assign micromatrizz[58][88] = 9'b111110010;
assign micromatrizz[58][89] = 9'b111110010;
assign micromatrizz[58][90] = 9'b111110010;
assign micromatrizz[58][91] = 9'b111110010;
assign micromatrizz[58][92] = 9'b111110011;
assign micromatrizz[58][93] = 9'b111110011;
assign micromatrizz[58][94] = 9'b111110011;
assign micromatrizz[58][95] = 9'b111111111;
assign micromatrizz[58][96] = 9'b111111111;
assign micromatrizz[58][97] = 9'b111111111;
assign micromatrizz[58][98] = 9'b111111111;
assign micromatrizz[58][99] = 9'b111111111;
assign micromatrizz[58][100] = 9'b111111111;
assign micromatrizz[58][101] = 9'b111111111;
assign micromatrizz[58][102] = 9'b111111111;
assign micromatrizz[58][103] = 9'b111111111;
assign micromatrizz[58][104] = 9'b111110010;
assign micromatrizz[58][105] = 9'b111110010;
assign micromatrizz[58][106] = 9'b111110010;
assign micromatrizz[58][107] = 9'b111110010;
assign micromatrizz[58][108] = 9'b111110011;
assign micromatrizz[58][109] = 9'b111110011;
assign micromatrizz[58][110] = 9'b111110011;
assign micromatrizz[58][111] = 9'b111110011;
assign micromatrizz[58][112] = 9'b111110011;
assign micromatrizz[58][113] = 9'b111111111;
assign micromatrizz[58][114] = 9'b111111111;
assign micromatrizz[58][115] = 9'b111111111;
assign micromatrizz[58][116] = 9'b111111111;
assign micromatrizz[58][117] = 9'b111111111;
assign micromatrizz[58][118] = 9'b111111111;
assign micromatrizz[58][119] = 9'b111110110;
assign micromatrizz[58][120] = 9'b111110010;
assign micromatrizz[58][121] = 9'b111110010;
assign micromatrizz[58][122] = 9'b111110010;
assign micromatrizz[58][123] = 9'b111110010;
assign micromatrizz[58][124] = 9'b111110011;
assign micromatrizz[58][125] = 9'b111110011;
assign micromatrizz[58][126] = 9'b111110011;
assign micromatrizz[58][127] = 9'b111111111;
assign micromatrizz[58][128] = 9'b111111111;
assign micromatrizz[58][129] = 9'b111111111;
assign micromatrizz[58][130] = 9'b111111111;
assign micromatrizz[58][131] = 9'b111111111;
assign micromatrizz[58][132] = 9'b111111111;
assign micromatrizz[58][133] = 9'b111111111;
assign micromatrizz[58][134] = 9'b111110110;
assign micromatrizz[58][135] = 9'b111111111;
assign micromatrizz[58][136] = 9'b111111111;
assign micromatrizz[58][137] = 9'b111111111;
assign micromatrizz[58][138] = 9'b111110111;
assign micromatrizz[58][139] = 9'b111110010;
assign micromatrizz[58][140] = 9'b111110010;
assign micromatrizz[58][141] = 9'b111110010;
assign micromatrizz[58][142] = 9'b111110010;
assign micromatrizz[58][143] = 9'b111110011;
assign micromatrizz[58][144] = 9'b111110011;
assign micromatrizz[58][145] = 9'b111110011;
assign micromatrizz[58][146] = 9'b111111111;
assign micromatrizz[58][147] = 9'b111111111;
assign micromatrizz[58][148] = 9'b111111111;
assign micromatrizz[58][149] = 9'b111111111;
assign micromatrizz[58][150] = 9'b111110111;
assign micromatrizz[58][151] = 9'b111110010;
assign micromatrizz[58][152] = 9'b111110011;
assign micromatrizz[58][153] = 9'b111110011;
assign micromatrizz[58][154] = 9'b111110011;
assign micromatrizz[58][155] = 9'b111110011;
assign micromatrizz[58][156] = 9'b111110011;
assign micromatrizz[58][157] = 9'b111110011;
assign micromatrizz[58][158] = 9'b111111111;
assign micromatrizz[58][159] = 9'b111111111;
assign micromatrizz[58][160] = 9'b111111111;
assign micromatrizz[58][161] = 9'b111111111;
assign micromatrizz[58][162] = 9'b111111111;
assign micromatrizz[58][163] = 9'b111111111;
assign micromatrizz[58][164] = 9'b111111111;
assign micromatrizz[58][165] = 9'b111111111;
assign micromatrizz[58][166] = 9'b111111111;
assign micromatrizz[58][167] = 9'b111111111;
assign micromatrizz[58][168] = 9'b111111111;
assign micromatrizz[58][169] = 9'b111111111;
assign micromatrizz[58][170] = 9'b111111111;
assign micromatrizz[58][171] = 9'b111111111;
assign micromatrizz[58][172] = 9'b111110010;
assign micromatrizz[58][173] = 9'b111110010;
assign micromatrizz[58][174] = 9'b111110010;
assign micromatrizz[58][175] = 9'b111110011;
assign micromatrizz[58][176] = 9'b111110011;
assign micromatrizz[58][177] = 9'b111110011;
assign micromatrizz[58][178] = 9'b111110011;
assign micromatrizz[58][179] = 9'b111110111;
assign micromatrizz[58][180] = 9'b111111111;
assign micromatrizz[58][181] = 9'b111111111;
assign micromatrizz[58][182] = 9'b111111111;
assign micromatrizz[58][183] = 9'b111110010;
assign micromatrizz[58][184] = 9'b111110010;
assign micromatrizz[58][185] = 9'b111110010;
assign micromatrizz[58][186] = 9'b111110010;
assign micromatrizz[58][187] = 9'b111110011;
assign micromatrizz[58][188] = 9'b111110010;
assign micromatrizz[58][189] = 9'b111110011;
assign micromatrizz[58][190] = 9'b111111111;
assign micromatrizz[58][191] = 9'b111111111;
assign micromatrizz[58][192] = 9'b111111111;
assign micromatrizz[58][193] = 9'b111111111;
assign micromatrizz[58][194] = 9'b111111111;
assign micromatrizz[58][195] = 9'b111110010;
assign micromatrizz[58][196] = 9'b111110010;
assign micromatrizz[58][197] = 9'b111110011;
assign micromatrizz[58][198] = 9'b111110011;
assign micromatrizz[58][199] = 9'b111110010;
assign micromatrizz[58][200] = 9'b111110010;
assign micromatrizz[58][201] = 9'b111110011;
assign micromatrizz[58][202] = 9'b111110111;
assign micromatrizz[58][203] = 9'b111111111;
assign micromatrizz[58][204] = 9'b111111111;
assign micromatrizz[58][205] = 9'b111111111;
assign micromatrizz[58][206] = 9'b111110010;
assign micromatrizz[58][207] = 9'b111110010;
assign micromatrizz[58][208] = 9'b111110010;
assign micromatrizz[58][209] = 9'b111110010;
assign micromatrizz[58][210] = 9'b111110011;
assign micromatrizz[58][211] = 9'b111110011;
assign micromatrizz[58][212] = 9'b111110011;
assign micromatrizz[58][213] = 9'b111110111;
assign micromatrizz[58][214] = 9'b111111111;
assign micromatrizz[58][215] = 9'b111111111;
assign micromatrizz[58][216] = 9'b111111111;
assign micromatrizz[58][217] = 9'b111111111;
assign micromatrizz[58][218] = 9'b111111111;
assign micromatrizz[58][219] = 9'b111111111;
assign micromatrizz[58][220] = 9'b111111111;
assign micromatrizz[58][221] = 9'b111110010;
assign micromatrizz[58][222] = 9'b111111111;
assign micromatrizz[58][223] = 9'b111111111;
assign micromatrizz[58][224] = 9'b111111111;
assign micromatrizz[58][225] = 9'b111110110;
assign micromatrizz[58][226] = 9'b111110010;
assign micromatrizz[58][227] = 9'b111110010;
assign micromatrizz[58][228] = 9'b111110010;
assign micromatrizz[58][229] = 9'b111110010;
assign micromatrizz[58][230] = 9'b111110011;
assign micromatrizz[58][231] = 9'b111110010;
assign micromatrizz[58][232] = 9'b111110111;
assign micromatrizz[58][233] = 9'b111111111;
assign micromatrizz[58][234] = 9'b111111111;
assign micromatrizz[58][235] = 9'b111111111;
assign micromatrizz[58][236] = 9'b111111111;
assign micromatrizz[58][237] = 9'b111111111;
assign micromatrizz[58][238] = 9'b111111111;
assign micromatrizz[58][239] = 9'b111111111;
assign micromatrizz[58][240] = 9'b111111111;
assign micromatrizz[58][241] = 9'b111110111;
assign micromatrizz[58][242] = 9'b111110010;
assign micromatrizz[58][243] = 9'b111110010;
assign micromatrizz[58][244] = 9'b111110011;
assign micromatrizz[58][245] = 9'b111110011;
assign micromatrizz[58][246] = 9'b111110011;
assign micromatrizz[58][247] = 9'b111110111;
assign micromatrizz[58][248] = 9'b111111111;
assign micromatrizz[58][249] = 9'b111111111;
assign micromatrizz[58][250] = 9'b111111111;
assign micromatrizz[58][251] = 9'b111110110;
assign micromatrizz[58][252] = 9'b111110010;
assign micromatrizz[58][253] = 9'b111110010;
assign micromatrizz[58][254] = 9'b111110011;
assign micromatrizz[58][255] = 9'b111110011;
assign micromatrizz[58][256] = 9'b111110010;
assign micromatrizz[58][257] = 9'b111111111;
assign micromatrizz[58][258] = 9'b111111111;
assign micromatrizz[58][259] = 9'b111110111;
assign micromatrizz[58][260] = 9'b111110010;
assign micromatrizz[58][261] = 9'b111110010;
assign micromatrizz[58][262] = 9'b111110011;
assign micromatrizz[58][263] = 9'b111110011;
assign micromatrizz[58][264] = 9'b111110011;
assign micromatrizz[58][265] = 9'b111110011;
assign micromatrizz[58][266] = 9'b111110011;
assign micromatrizz[58][267] = 9'b111110011;
assign micromatrizz[58][268] = 9'b111110111;
assign micromatrizz[58][269] = 9'b111111111;
assign micromatrizz[58][270] = 9'b111111111;
assign micromatrizz[58][271] = 9'b111111111;
assign micromatrizz[58][272] = 9'b111111111;
assign micromatrizz[58][273] = 9'b111111111;
assign micromatrizz[58][274] = 9'b111111111;
assign micromatrizz[58][275] = 9'b111111111;
assign micromatrizz[58][276] = 9'b111111111;
assign micromatrizz[58][277] = 9'b111111111;
assign micromatrizz[58][278] = 9'b111111111;
assign micromatrizz[58][279] = 9'b111111111;
assign micromatrizz[58][280] = 9'b111111111;
assign micromatrizz[58][281] = 9'b111111111;
assign micromatrizz[58][282] = 9'b111111111;
assign micromatrizz[58][283] = 9'b111111111;
assign micromatrizz[58][284] = 9'b111111111;
assign micromatrizz[58][285] = 9'b111111111;
assign micromatrizz[58][286] = 9'b111110010;
assign micromatrizz[58][287] = 9'b111110010;
assign micromatrizz[58][288] = 9'b111110011;
assign micromatrizz[58][289] = 9'b111110010;
assign micromatrizz[58][290] = 9'b111110010;
assign micromatrizz[58][291] = 9'b111110011;
assign micromatrizz[58][292] = 9'b111110010;
assign micromatrizz[58][293] = 9'b111111111;
assign micromatrizz[58][294] = 9'b111111111;
assign micromatrizz[58][295] = 9'b111111111;
assign micromatrizz[58][296] = 9'b111111111;
assign micromatrizz[58][297] = 9'b111111111;
assign micromatrizz[58][298] = 9'b111111111;
assign micromatrizz[58][299] = 9'b111110010;
assign micromatrizz[58][300] = 9'b111110010;
assign micromatrizz[58][301] = 9'b111110010;
assign micromatrizz[58][302] = 9'b111110011;
assign micromatrizz[58][303] = 9'b111110011;
assign micromatrizz[58][304] = 9'b111110011;
assign micromatrizz[58][305] = 9'b111110011;
assign micromatrizz[58][306] = 9'b111110011;
assign micromatrizz[58][307] = 9'b111110111;
assign micromatrizz[58][308] = 9'b111111111;
assign micromatrizz[58][309] = 9'b111111111;
assign micromatrizz[58][310] = 9'b111110111;
assign micromatrizz[58][311] = 9'b111110010;
assign micromatrizz[58][312] = 9'b111111111;
assign micromatrizz[58][313] = 9'b111111111;
assign micromatrizz[58][314] = 9'b111111111;
assign micromatrizz[58][315] = 9'b111111111;
assign micromatrizz[58][316] = 9'b111110010;
assign micromatrizz[58][317] = 9'b111110010;
assign micromatrizz[58][318] = 9'b111110010;
assign micromatrizz[58][319] = 9'b111110010;
assign micromatrizz[58][320] = 9'b111110010;
assign micromatrizz[58][321] = 9'b111110011;
assign micromatrizz[58][322] = 9'b111111111;
assign micromatrizz[58][323] = 9'b111111111;
assign micromatrizz[58][324] = 9'b111111111;
assign micromatrizz[58][325] = 9'b111111111;
assign micromatrizz[58][326] = 9'b111110010;
assign micromatrizz[58][327] = 9'b111110010;
assign micromatrizz[58][328] = 9'b111110010;
assign micromatrizz[58][329] = 9'b111110010;
assign micromatrizz[58][330] = 9'b111110010;
assign micromatrizz[58][331] = 9'b111110111;
assign micromatrizz[58][332] = 9'b111111111;
assign micromatrizz[58][333] = 9'b111111111;
assign micromatrizz[58][334] = 9'b111111111;
assign micromatrizz[58][335] = 9'b111110010;
assign micromatrizz[58][336] = 9'b111110010;
assign micromatrizz[58][337] = 9'b111110011;
assign micromatrizz[58][338] = 9'b111110011;
assign micromatrizz[58][339] = 9'b111110011;
assign micromatrizz[58][340] = 9'b111110011;
assign micromatrizz[58][341] = 9'b111110011;
assign micromatrizz[58][342] = 9'b111111111;
assign micromatrizz[58][343] = 9'b111111111;
assign micromatrizz[58][344] = 9'b111111111;
assign micromatrizz[58][345] = 9'b111111111;
assign micromatrizz[58][346] = 9'b111111111;
assign micromatrizz[58][347] = 9'b111110010;
assign micromatrizz[58][348] = 9'b111110010;
assign micromatrizz[58][349] = 9'b111110010;
assign micromatrizz[58][350] = 9'b111110010;
assign micromatrizz[58][351] = 9'b111110011;
assign micromatrizz[58][352] = 9'b111110011;
assign micromatrizz[58][353] = 9'b111110011;
assign micromatrizz[58][354] = 9'b111111111;
assign micromatrizz[58][355] = 9'b111111111;
assign micromatrizz[58][356] = 9'b111111111;
assign micromatrizz[58][357] = 9'b111111111;
assign micromatrizz[58][358] = 9'b111111111;
assign micromatrizz[58][359] = 9'b111110010;
assign micromatrizz[58][360] = 9'b111110011;
assign micromatrizz[58][361] = 9'b111110010;
assign micromatrizz[58][362] = 9'b111110010;
assign micromatrizz[58][363] = 9'b111110011;
assign micromatrizz[58][364] = 9'b111110011;
assign micromatrizz[58][365] = 9'b111110011;
assign micromatrizz[58][366] = 9'b111111111;
assign micromatrizz[58][367] = 9'b111111111;
assign micromatrizz[58][368] = 9'b111111111;
assign micromatrizz[58][369] = 9'b111111111;
assign micromatrizz[58][370] = 9'b111111111;
assign micromatrizz[58][371] = 9'b111111111;
assign micromatrizz[58][372] = 9'b111110010;
assign micromatrizz[58][373] = 9'b111110011;
assign micromatrizz[58][374] = 9'b111110011;
assign micromatrizz[58][375] = 9'b111110011;
assign micromatrizz[58][376] = 9'b111110011;
assign micromatrizz[58][377] = 9'b111110011;
assign micromatrizz[58][378] = 9'b111110011;
assign micromatrizz[58][379] = 9'b111111111;
assign micromatrizz[58][380] = 9'b111111111;
assign micromatrizz[58][381] = 9'b111111111;
assign micromatrizz[58][382] = 9'b111111111;
assign micromatrizz[58][383] = 9'b111110111;
assign micromatrizz[58][384] = 9'b111110010;
assign micromatrizz[58][385] = 9'b111110010;
assign micromatrizz[58][386] = 9'b111110011;
assign micromatrizz[58][387] = 9'b111110011;
assign micromatrizz[58][388] = 9'b111110011;
assign micromatrizz[58][389] = 9'b111110011;
assign micromatrizz[58][390] = 9'b111110011;
assign micromatrizz[58][391] = 9'b111111111;
assign micromatrizz[58][392] = 9'b111111111;
assign micromatrizz[58][393] = 9'b111111111;
assign micromatrizz[58][394] = 9'b111111111;
assign micromatrizz[58][395] = 9'b111110010;
assign micromatrizz[58][396] = 9'b111110010;
assign micromatrizz[58][397] = 9'b111110010;
assign micromatrizz[58][398] = 9'b111110010;
assign micromatrizz[58][399] = 9'b111110011;
assign micromatrizz[58][400] = 9'b111110011;
assign micromatrizz[58][401] = 9'b111110010;
assign micromatrizz[58][402] = 9'b111110111;
assign micromatrizz[58][403] = 9'b111111111;
assign micromatrizz[58][404] = 9'b111111111;
assign micromatrizz[58][405] = 9'b111111111;
assign micromatrizz[58][406] = 9'b111111111;
assign micromatrizz[58][407] = 9'b111111111;
assign micromatrizz[58][408] = 9'b111111111;
assign micromatrizz[58][409] = 9'b111111111;
assign micromatrizz[58][410] = 9'b111111111;
assign micromatrizz[58][411] = 9'b111110111;
assign micromatrizz[58][412] = 9'b111110010;
assign micromatrizz[58][413] = 9'b111110010;
assign micromatrizz[58][414] = 9'b111110011;
assign micromatrizz[58][415] = 9'b111110011;
assign micromatrizz[58][416] = 9'b111110011;
assign micromatrizz[58][417] = 9'b111110111;
assign micromatrizz[58][418] = 9'b111111111;
assign micromatrizz[58][419] = 9'b111111111;
assign micromatrizz[58][420] = 9'b111111111;
assign micromatrizz[58][421] = 9'b111110111;
assign micromatrizz[58][422] = 9'b111110010;
assign micromatrizz[58][423] = 9'b111110011;
assign micromatrizz[58][424] = 9'b111110011;
assign micromatrizz[58][425] = 9'b111110011;
assign micromatrizz[58][426] = 9'b111110010;
assign micromatrizz[58][427] = 9'b111111111;
assign micromatrizz[58][428] = 9'b111111111;
assign micromatrizz[58][429] = 9'b111111111;
assign micromatrizz[58][430] = 9'b111110111;
assign micromatrizz[58][431] = 9'b111110010;
assign micromatrizz[58][432] = 9'b111110010;
assign micromatrizz[58][433] = 9'b111110010;
assign micromatrizz[58][434] = 9'b111110011;
assign micromatrizz[58][435] = 9'b111110011;
assign micromatrizz[58][436] = 9'b111110011;
assign micromatrizz[58][437] = 9'b111110111;
assign micromatrizz[58][438] = 9'b111111111;
assign micromatrizz[58][439] = 9'b111111111;
assign micromatrizz[58][440] = 9'b111111111;
assign micromatrizz[58][441] = 9'b111111111;
assign micromatrizz[58][442] = 9'b111111111;
assign micromatrizz[58][443] = 9'b111111111;
assign micromatrizz[58][444] = 9'b111111111;
assign micromatrizz[58][445] = 9'b111111111;
assign micromatrizz[58][446] = 9'b111110111;
assign micromatrizz[58][447] = 9'b111110010;
assign micromatrizz[58][448] = 9'b111110010;
assign micromatrizz[58][449] = 9'b111110010;
assign micromatrizz[58][450] = 9'b111110011;
assign micromatrizz[58][451] = 9'b111110011;
assign micromatrizz[58][452] = 9'b111110011;
assign micromatrizz[58][453] = 9'b111110011;
assign micromatrizz[58][454] = 9'b111111111;
assign micromatrizz[58][455] = 9'b111111111;
assign micromatrizz[58][456] = 9'b111111111;
assign micromatrizz[58][457] = 9'b111111111;
assign micromatrizz[58][458] = 9'b111111111;
assign micromatrizz[58][459] = 9'b111111111;
assign micromatrizz[58][460] = 9'b111111111;
assign micromatrizz[58][461] = 9'b111110111;
assign micromatrizz[58][462] = 9'b111111111;
assign micromatrizz[58][463] = 9'b111111111;
assign micromatrizz[58][464] = 9'b111111111;
assign micromatrizz[58][465] = 9'b111110010;
assign micromatrizz[58][466] = 9'b111110010;
assign micromatrizz[58][467] = 9'b111110010;
assign micromatrizz[58][468] = 9'b111110011;
assign micromatrizz[58][469] = 9'b111110011;
assign micromatrizz[58][470] = 9'b111110011;
assign micromatrizz[58][471] = 9'b111110011;
assign micromatrizz[58][472] = 9'b111110011;
assign micromatrizz[58][473] = 9'b111110011;
assign micromatrizz[58][474] = 9'b111111111;
assign micromatrizz[58][475] = 9'b111111111;
assign micromatrizz[58][476] = 9'b111111111;
assign micromatrizz[58][477] = 9'b111111111;
assign micromatrizz[58][478] = 9'b111111111;
assign micromatrizz[58][479] = 9'b111111111;
assign micromatrizz[58][480] = 9'b111111111;
assign micromatrizz[58][481] = 9'b111110010;
assign micromatrizz[58][482] = 9'b111110010;
assign micromatrizz[58][483] = 9'b111110010;
assign micromatrizz[58][484] = 9'b111110010;
assign micromatrizz[58][485] = 9'b111110011;
assign micromatrizz[58][486] = 9'b111110011;
assign micromatrizz[58][487] = 9'b111110011;
assign micromatrizz[58][488] = 9'b111111111;
assign micromatrizz[58][489] = 9'b111111111;
assign micromatrizz[58][490] = 9'b111111111;
assign micromatrizz[58][491] = 9'b111111111;
assign micromatrizz[58][492] = 9'b111111111;
assign micromatrizz[58][493] = 9'b111111111;
assign micromatrizz[58][494] = 9'b111111111;
assign micromatrizz[58][495] = 9'b111111111;
assign micromatrizz[58][496] = 9'b111111111;
assign micromatrizz[58][497] = 9'b111110011;
assign micromatrizz[58][498] = 9'b111110010;
assign micromatrizz[58][499] = 9'b111110011;
assign micromatrizz[58][500] = 9'b111110010;
assign micromatrizz[58][501] = 9'b111110011;
assign micromatrizz[58][502] = 9'b111110010;
assign micromatrizz[58][503] = 9'b111110111;
assign micromatrizz[58][504] = 9'b111111111;
assign micromatrizz[58][505] = 9'b111111111;
assign micromatrizz[58][506] = 9'b111111111;
assign micromatrizz[58][507] = 9'b111110010;
assign micromatrizz[58][508] = 9'b111110010;
assign micromatrizz[58][509] = 9'b111110011;
assign micromatrizz[58][510] = 9'b111110011;
assign micromatrizz[58][511] = 9'b111110011;
assign micromatrizz[58][512] = 9'b111110011;
assign micromatrizz[58][513] = 9'b111111111;
assign micromatrizz[58][514] = 9'b111111111;
assign micromatrizz[58][515] = 9'b111111111;
assign micromatrizz[58][516] = 9'b111110111;
assign micromatrizz[58][517] = 9'b111110011;
assign micromatrizz[58][518] = 9'b111110011;
assign micromatrizz[58][519] = 9'b111110011;
assign micromatrizz[58][520] = 9'b111110010;
assign micromatrizz[58][521] = 9'b111110011;
assign micromatrizz[58][522] = 9'b111110011;
assign micromatrizz[58][523] = 9'b111110111;
assign micromatrizz[58][524] = 9'b111111111;
assign micromatrizz[58][525] = 9'b111111111;
assign micromatrizz[58][526] = 9'b111111111;
assign micromatrizz[58][527] = 9'b111111111;
assign micromatrizz[58][528] = 9'b111110111;
assign micromatrizz[58][529] = 9'b111110010;
assign micromatrizz[58][530] = 9'b111110010;
assign micromatrizz[58][531] = 9'b111110011;
assign micromatrizz[58][532] = 9'b111110011;
assign micromatrizz[58][533] = 9'b111110011;
assign micromatrizz[58][534] = 9'b111110011;
assign micromatrizz[58][535] = 9'b111110010;
assign micromatrizz[58][536] = 9'b111111111;
assign micromatrizz[58][537] = 9'b111111111;
assign micromatrizz[58][538] = 9'b111111111;
assign micromatrizz[58][539] = 9'b111110010;
assign micromatrizz[58][540] = 9'b111110011;
assign micromatrizz[58][541] = 9'b111110011;
assign micromatrizz[58][542] = 9'b111110010;
assign micromatrizz[58][543] = 9'b111110011;
assign micromatrizz[58][544] = 9'b111110010;
assign micromatrizz[58][545] = 9'b111111111;
assign micromatrizz[58][546] = 9'b111111111;
assign micromatrizz[58][547] = 9'b111111111;
assign micromatrizz[58][548] = 9'b111111111;
assign micromatrizz[58][549] = 9'b111110010;
assign micromatrizz[58][550] = 9'b111110010;
assign micromatrizz[58][551] = 9'b111110011;
assign micromatrizz[58][552] = 9'b111110011;
assign micromatrizz[58][553] = 9'b111110011;
assign micromatrizz[58][554] = 9'b111110111;
assign micromatrizz[58][555] = 9'b111111111;
assign micromatrizz[58][556] = 9'b111111111;
assign micromatrizz[58][557] = 9'b111111111;
assign micromatrizz[58][558] = 9'b111110010;
assign micromatrizz[58][559] = 9'b111110010;
assign micromatrizz[58][560] = 9'b111110010;
assign micromatrizz[58][561] = 9'b111110010;
assign micromatrizz[58][562] = 9'b111110011;
assign micromatrizz[58][563] = 9'b111110011;
assign micromatrizz[58][564] = 9'b111110011;
assign micromatrizz[58][565] = 9'b111111111;
assign micromatrizz[58][566] = 9'b111111111;
assign micromatrizz[58][567] = 9'b111111111;
assign micromatrizz[58][568] = 9'b111110111;
assign micromatrizz[58][569] = 9'b111110010;
assign micromatrizz[58][570] = 9'b111110010;
assign micromatrizz[58][571] = 9'b111110010;
assign micromatrizz[58][572] = 9'b111110010;
assign micromatrizz[58][573] = 9'b111110011;
assign micromatrizz[58][574] = 9'b111110011;
assign micromatrizz[58][575] = 9'b111110011;
assign micromatrizz[58][576] = 9'b111111111;
assign micromatrizz[58][577] = 9'b111111111;
assign micromatrizz[58][578] = 9'b111111111;
assign micromatrizz[58][579] = 9'b111111111;
assign micromatrizz[58][580] = 9'b111111111;
assign micromatrizz[58][581] = 9'b111110010;
assign micromatrizz[58][582] = 9'b111110011;
assign micromatrizz[58][583] = 9'b111110011;
assign micromatrizz[58][584] = 9'b111110010;
assign micromatrizz[58][585] = 9'b111110010;
assign micromatrizz[58][586] = 9'b111110011;
assign micromatrizz[58][587] = 9'b111110011;
assign micromatrizz[58][588] = 9'b111111111;
assign micromatrizz[58][589] = 9'b111111111;
assign micromatrizz[58][590] = 9'b111111111;
assign micromatrizz[58][591] = 9'b111111111;
assign micromatrizz[58][592] = 9'b111110010;
assign micromatrizz[58][593] = 9'b111110010;
assign micromatrizz[58][594] = 9'b111110011;
assign micromatrizz[58][595] = 9'b111110011;
assign micromatrizz[58][596] = 9'b111110011;
assign micromatrizz[58][597] = 9'b111110010;
assign micromatrizz[58][598] = 9'b111111111;
assign micromatrizz[58][599] = 9'b111111111;
assign micromatrizz[58][600] = 9'b111111111;
assign micromatrizz[58][601] = 9'b111111111;
assign micromatrizz[58][602] = 9'b111110010;
assign micromatrizz[58][603] = 9'b111110011;
assign micromatrizz[58][604] = 9'b111110011;
assign micromatrizz[58][605] = 9'b111110011;
assign micromatrizz[58][606] = 9'b111110011;
assign micromatrizz[58][607] = 9'b111110111;
assign micromatrizz[58][608] = 9'b111111111;
assign micromatrizz[58][609] = 9'b111111111;
assign micromatrizz[58][610] = 9'b111110011;
assign micromatrizz[58][611] = 9'b111110010;
assign micromatrizz[58][612] = 9'b111110010;
assign micromatrizz[58][613] = 9'b111110010;
assign micromatrizz[58][614] = 9'b111110010;
assign micromatrizz[58][615] = 9'b111110011;
assign micromatrizz[58][616] = 9'b111110011;
assign micromatrizz[58][617] = 9'b111110011;
assign micromatrizz[58][618] = 9'b111110011;
assign micromatrizz[58][619] = 9'b111111111;
assign micromatrizz[58][620] = 9'b111111111;
assign micromatrizz[58][621] = 9'b111111111;
assign micromatrizz[58][622] = 9'b111111111;
assign micromatrizz[58][623] = 9'b111111111;
assign micromatrizz[58][624] = 9'b111111111;
assign micromatrizz[58][625] = 9'b111111111;
assign micromatrizz[58][626] = 9'b111111111;
assign micromatrizz[58][627] = 9'b111111111;
assign micromatrizz[58][628] = 9'b111111111;
assign micromatrizz[58][629] = 9'b111111111;
assign micromatrizz[58][630] = 9'b111111111;
assign micromatrizz[58][631] = 9'b111111111;
assign micromatrizz[58][632] = 9'b111111111;
assign micromatrizz[58][633] = 9'b111111111;
assign micromatrizz[58][634] = 9'b111111111;
assign micromatrizz[58][635] = 9'b111111111;
assign micromatrizz[58][636] = 9'b111111111;
assign micromatrizz[58][637] = 9'b111111111;
assign micromatrizz[58][638] = 9'b111111111;
assign micromatrizz[58][639] = 9'b111111111;
assign micromatrizz[59][0] = 9'b111111111;
assign micromatrizz[59][1] = 9'b111111111;
assign micromatrizz[59][2] = 9'b111111111;
assign micromatrizz[59][3] = 9'b111111111;
assign micromatrizz[59][4] = 9'b111111111;
assign micromatrizz[59][5] = 9'b111111111;
assign micromatrizz[59][6] = 9'b111111111;
assign micromatrizz[59][7] = 9'b111111111;
assign micromatrizz[59][8] = 9'b111110110;
assign micromatrizz[59][9] = 9'b111110010;
assign micromatrizz[59][10] = 9'b111110010;
assign micromatrizz[59][11] = 9'b111110010;
assign micromatrizz[59][12] = 9'b111110010;
assign micromatrizz[59][13] = 9'b111110011;
assign micromatrizz[59][14] = 9'b111110010;
assign micromatrizz[59][15] = 9'b111110011;
assign micromatrizz[59][16] = 9'b111110011;
assign micromatrizz[59][17] = 9'b111110111;
assign micromatrizz[59][18] = 9'b111111111;
assign micromatrizz[59][19] = 9'b111111111;
assign micromatrizz[59][20] = 9'b111111111;
assign micromatrizz[59][21] = 9'b111111111;
assign micromatrizz[59][22] = 9'b111111111;
assign micromatrizz[59][23] = 9'b111110111;
assign micromatrizz[59][24] = 9'b111110010;
assign micromatrizz[59][25] = 9'b111110010;
assign micromatrizz[59][26] = 9'b111110010;
assign micromatrizz[59][27] = 9'b111110011;
assign micromatrizz[59][28] = 9'b111110011;
assign micromatrizz[59][29] = 9'b111110011;
assign micromatrizz[59][30] = 9'b111110011;
assign micromatrizz[59][31] = 9'b111111111;
assign micromatrizz[59][32] = 9'b111111111;
assign micromatrizz[59][33] = 9'b111111111;
assign micromatrizz[59][34] = 9'b111111111;
assign micromatrizz[59][35] = 9'b111110111;
assign micromatrizz[59][36] = 9'b111110010;
assign micromatrizz[59][37] = 9'b111110010;
assign micromatrizz[59][38] = 9'b111110010;
assign micromatrizz[59][39] = 9'b111110011;
assign micromatrizz[59][40] = 9'b111110011;
assign micromatrizz[59][41] = 9'b111110011;
assign micromatrizz[59][42] = 9'b111110011;
assign micromatrizz[59][43] = 9'b111111111;
assign micromatrizz[59][44] = 9'b111111111;
assign micromatrizz[59][45] = 9'b111111111;
assign micromatrizz[59][46] = 9'b111111111;
assign micromatrizz[59][47] = 9'b111110010;
assign micromatrizz[59][48] = 9'b111110010;
assign micromatrizz[59][49] = 9'b111110010;
assign micromatrizz[59][50] = 9'b111110011;
assign micromatrizz[59][51] = 9'b111110011;
assign micromatrizz[59][52] = 9'b111110011;
assign micromatrizz[59][53] = 9'b111110011;
assign micromatrizz[59][54] = 9'b111111111;
assign micromatrizz[59][55] = 9'b111111111;
assign micromatrizz[59][56] = 9'b111111111;
assign micromatrizz[59][57] = 9'b111111111;
assign micromatrizz[59][58] = 9'b111111111;
assign micromatrizz[59][59] = 9'b111110010;
assign micromatrizz[59][60] = 9'b111110010;
assign micromatrizz[59][61] = 9'b111110010;
assign micromatrizz[59][62] = 9'b111110011;
assign micromatrizz[59][63] = 9'b111110011;
assign micromatrizz[59][64] = 9'b111110011;
assign micromatrizz[59][65] = 9'b111110011;
assign micromatrizz[59][66] = 9'b111110111;
assign micromatrizz[59][67] = 9'b111111111;
assign micromatrizz[59][68] = 9'b111110111;
assign micromatrizz[59][69] = 9'b111110010;
assign micromatrizz[59][70] = 9'b111110010;
assign micromatrizz[59][71] = 9'b111110010;
assign micromatrizz[59][72] = 9'b111110011;
assign micromatrizz[59][73] = 9'b111110011;
assign micromatrizz[59][74] = 9'b111110010;
assign micromatrizz[59][75] = 9'b111111111;
assign micromatrizz[59][76] = 9'b111111111;
assign micromatrizz[59][77] = 9'b111111111;
assign micromatrizz[59][78] = 9'b111111111;
assign micromatrizz[59][79] = 9'b111110010;
assign micromatrizz[59][80] = 9'b111110011;
assign micromatrizz[59][81] = 9'b111110011;
assign micromatrizz[59][82] = 9'b111110011;
assign micromatrizz[59][83] = 9'b111110011;
assign micromatrizz[59][84] = 9'b111110011;
assign micromatrizz[59][85] = 9'b111111111;
assign micromatrizz[59][86] = 9'b111111111;
assign micromatrizz[59][87] = 9'b111111111;
assign micromatrizz[59][88] = 9'b111110110;
assign micromatrizz[59][89] = 9'b111110010;
assign micromatrizz[59][90] = 9'b111110010;
assign micromatrizz[59][91] = 9'b111110010;
assign micromatrizz[59][92] = 9'b111110011;
assign micromatrizz[59][93] = 9'b111110011;
assign micromatrizz[59][94] = 9'b111110011;
assign micromatrizz[59][95] = 9'b111110111;
assign micromatrizz[59][96] = 9'b111111111;
assign micromatrizz[59][97] = 9'b111111111;
assign micromatrizz[59][98] = 9'b111111111;
assign micromatrizz[59][99] = 9'b111111111;
assign micromatrizz[59][100] = 9'b111111111;
assign micromatrizz[59][101] = 9'b111111111;
assign micromatrizz[59][102] = 9'b111111111;
assign micromatrizz[59][103] = 9'b111111111;
assign micromatrizz[59][104] = 9'b111110111;
assign micromatrizz[59][105] = 9'b111110010;
assign micromatrizz[59][106] = 9'b111110010;
assign micromatrizz[59][107] = 9'b111110010;
assign micromatrizz[59][108] = 9'b111110010;
assign micromatrizz[59][109] = 9'b111110011;
assign micromatrizz[59][110] = 9'b111110010;
assign micromatrizz[59][111] = 9'b111110011;
assign micromatrizz[59][112] = 9'b111110011;
assign micromatrizz[59][113] = 9'b111110010;
assign micromatrizz[59][114] = 9'b111111111;
assign micromatrizz[59][115] = 9'b111111111;
assign micromatrizz[59][116] = 9'b111111111;
assign micromatrizz[59][117] = 9'b111111111;
assign micromatrizz[59][118] = 9'b111111111;
assign micromatrizz[59][119] = 9'b111110010;
assign micromatrizz[59][120] = 9'b111110010;
assign micromatrizz[59][121] = 9'b111110010;
assign micromatrizz[59][122] = 9'b111110010;
assign micromatrizz[59][123] = 9'b111110010;
assign micromatrizz[59][124] = 9'b111110011;
assign micromatrizz[59][125] = 9'b111110011;
assign micromatrizz[59][126] = 9'b111110011;
assign micromatrizz[59][127] = 9'b111111111;
assign micromatrizz[59][128] = 9'b111111111;
assign micromatrizz[59][129] = 9'b111111111;
assign micromatrizz[59][130] = 9'b111111111;
assign micromatrizz[59][131] = 9'b111111111;
assign micromatrizz[59][132] = 9'b111111111;
assign micromatrizz[59][133] = 9'b111111111;
assign micromatrizz[59][134] = 9'b111110111;
assign micromatrizz[59][135] = 9'b111111111;
assign micromatrizz[59][136] = 9'b111111111;
assign micromatrizz[59][137] = 9'b111111111;
assign micromatrizz[59][138] = 9'b111110111;
assign micromatrizz[59][139] = 9'b111110010;
assign micromatrizz[59][140] = 9'b111110010;
assign micromatrizz[59][141] = 9'b111110010;
assign micromatrizz[59][142] = 9'b111110010;
assign micromatrizz[59][143] = 9'b111110011;
assign micromatrizz[59][144] = 9'b111110011;
assign micromatrizz[59][145] = 9'b111110011;
assign micromatrizz[59][146] = 9'b111111111;
assign micromatrizz[59][147] = 9'b111111111;
assign micromatrizz[59][148] = 9'b111111111;
assign micromatrizz[59][149] = 9'b111111111;
assign micromatrizz[59][150] = 9'b111110111;
assign micromatrizz[59][151] = 9'b111110010;
assign micromatrizz[59][152] = 9'b111110011;
assign micromatrizz[59][153] = 9'b111110011;
assign micromatrizz[59][154] = 9'b111110011;
assign micromatrizz[59][155] = 9'b111110011;
assign micromatrizz[59][156] = 9'b111110011;
assign micromatrizz[59][157] = 9'b111110011;
assign micromatrizz[59][158] = 9'b111111111;
assign micromatrizz[59][159] = 9'b111111111;
assign micromatrizz[59][160] = 9'b111111111;
assign micromatrizz[59][161] = 9'b111111111;
assign micromatrizz[59][162] = 9'b111111111;
assign micromatrizz[59][163] = 9'b111110111;
assign micromatrizz[59][164] = 9'b111110111;
assign micromatrizz[59][165] = 9'b111110011;
assign micromatrizz[59][166] = 9'b111110010;
assign micromatrizz[59][167] = 9'b111110010;
assign micromatrizz[59][168] = 9'b111110010;
assign micromatrizz[59][169] = 9'b111110110;
assign micromatrizz[59][170] = 9'b111110111;
assign micromatrizz[59][171] = 9'b111110111;
assign micromatrizz[59][172] = 9'b111110010;
assign micromatrizz[59][173] = 9'b111110010;
assign micromatrizz[59][174] = 9'b111110010;
assign micromatrizz[59][175] = 9'b111110011;
assign micromatrizz[59][176] = 9'b111110011;
assign micromatrizz[59][177] = 9'b111110011;
assign micromatrizz[59][178] = 9'b111110011;
assign micromatrizz[59][179] = 9'b111110111;
assign micromatrizz[59][180] = 9'b111111111;
assign micromatrizz[59][181] = 9'b111111111;
assign micromatrizz[59][182] = 9'b111110111;
assign micromatrizz[59][183] = 9'b111110010;
assign micromatrizz[59][184] = 9'b111110010;
assign micromatrizz[59][185] = 9'b111110011;
assign micromatrizz[59][186] = 9'b111110010;
assign micromatrizz[59][187] = 9'b111110011;
assign micromatrizz[59][188] = 9'b111110011;
assign micromatrizz[59][189] = 9'b111110011;
assign micromatrizz[59][190] = 9'b111111111;
assign micromatrizz[59][191] = 9'b111111111;
assign micromatrizz[59][192] = 9'b111111111;
assign micromatrizz[59][193] = 9'b111111111;
assign micromatrizz[59][194] = 9'b111111111;
assign micromatrizz[59][195] = 9'b111110010;
assign micromatrizz[59][196] = 9'b111110011;
assign micromatrizz[59][197] = 9'b111110011;
assign micromatrizz[59][198] = 9'b111110011;
assign micromatrizz[59][199] = 9'b111110010;
assign micromatrizz[59][200] = 9'b111110010;
assign micromatrizz[59][201] = 9'b111110011;
assign micromatrizz[59][202] = 9'b111110111;
assign micromatrizz[59][203] = 9'b111111111;
assign micromatrizz[59][204] = 9'b111111111;
assign micromatrizz[59][205] = 9'b111111111;
assign micromatrizz[59][206] = 9'b111110010;
assign micromatrizz[59][207] = 9'b111110010;
assign micromatrizz[59][208] = 9'b111110010;
assign micromatrizz[59][209] = 9'b111110011;
assign micromatrizz[59][210] = 9'b111110010;
assign micromatrizz[59][211] = 9'b111110011;
assign micromatrizz[59][212] = 9'b111110011;
assign micromatrizz[59][213] = 9'b111110111;
assign micromatrizz[59][214] = 9'b111111111;
assign micromatrizz[59][215] = 9'b111111111;
assign micromatrizz[59][216] = 9'b111111111;
assign micromatrizz[59][217] = 9'b111111111;
assign micromatrizz[59][218] = 9'b111111111;
assign micromatrizz[59][219] = 9'b111111111;
assign micromatrizz[59][220] = 9'b111111111;
assign micromatrizz[59][221] = 9'b111110110;
assign micromatrizz[59][222] = 9'b111111111;
assign micromatrizz[59][223] = 9'b111111111;
assign micromatrizz[59][224] = 9'b111111111;
assign micromatrizz[59][225] = 9'b111110110;
assign micromatrizz[59][226] = 9'b111110010;
assign micromatrizz[59][227] = 9'b111110010;
assign micromatrizz[59][228] = 9'b111110010;
assign micromatrizz[59][229] = 9'b111110010;
assign micromatrizz[59][230] = 9'b111110011;
assign micromatrizz[59][231] = 9'b111110011;
assign micromatrizz[59][232] = 9'b111110111;
assign micromatrizz[59][233] = 9'b111111111;
assign micromatrizz[59][234] = 9'b111111111;
assign micromatrizz[59][235] = 9'b111111111;
assign micromatrizz[59][236] = 9'b111111111;
assign micromatrizz[59][237] = 9'b111111111;
assign micromatrizz[59][238] = 9'b111111111;
assign micromatrizz[59][239] = 9'b111111111;
assign micromatrizz[59][240] = 9'b111111111;
assign micromatrizz[59][241] = 9'b111110010;
assign micromatrizz[59][242] = 9'b111110010;
assign micromatrizz[59][243] = 9'b111110010;
assign micromatrizz[59][244] = 9'b111110011;
assign micromatrizz[59][245] = 9'b111110011;
assign micromatrizz[59][246] = 9'b111110011;
assign micromatrizz[59][247] = 9'b111110111;
assign micromatrizz[59][248] = 9'b111111111;
assign micromatrizz[59][249] = 9'b111111111;
assign micromatrizz[59][250] = 9'b111111111;
assign micromatrizz[59][251] = 9'b111110110;
assign micromatrizz[59][252] = 9'b111110010;
assign micromatrizz[59][253] = 9'b111110010;
assign micromatrizz[59][254] = 9'b111110010;
assign micromatrizz[59][255] = 9'b111110011;
assign micromatrizz[59][256] = 9'b111110010;
assign micromatrizz[59][257] = 9'b111111111;
assign micromatrizz[59][258] = 9'b111111111;
assign micromatrizz[59][259] = 9'b111111111;
assign micromatrizz[59][260] = 9'b111110010;
assign micromatrizz[59][261] = 9'b111110010;
assign micromatrizz[59][262] = 9'b111110010;
assign micromatrizz[59][263] = 9'b111110010;
assign micromatrizz[59][264] = 9'b111110010;
assign micromatrizz[59][265] = 9'b111110011;
assign micromatrizz[59][266] = 9'b111110011;
assign micromatrizz[59][267] = 9'b111110011;
assign micromatrizz[59][268] = 9'b111110010;
assign micromatrizz[59][269] = 9'b111110111;
assign micromatrizz[59][270] = 9'b111111111;
assign micromatrizz[59][271] = 9'b111111111;
assign micromatrizz[59][272] = 9'b111111111;
assign micromatrizz[59][273] = 9'b111111111;
assign micromatrizz[59][274] = 9'b111111111;
assign micromatrizz[59][275] = 9'b111111111;
assign micromatrizz[59][276] = 9'b111111111;
assign micromatrizz[59][277] = 9'b111111111;
assign micromatrizz[59][278] = 9'b111110111;
assign micromatrizz[59][279] = 9'b111110011;
assign micromatrizz[59][280] = 9'b111110010;
assign micromatrizz[59][281] = 9'b111110010;
assign micromatrizz[59][282] = 9'b111110010;
assign micromatrizz[59][283] = 9'b111110110;
assign micromatrizz[59][284] = 9'b111110111;
assign micromatrizz[59][285] = 9'b111110111;
assign micromatrizz[59][286] = 9'b111110011;
assign micromatrizz[59][287] = 9'b111110010;
assign micromatrizz[59][288] = 9'b111110011;
assign micromatrizz[59][289] = 9'b111110011;
assign micromatrizz[59][290] = 9'b111110011;
assign micromatrizz[59][291] = 9'b111110011;
assign micromatrizz[59][292] = 9'b111110010;
assign micromatrizz[59][293] = 9'b111111111;
assign micromatrizz[59][294] = 9'b111111111;
assign micromatrizz[59][295] = 9'b111111111;
assign micromatrizz[59][296] = 9'b111111111;
assign micromatrizz[59][297] = 9'b111111111;
assign micromatrizz[59][298] = 9'b111111111;
assign micromatrizz[59][299] = 9'b111110111;
assign micromatrizz[59][300] = 9'b111110010;
assign micromatrizz[59][301] = 9'b111110010;
assign micromatrizz[59][302] = 9'b111110011;
assign micromatrizz[59][303] = 9'b111110010;
assign micromatrizz[59][304] = 9'b111110011;
assign micromatrizz[59][305] = 9'b111110011;
assign micromatrizz[59][306] = 9'b111110011;
assign micromatrizz[59][307] = 9'b111110011;
assign micromatrizz[59][308] = 9'b111111111;
assign micromatrizz[59][309] = 9'b111111111;
assign micromatrizz[59][310] = 9'b111110010;
assign micromatrizz[59][311] = 9'b111111111;
assign micromatrizz[59][312] = 9'b111111111;
assign micromatrizz[59][313] = 9'b111111111;
assign micromatrizz[59][314] = 9'b111111111;
assign micromatrizz[59][315] = 9'b111110111;
assign micromatrizz[59][316] = 9'b111110010;
assign micromatrizz[59][317] = 9'b111110010;
assign micromatrizz[59][318] = 9'b111110011;
assign micromatrizz[59][319] = 9'b111110010;
assign micromatrizz[59][320] = 9'b111110011;
assign micromatrizz[59][321] = 9'b111110010;
assign micromatrizz[59][322] = 9'b111111111;
assign micromatrizz[59][323] = 9'b111111111;
assign micromatrizz[59][324] = 9'b111111111;
assign micromatrizz[59][325] = 9'b111111111;
assign micromatrizz[59][326] = 9'b111110010;
assign micromatrizz[59][327] = 9'b111110011;
assign micromatrizz[59][328] = 9'b111110011;
assign micromatrizz[59][329] = 9'b111110011;
assign micromatrizz[59][330] = 9'b111110011;
assign micromatrizz[59][331] = 9'b111110011;
assign micromatrizz[59][332] = 9'b111111111;
assign micromatrizz[59][333] = 9'b111111111;
assign micromatrizz[59][334] = 9'b111111111;
assign micromatrizz[59][335] = 9'b111110010;
assign micromatrizz[59][336] = 9'b111110010;
assign micromatrizz[59][337] = 9'b111110011;
assign micromatrizz[59][338] = 9'b111110011;
assign micromatrizz[59][339] = 9'b111110011;
assign micromatrizz[59][340] = 9'b111110011;
assign micromatrizz[59][341] = 9'b111110011;
assign micromatrizz[59][342] = 9'b111110111;
assign micromatrizz[59][343] = 9'b111111111;
assign micromatrizz[59][344] = 9'b111111111;
assign micromatrizz[59][345] = 9'b111111111;
assign micromatrizz[59][346] = 9'b111111111;
assign micromatrizz[59][347] = 9'b111110010;
assign micromatrizz[59][348] = 9'b111110010;
assign micromatrizz[59][349] = 9'b111110010;
assign micromatrizz[59][350] = 9'b111110011;
assign micromatrizz[59][351] = 9'b111110011;
assign micromatrizz[59][352] = 9'b111110011;
assign micromatrizz[59][353] = 9'b111110011;
assign micromatrizz[59][354] = 9'b111111111;
assign micromatrizz[59][355] = 9'b111111111;
assign micromatrizz[59][356] = 9'b111111111;
assign micromatrizz[59][357] = 9'b111111111;
assign micromatrizz[59][358] = 9'b111111111;
assign micromatrizz[59][359] = 9'b111110010;
assign micromatrizz[59][360] = 9'b111110011;
assign micromatrizz[59][361] = 9'b111110010;
assign micromatrizz[59][362] = 9'b111110010;
assign micromatrizz[59][363] = 9'b111110011;
assign micromatrizz[59][364] = 9'b111110011;
assign micromatrizz[59][365] = 9'b111110011;
assign micromatrizz[59][366] = 9'b111111111;
assign micromatrizz[59][367] = 9'b111111111;
assign micromatrizz[59][368] = 9'b111111111;
assign micromatrizz[59][369] = 9'b111111111;
assign micromatrizz[59][370] = 9'b111111111;
assign micromatrizz[59][371] = 9'b111111111;
assign micromatrizz[59][372] = 9'b111110010;
assign micromatrizz[59][373] = 9'b111110010;
assign micromatrizz[59][374] = 9'b111110011;
assign micromatrizz[59][375] = 9'b111110011;
assign micromatrizz[59][376] = 9'b111110011;
assign micromatrizz[59][377] = 9'b111110011;
assign micromatrizz[59][378] = 9'b111110011;
assign micromatrizz[59][379] = 9'b111111111;
assign micromatrizz[59][380] = 9'b111111111;
assign micromatrizz[59][381] = 9'b111111111;
assign micromatrizz[59][382] = 9'b111111111;
assign micromatrizz[59][383] = 9'b111110111;
assign micromatrizz[59][384] = 9'b111110010;
assign micromatrizz[59][385] = 9'b111110010;
assign micromatrizz[59][386] = 9'b111110011;
assign micromatrizz[59][387] = 9'b111110011;
assign micromatrizz[59][388] = 9'b111110011;
assign micromatrizz[59][389] = 9'b111110011;
assign micromatrizz[59][390] = 9'b111110011;
assign micromatrizz[59][391] = 9'b111111111;
assign micromatrizz[59][392] = 9'b111111111;
assign micromatrizz[59][393] = 9'b111111111;
assign micromatrizz[59][394] = 9'b111111111;
assign micromatrizz[59][395] = 9'b111110010;
assign micromatrizz[59][396] = 9'b111110010;
assign micromatrizz[59][397] = 9'b111110010;
assign micromatrizz[59][398] = 9'b111110010;
assign micromatrizz[59][399] = 9'b111110011;
assign micromatrizz[59][400] = 9'b111110011;
assign micromatrizz[59][401] = 9'b111110010;
assign micromatrizz[59][402] = 9'b111110111;
assign micromatrizz[59][403] = 9'b111111111;
assign micromatrizz[59][404] = 9'b111111111;
assign micromatrizz[59][405] = 9'b111111111;
assign micromatrizz[59][406] = 9'b111111111;
assign micromatrizz[59][407] = 9'b111111111;
assign micromatrizz[59][408] = 9'b111111111;
assign micromatrizz[59][409] = 9'b111111111;
assign micromatrizz[59][410] = 9'b111111111;
assign micromatrizz[59][411] = 9'b111110010;
assign micromatrizz[59][412] = 9'b111110010;
assign micromatrizz[59][413] = 9'b111110010;
assign micromatrizz[59][414] = 9'b111110011;
assign micromatrizz[59][415] = 9'b111110011;
assign micromatrizz[59][416] = 9'b111110011;
assign micromatrizz[59][417] = 9'b111110111;
assign micromatrizz[59][418] = 9'b111111111;
assign micromatrizz[59][419] = 9'b111111111;
assign micromatrizz[59][420] = 9'b111111111;
assign micromatrizz[59][421] = 9'b111110111;
assign micromatrizz[59][422] = 9'b111110010;
assign micromatrizz[59][423] = 9'b111110010;
assign micromatrizz[59][424] = 9'b111110011;
assign micromatrizz[59][425] = 9'b111110011;
assign micromatrizz[59][426] = 9'b111110010;
assign micromatrizz[59][427] = 9'b111111111;
assign micromatrizz[59][428] = 9'b111111111;
assign micromatrizz[59][429] = 9'b111111111;
assign micromatrizz[59][430] = 9'b111110111;
assign micromatrizz[59][431] = 9'b111110010;
assign micromatrizz[59][432] = 9'b111110010;
assign micromatrizz[59][433] = 9'b111110010;
assign micromatrizz[59][434] = 9'b111110011;
assign micromatrizz[59][435] = 9'b111110011;
assign micromatrizz[59][436] = 9'b111110011;
assign micromatrizz[59][437] = 9'b111110111;
assign micromatrizz[59][438] = 9'b111111111;
assign micromatrizz[59][439] = 9'b111111111;
assign micromatrizz[59][440] = 9'b111111111;
assign micromatrizz[59][441] = 9'b111111111;
assign micromatrizz[59][442] = 9'b111111111;
assign micromatrizz[59][443] = 9'b111111111;
assign micromatrizz[59][444] = 9'b111111111;
assign micromatrizz[59][445] = 9'b111111111;
assign micromatrizz[59][446] = 9'b111110010;
assign micromatrizz[59][447] = 9'b111110010;
assign micromatrizz[59][448] = 9'b111110010;
assign micromatrizz[59][449] = 9'b111110010;
assign micromatrizz[59][450] = 9'b111110010;
assign micromatrizz[59][451] = 9'b111110011;
assign micromatrizz[59][452] = 9'b111110011;
assign micromatrizz[59][453] = 9'b111110011;
assign micromatrizz[59][454] = 9'b111111111;
assign micromatrizz[59][455] = 9'b111111111;
assign micromatrizz[59][456] = 9'b111111111;
assign micromatrizz[59][457] = 9'b111111111;
assign micromatrizz[59][458] = 9'b111111111;
assign micromatrizz[59][459] = 9'b111111111;
assign micromatrizz[59][460] = 9'b111111111;
assign micromatrizz[59][461] = 9'b111111111;
assign micromatrizz[59][462] = 9'b111110111;
assign micromatrizz[59][463] = 9'b111111111;
assign micromatrizz[59][464] = 9'b111111111;
assign micromatrizz[59][465] = 9'b111110111;
assign micromatrizz[59][466] = 9'b111110010;
assign micromatrizz[59][467] = 9'b111110010;
assign micromatrizz[59][468] = 9'b111110010;
assign micromatrizz[59][469] = 9'b111110010;
assign micromatrizz[59][470] = 9'b111110010;
assign micromatrizz[59][471] = 9'b111110011;
assign micromatrizz[59][472] = 9'b111110011;
assign micromatrizz[59][473] = 9'b111110011;
assign micromatrizz[59][474] = 9'b111110011;
assign micromatrizz[59][475] = 9'b111111111;
assign micromatrizz[59][476] = 9'b111111111;
assign micromatrizz[59][477] = 9'b111111111;
assign micromatrizz[59][478] = 9'b111111111;
assign micromatrizz[59][479] = 9'b111111111;
assign micromatrizz[59][480] = 9'b111111111;
assign micromatrizz[59][481] = 9'b111110110;
assign micromatrizz[59][482] = 9'b111110010;
assign micromatrizz[59][483] = 9'b111110010;
assign micromatrizz[59][484] = 9'b111110010;
assign micromatrizz[59][485] = 9'b111110011;
assign micromatrizz[59][486] = 9'b111110011;
assign micromatrizz[59][487] = 9'b111110010;
assign micromatrizz[59][488] = 9'b111110111;
assign micromatrizz[59][489] = 9'b111111111;
assign micromatrizz[59][490] = 9'b111111111;
assign micromatrizz[59][491] = 9'b111111111;
assign micromatrizz[59][492] = 9'b111111111;
assign micromatrizz[59][493] = 9'b111111111;
assign micromatrizz[59][494] = 9'b111111111;
assign micromatrizz[59][495] = 9'b111111111;
assign micromatrizz[59][496] = 9'b111111111;
assign micromatrizz[59][497] = 9'b111110010;
assign micromatrizz[59][498] = 9'b111110010;
assign micromatrizz[59][499] = 9'b111110011;
assign micromatrizz[59][500] = 9'b111110010;
assign micromatrizz[59][501] = 9'b111110011;
assign micromatrizz[59][502] = 9'b111110010;
assign micromatrizz[59][503] = 9'b111110111;
assign micromatrizz[59][504] = 9'b111111111;
assign micromatrizz[59][505] = 9'b111111111;
assign micromatrizz[59][506] = 9'b111111111;
assign micromatrizz[59][507] = 9'b111110010;
assign micromatrizz[59][508] = 9'b111110010;
assign micromatrizz[59][509] = 9'b111110010;
assign micromatrizz[59][510] = 9'b111110011;
assign micromatrizz[59][511] = 9'b111110011;
assign micromatrizz[59][512] = 9'b111110011;
assign micromatrizz[59][513] = 9'b111111111;
assign micromatrizz[59][514] = 9'b111111111;
assign micromatrizz[59][515] = 9'b111111111;
assign micromatrizz[59][516] = 9'b111110111;
assign micromatrizz[59][517] = 9'b111110011;
assign micromatrizz[59][518] = 9'b111110011;
assign micromatrizz[59][519] = 9'b111110011;
assign micromatrizz[59][520] = 9'b111110010;
assign micromatrizz[59][521] = 9'b111110010;
assign micromatrizz[59][522] = 9'b111110011;
assign micromatrizz[59][523] = 9'b111110111;
assign micromatrizz[59][524] = 9'b111111111;
assign micromatrizz[59][525] = 9'b111111111;
assign micromatrizz[59][526] = 9'b111111111;
assign micromatrizz[59][527] = 9'b111111111;
assign micromatrizz[59][528] = 9'b111110111;
assign micromatrizz[59][529] = 9'b111110010;
assign micromatrizz[59][530] = 9'b111110010;
assign micromatrizz[59][531] = 9'b111110010;
assign micromatrizz[59][532] = 9'b111110011;
assign micromatrizz[59][533] = 9'b111110011;
assign micromatrizz[59][534] = 9'b111110011;
assign micromatrizz[59][535] = 9'b111110010;
assign micromatrizz[59][536] = 9'b111111111;
assign micromatrizz[59][537] = 9'b111111111;
assign micromatrizz[59][538] = 9'b111110111;
assign micromatrizz[59][539] = 9'b111110010;
assign micromatrizz[59][540] = 9'b111110010;
assign micromatrizz[59][541] = 9'b111110010;
assign micromatrizz[59][542] = 9'b111110011;
assign micromatrizz[59][543] = 9'b111110011;
assign micromatrizz[59][544] = 9'b111110010;
assign micromatrizz[59][545] = 9'b111111111;
assign micromatrizz[59][546] = 9'b111111111;
assign micromatrizz[59][547] = 9'b111111111;
assign micromatrizz[59][548] = 9'b111111111;
assign micromatrizz[59][549] = 9'b111110010;
assign micromatrizz[59][550] = 9'b111110011;
assign micromatrizz[59][551] = 9'b111110011;
assign micromatrizz[59][552] = 9'b111110011;
assign micromatrizz[59][553] = 9'b111110010;
assign micromatrizz[59][554] = 9'b111110111;
assign micromatrizz[59][555] = 9'b111111111;
assign micromatrizz[59][556] = 9'b111111111;
assign micromatrizz[59][557] = 9'b111111111;
assign micromatrizz[59][558] = 9'b111110010;
assign micromatrizz[59][559] = 9'b111110010;
assign micromatrizz[59][560] = 9'b111110010;
assign micromatrizz[59][561] = 9'b111110010;
assign micromatrizz[59][562] = 9'b111110011;
assign micromatrizz[59][563] = 9'b111110011;
assign micromatrizz[59][564] = 9'b111110010;
assign micromatrizz[59][565] = 9'b111111111;
assign micromatrizz[59][566] = 9'b111111111;
assign micromatrizz[59][567] = 9'b111111111;
assign micromatrizz[59][568] = 9'b111110111;
assign micromatrizz[59][569] = 9'b111110010;
assign micromatrizz[59][570] = 9'b111110010;
assign micromatrizz[59][571] = 9'b111110010;
assign micromatrizz[59][572] = 9'b111110011;
assign micromatrizz[59][573] = 9'b111110011;
assign micromatrizz[59][574] = 9'b111110011;
assign micromatrizz[59][575] = 9'b111110011;
assign micromatrizz[59][576] = 9'b111111111;
assign micromatrizz[59][577] = 9'b111111111;
assign micromatrizz[59][578] = 9'b111111111;
assign micromatrizz[59][579] = 9'b111111111;
assign micromatrizz[59][580] = 9'b111111111;
assign micromatrizz[59][581] = 9'b111110010;
assign micromatrizz[59][582] = 9'b111110011;
assign micromatrizz[59][583] = 9'b111110011;
assign micromatrizz[59][584] = 9'b111110010;
assign micromatrizz[59][585] = 9'b111110011;
assign micromatrizz[59][586] = 9'b111110011;
assign micromatrizz[59][587] = 9'b111110011;
assign micromatrizz[59][588] = 9'b111111111;
assign micromatrizz[59][589] = 9'b111111111;
assign micromatrizz[59][590] = 9'b111111111;
assign micromatrizz[59][591] = 9'b111110111;
assign micromatrizz[59][592] = 9'b111110010;
assign micromatrizz[59][593] = 9'b111110010;
assign micromatrizz[59][594] = 9'b111110011;
assign micromatrizz[59][595] = 9'b111110011;
assign micromatrizz[59][596] = 9'b111110011;
assign micromatrizz[59][597] = 9'b111110011;
assign micromatrizz[59][598] = 9'b111111111;
assign micromatrizz[59][599] = 9'b111111111;
assign micromatrizz[59][600] = 9'b111111111;
assign micromatrizz[59][601] = 9'b111111111;
assign micromatrizz[59][602] = 9'b111110010;
assign micromatrizz[59][603] = 9'b111110011;
assign micromatrizz[59][604] = 9'b111110011;
assign micromatrizz[59][605] = 9'b111110011;
assign micromatrizz[59][606] = 9'b111110011;
assign micromatrizz[59][607] = 9'b111110111;
assign micromatrizz[59][608] = 9'b111111111;
assign micromatrizz[59][609] = 9'b111111111;
assign micromatrizz[59][610] = 9'b111110111;
assign micromatrizz[59][611] = 9'b111110010;
assign micromatrizz[59][612] = 9'b111110011;
assign micromatrizz[59][613] = 9'b111110010;
assign micromatrizz[59][614] = 9'b111110010;
assign micromatrizz[59][615] = 9'b111110011;
assign micromatrizz[59][616] = 9'b111110011;
assign micromatrizz[59][617] = 9'b111110011;
assign micromatrizz[59][618] = 9'b111110011;
assign micromatrizz[59][619] = 9'b111110011;
assign micromatrizz[59][620] = 9'b111111111;
assign micromatrizz[59][621] = 9'b111111111;
assign micromatrizz[59][622] = 9'b111111111;
assign micromatrizz[59][623] = 9'b111111111;
assign micromatrizz[59][624] = 9'b111111111;
assign micromatrizz[59][625] = 9'b111111111;
assign micromatrizz[59][626] = 9'b111111111;
assign micromatrizz[59][627] = 9'b111111111;
assign micromatrizz[59][628] = 9'b111111111;
assign micromatrizz[59][629] = 9'b111111111;
assign micromatrizz[59][630] = 9'b111111111;
assign micromatrizz[59][631] = 9'b111111111;
assign micromatrizz[59][632] = 9'b111111111;
assign micromatrizz[59][633] = 9'b111111111;
assign micromatrizz[59][634] = 9'b111111111;
assign micromatrizz[59][635] = 9'b111111111;
assign micromatrizz[59][636] = 9'b111111111;
assign micromatrizz[59][637] = 9'b111111111;
assign micromatrizz[59][638] = 9'b111111111;
assign micromatrizz[59][639] = 9'b111111111;
assign micromatrizz[60][0] = 9'b111111111;
assign micromatrizz[60][1] = 9'b111111111;
assign micromatrizz[60][2] = 9'b111111111;
assign micromatrizz[60][3] = 9'b111111111;
assign micromatrizz[60][4] = 9'b111111111;
assign micromatrizz[60][5] = 9'b111111111;
assign micromatrizz[60][6] = 9'b111111111;
assign micromatrizz[60][7] = 9'b111111111;
assign micromatrizz[60][8] = 9'b111110111;
assign micromatrizz[60][9] = 9'b111110010;
assign micromatrizz[60][10] = 9'b111110010;
assign micromatrizz[60][11] = 9'b111110010;
assign micromatrizz[60][12] = 9'b111110010;
assign micromatrizz[60][13] = 9'b111110010;
assign micromatrizz[60][14] = 9'b111110010;
assign micromatrizz[60][15] = 9'b111110010;
assign micromatrizz[60][16] = 9'b111110011;
assign micromatrizz[60][17] = 9'b111110010;
assign micromatrizz[60][18] = 9'b111110111;
assign micromatrizz[60][19] = 9'b111111111;
assign micromatrizz[60][20] = 9'b111111111;
assign micromatrizz[60][21] = 9'b111111111;
assign micromatrizz[60][22] = 9'b111111111;
assign micromatrizz[60][23] = 9'b111111111;
assign micromatrizz[60][24] = 9'b111110010;
assign micromatrizz[60][25] = 9'b111110010;
assign micromatrizz[60][26] = 9'b111110010;
assign micromatrizz[60][27] = 9'b111110011;
assign micromatrizz[60][28] = 9'b111110011;
assign micromatrizz[60][29] = 9'b111110011;
assign micromatrizz[60][30] = 9'b111110011;
assign micromatrizz[60][31] = 9'b111111111;
assign micromatrizz[60][32] = 9'b111111111;
assign micromatrizz[60][33] = 9'b111111111;
assign micromatrizz[60][34] = 9'b111111111;
assign micromatrizz[60][35] = 9'b111110111;
assign micromatrizz[60][36] = 9'b111110010;
assign micromatrizz[60][37] = 9'b111110010;
assign micromatrizz[60][38] = 9'b111110011;
assign micromatrizz[60][39] = 9'b111110011;
assign micromatrizz[60][40] = 9'b111110011;
assign micromatrizz[60][41] = 9'b111110011;
assign micromatrizz[60][42] = 9'b111110011;
assign micromatrizz[60][43] = 9'b111111111;
assign micromatrizz[60][44] = 9'b111111111;
assign micromatrizz[60][45] = 9'b111111111;
assign micromatrizz[60][46] = 9'b111111111;
assign micromatrizz[60][47] = 9'b111110010;
assign micromatrizz[60][48] = 9'b111110010;
assign micromatrizz[60][49] = 9'b111110010;
assign micromatrizz[60][50] = 9'b111110011;
assign micromatrizz[60][51] = 9'b111110011;
assign micromatrizz[60][52] = 9'b111110011;
assign micromatrizz[60][53] = 9'b111110011;
assign micromatrizz[60][54] = 9'b111110111;
assign micromatrizz[60][55] = 9'b111111111;
assign micromatrizz[60][56] = 9'b111111111;
assign micromatrizz[60][57] = 9'b111111111;
assign micromatrizz[60][58] = 9'b111111111;
assign micromatrizz[60][59] = 9'b111110010;
assign micromatrizz[60][60] = 9'b111110010;
assign micromatrizz[60][61] = 9'b111110010;
assign micromatrizz[60][62] = 9'b111110011;
assign micromatrizz[60][63] = 9'b111110011;
assign micromatrizz[60][64] = 9'b111110011;
assign micromatrizz[60][65] = 9'b111110011;
assign micromatrizz[60][66] = 9'b111110111;
assign micromatrizz[60][67] = 9'b111111111;
assign micromatrizz[60][68] = 9'b111110111;
assign micromatrizz[60][69] = 9'b111110010;
assign micromatrizz[60][70] = 9'b111110010;
assign micromatrizz[60][71] = 9'b111110010;
assign micromatrizz[60][72] = 9'b111110010;
assign micromatrizz[60][73] = 9'b111110011;
assign micromatrizz[60][74] = 9'b111110011;
assign micromatrizz[60][75] = 9'b111111111;
assign micromatrizz[60][76] = 9'b111111111;
assign micromatrizz[60][77] = 9'b111111111;
assign micromatrizz[60][78] = 9'b111111111;
assign micromatrizz[60][79] = 9'b111110010;
assign micromatrizz[60][80] = 9'b111110010;
assign micromatrizz[60][81] = 9'b111110010;
assign micromatrizz[60][82] = 9'b111110011;
assign micromatrizz[60][83] = 9'b111110011;
assign micromatrizz[60][84] = 9'b111110011;
assign micromatrizz[60][85] = 9'b111111111;
assign micromatrizz[60][86] = 9'b111111111;
assign micromatrizz[60][87] = 9'b111111111;
assign micromatrizz[60][88] = 9'b111110010;
assign micromatrizz[60][89] = 9'b111110010;
assign micromatrizz[60][90] = 9'b111110010;
assign micromatrizz[60][91] = 9'b111110010;
assign micromatrizz[60][92] = 9'b111110011;
assign micromatrizz[60][93] = 9'b111110011;
assign micromatrizz[60][94] = 9'b111110011;
assign micromatrizz[60][95] = 9'b111110111;
assign micromatrizz[60][96] = 9'b111111111;
assign micromatrizz[60][97] = 9'b111111111;
assign micromatrizz[60][98] = 9'b111111111;
assign micromatrizz[60][99] = 9'b111111111;
assign micromatrizz[60][100] = 9'b111111111;
assign micromatrizz[60][101] = 9'b111111111;
assign micromatrizz[60][102] = 9'b111111111;
assign micromatrizz[60][103] = 9'b111111111;
assign micromatrizz[60][104] = 9'b111111111;
assign micromatrizz[60][105] = 9'b111110010;
assign micromatrizz[60][106] = 9'b111110010;
assign micromatrizz[60][107] = 9'b111110010;
assign micromatrizz[60][108] = 9'b111110010;
assign micromatrizz[60][109] = 9'b111110010;
assign micromatrizz[60][110] = 9'b111110010;
assign micromatrizz[60][111] = 9'b111110010;
assign micromatrizz[60][112] = 9'b111110011;
assign micromatrizz[60][113] = 9'b111110011;
assign micromatrizz[60][114] = 9'b111110011;
assign micromatrizz[60][115] = 9'b111111111;
assign micromatrizz[60][116] = 9'b111111111;
assign micromatrizz[60][117] = 9'b111111111;
assign micromatrizz[60][118] = 9'b111111111;
assign micromatrizz[60][119] = 9'b111110010;
assign micromatrizz[60][120] = 9'b111110010;
assign micromatrizz[60][121] = 9'b111110010;
assign micromatrizz[60][122] = 9'b111110010;
assign micromatrizz[60][123] = 9'b111110010;
assign micromatrizz[60][124] = 9'b111110011;
assign micromatrizz[60][125] = 9'b111110011;
assign micromatrizz[60][126] = 9'b111110011;
assign micromatrizz[60][127] = 9'b111111111;
assign micromatrizz[60][128] = 9'b111111111;
assign micromatrizz[60][129] = 9'b111111111;
assign micromatrizz[60][130] = 9'b111111111;
assign micromatrizz[60][131] = 9'b111111111;
assign micromatrizz[60][132] = 9'b111111111;
assign micromatrizz[60][133] = 9'b111111111;
assign micromatrizz[60][134] = 9'b111110111;
assign micromatrizz[60][135] = 9'b111110111;
assign micromatrizz[60][136] = 9'b111111111;
assign micromatrizz[60][137] = 9'b111111111;
assign micromatrizz[60][138] = 9'b111110111;
assign micromatrizz[60][139] = 9'b111110010;
assign micromatrizz[60][140] = 9'b111110010;
assign micromatrizz[60][141] = 9'b111110010;
assign micromatrizz[60][142] = 9'b111110010;
assign micromatrizz[60][143] = 9'b111110011;
assign micromatrizz[60][144] = 9'b111110011;
assign micromatrizz[60][145] = 9'b111110011;
assign micromatrizz[60][146] = 9'b111111111;
assign micromatrizz[60][147] = 9'b111111111;
assign micromatrizz[60][148] = 9'b111111111;
assign micromatrizz[60][149] = 9'b111111111;
assign micromatrizz[60][150] = 9'b111110111;
assign micromatrizz[60][151] = 9'b111110010;
assign micromatrizz[60][152] = 9'b111110010;
assign micromatrizz[60][153] = 9'b111110010;
assign micromatrizz[60][154] = 9'b111110011;
assign micromatrizz[60][155] = 9'b111110011;
assign micromatrizz[60][156] = 9'b111110011;
assign micromatrizz[60][157] = 9'b111110011;
assign micromatrizz[60][158] = 9'b111111111;
assign micromatrizz[60][159] = 9'b111111111;
assign micromatrizz[60][160] = 9'b111111111;
assign micromatrizz[60][161] = 9'b111111111;
assign micromatrizz[60][162] = 9'b111110111;
assign micromatrizz[60][163] = 9'b111110010;
assign micromatrizz[60][164] = 9'b111110010;
assign micromatrizz[60][165] = 9'b111110010;
assign micromatrizz[60][166] = 9'b111110011;
assign micromatrizz[60][167] = 9'b111110011;
assign micromatrizz[60][168] = 9'b111110111;
assign micromatrizz[60][169] = 9'b111111111;
assign micromatrizz[60][170] = 9'b111111111;
assign micromatrizz[60][171] = 9'b111110010;
assign micromatrizz[60][172] = 9'b111110010;
assign micromatrizz[60][173] = 9'b111110011;
assign micromatrizz[60][174] = 9'b111110011;
assign micromatrizz[60][175] = 9'b111110011;
assign micromatrizz[60][176] = 9'b111110011;
assign micromatrizz[60][177] = 9'b111110011;
assign micromatrizz[60][178] = 9'b111110010;
assign micromatrizz[60][179] = 9'b111110111;
assign micromatrizz[60][180] = 9'b111111111;
assign micromatrizz[60][181] = 9'b111111111;
assign micromatrizz[60][182] = 9'b111110111;
assign micromatrizz[60][183] = 9'b111110010;
assign micromatrizz[60][184] = 9'b111110010;
assign micromatrizz[60][185] = 9'b111110011;
assign micromatrizz[60][186] = 9'b111110010;
assign micromatrizz[60][187] = 9'b111110010;
assign micromatrizz[60][188] = 9'b111110011;
assign micromatrizz[60][189] = 9'b111110011;
assign micromatrizz[60][190] = 9'b111110111;
assign micromatrizz[60][191] = 9'b111111111;
assign micromatrizz[60][192] = 9'b111111111;
assign micromatrizz[60][193] = 9'b111111111;
assign micromatrizz[60][194] = 9'b111111111;
assign micromatrizz[60][195] = 9'b111110010;
assign micromatrizz[60][196] = 9'b111110010;
assign micromatrizz[60][197] = 9'b111110011;
assign micromatrizz[60][198] = 9'b111110011;
assign micromatrizz[60][199] = 9'b111110010;
assign micromatrizz[60][200] = 9'b111110010;
assign micromatrizz[60][201] = 9'b111110011;
assign micromatrizz[60][202] = 9'b111110111;
assign micromatrizz[60][203] = 9'b111111111;
assign micromatrizz[60][204] = 9'b111111111;
assign micromatrizz[60][205] = 9'b111110111;
assign micromatrizz[60][206] = 9'b111110010;
assign micromatrizz[60][207] = 9'b111110010;
assign micromatrizz[60][208] = 9'b111110010;
assign micromatrizz[60][209] = 9'b111110010;
assign micromatrizz[60][210] = 9'b111110011;
assign micromatrizz[60][211] = 9'b111110011;
assign micromatrizz[60][212] = 9'b111110011;
assign micromatrizz[60][213] = 9'b111110111;
assign micromatrizz[60][214] = 9'b111111111;
assign micromatrizz[60][215] = 9'b111111111;
assign micromatrizz[60][216] = 9'b111111111;
assign micromatrizz[60][217] = 9'b111111111;
assign micromatrizz[60][218] = 9'b111111111;
assign micromatrizz[60][219] = 9'b111111111;
assign micromatrizz[60][220] = 9'b111111111;
assign micromatrizz[60][221] = 9'b111110111;
assign micromatrizz[60][222] = 9'b111111111;
assign micromatrizz[60][223] = 9'b111111111;
assign micromatrizz[60][224] = 9'b111111111;
assign micromatrizz[60][225] = 9'b111110010;
assign micromatrizz[60][226] = 9'b111110010;
assign micromatrizz[60][227] = 9'b111110010;
assign micromatrizz[60][228] = 9'b111110010;
assign micromatrizz[60][229] = 9'b111110011;
assign micromatrizz[60][230] = 9'b111110011;
assign micromatrizz[60][231] = 9'b111110011;
assign micromatrizz[60][232] = 9'b111110111;
assign micromatrizz[60][233] = 9'b111111111;
assign micromatrizz[60][234] = 9'b111111111;
assign micromatrizz[60][235] = 9'b111111111;
assign micromatrizz[60][236] = 9'b111111111;
assign micromatrizz[60][237] = 9'b111111111;
assign micromatrizz[60][238] = 9'b111111111;
assign micromatrizz[60][239] = 9'b111111111;
assign micromatrizz[60][240] = 9'b111111111;
assign micromatrizz[60][241] = 9'b111110010;
assign micromatrizz[60][242] = 9'b111110010;
assign micromatrizz[60][243] = 9'b111110010;
assign micromatrizz[60][244] = 9'b111110010;
assign micromatrizz[60][245] = 9'b111110011;
assign micromatrizz[60][246] = 9'b111110011;
assign micromatrizz[60][247] = 9'b111110111;
assign micromatrizz[60][248] = 9'b111111111;
assign micromatrizz[60][249] = 9'b111111111;
assign micromatrizz[60][250] = 9'b111111111;
assign micromatrizz[60][251] = 9'b111110111;
assign micromatrizz[60][252] = 9'b111110010;
assign micromatrizz[60][253] = 9'b111110010;
assign micromatrizz[60][254] = 9'b111110010;
assign micromatrizz[60][255] = 9'b111110011;
assign micromatrizz[60][256] = 9'b111110010;
assign micromatrizz[60][257] = 9'b111111111;
assign micromatrizz[60][258] = 9'b111111111;
assign micromatrizz[60][259] = 9'b111111111;
assign micromatrizz[60][260] = 9'b111110111;
assign micromatrizz[60][261] = 9'b111110010;
assign micromatrizz[60][262] = 9'b111110010;
assign micromatrizz[60][263] = 9'b111110010;
assign micromatrizz[60][264] = 9'b111110010;
assign micromatrizz[60][265] = 9'b111110010;
assign micromatrizz[60][266] = 9'b111110010;
assign micromatrizz[60][267] = 9'b111110011;
assign micromatrizz[60][268] = 9'b111110011;
assign micromatrizz[60][269] = 9'b111110011;
assign micromatrizz[60][270] = 9'b111110111;
assign micromatrizz[60][271] = 9'b111111111;
assign micromatrizz[60][272] = 9'b111111111;
assign micromatrizz[60][273] = 9'b111111111;
assign micromatrizz[60][274] = 9'b111111111;
assign micromatrizz[60][275] = 9'b111111111;
assign micromatrizz[60][276] = 9'b111110111;
assign micromatrizz[60][277] = 9'b111110010;
assign micromatrizz[60][278] = 9'b111110010;
assign micromatrizz[60][279] = 9'b111110011;
assign micromatrizz[60][280] = 9'b111110011;
assign micromatrizz[60][281] = 9'b111110011;
assign micromatrizz[60][282] = 9'b111111111;
assign micromatrizz[60][283] = 9'b111111111;
assign micromatrizz[60][284] = 9'b111111111;
assign micromatrizz[60][285] = 9'b111110010;
assign micromatrizz[60][286] = 9'b111110010;
assign micromatrizz[60][287] = 9'b111110011;
assign micromatrizz[60][288] = 9'b111110011;
assign micromatrizz[60][289] = 9'b111110011;
assign micromatrizz[60][290] = 9'b111110011;
assign micromatrizz[60][291] = 9'b111110011;
assign micromatrizz[60][292] = 9'b111110010;
assign micromatrizz[60][293] = 9'b111111111;
assign micromatrizz[60][294] = 9'b111111111;
assign micromatrizz[60][295] = 9'b111111111;
assign micromatrizz[60][296] = 9'b111111111;
assign micromatrizz[60][297] = 9'b111111111;
assign micromatrizz[60][298] = 9'b111111111;
assign micromatrizz[60][299] = 9'b111111111;
assign micromatrizz[60][300] = 9'b111110010;
assign micromatrizz[60][301] = 9'b111110010;
assign micromatrizz[60][302] = 9'b111110010;
assign micromatrizz[60][303] = 9'b111110010;
assign micromatrizz[60][304] = 9'b111110010;
assign micromatrizz[60][305] = 9'b111110010;
assign micromatrizz[60][306] = 9'b111110011;
assign micromatrizz[60][307] = 9'b111110011;
assign micromatrizz[60][308] = 9'b111110011;
assign micromatrizz[60][309] = 9'b111110111;
assign micromatrizz[60][310] = 9'b111110111;
assign micromatrizz[60][311] = 9'b111111111;
assign micromatrizz[60][312] = 9'b111111111;
assign micromatrizz[60][313] = 9'b111111111;
assign micromatrizz[60][314] = 9'b111111111;
assign micromatrizz[60][315] = 9'b111110111;
assign micromatrizz[60][316] = 9'b111110010;
assign micromatrizz[60][317] = 9'b111110010;
assign micromatrizz[60][318] = 9'b111110011;
assign micromatrizz[60][319] = 9'b111110011;
assign micromatrizz[60][320] = 9'b111110011;
assign micromatrizz[60][321] = 9'b111110011;
assign micromatrizz[60][322] = 9'b111111111;
assign micromatrizz[60][323] = 9'b111111111;
assign micromatrizz[60][324] = 9'b111111111;
assign micromatrizz[60][325] = 9'b111111111;
assign micromatrizz[60][326] = 9'b111110010;
assign micromatrizz[60][327] = 9'b111110010;
assign micromatrizz[60][328] = 9'b111110011;
assign micromatrizz[60][329] = 9'b111110011;
assign micromatrizz[60][330] = 9'b111110011;
assign micromatrizz[60][331] = 9'b111110011;
assign micromatrizz[60][332] = 9'b111111111;
assign micromatrizz[60][333] = 9'b111111111;
assign micromatrizz[60][334] = 9'b111111111;
assign micromatrizz[60][335] = 9'b111110010;
assign micromatrizz[60][336] = 9'b111110011;
assign micromatrizz[60][337] = 9'b111110011;
assign micromatrizz[60][338] = 9'b111110011;
assign micromatrizz[60][339] = 9'b111110011;
assign micromatrizz[60][340] = 9'b111110011;
assign micromatrizz[60][341] = 9'b111110011;
assign micromatrizz[60][342] = 9'b111111111;
assign micromatrizz[60][343] = 9'b111111111;
assign micromatrizz[60][344] = 9'b111111111;
assign micromatrizz[60][345] = 9'b111111111;
assign micromatrizz[60][346] = 9'b111111111;
assign micromatrizz[60][347] = 9'b111110010;
assign micromatrizz[60][348] = 9'b111110010;
assign micromatrizz[60][349] = 9'b111110010;
assign micromatrizz[60][350] = 9'b111110010;
assign micromatrizz[60][351] = 9'b111110011;
assign micromatrizz[60][352] = 9'b111110011;
assign micromatrizz[60][353] = 9'b111110011;
assign micromatrizz[60][354] = 9'b111111111;
assign micromatrizz[60][355] = 9'b111111111;
assign micromatrizz[60][356] = 9'b111111111;
assign micromatrizz[60][357] = 9'b111111111;
assign micromatrizz[60][358] = 9'b111111111;
assign micromatrizz[60][359] = 9'b111110010;
assign micromatrizz[60][360] = 9'b111110011;
assign micromatrizz[60][361] = 9'b111110010;
assign micromatrizz[60][362] = 9'b111110010;
assign micromatrizz[60][363] = 9'b111110011;
assign micromatrizz[60][364] = 9'b111110011;
assign micromatrizz[60][365] = 9'b111110011;
assign micromatrizz[60][366] = 9'b111111111;
assign micromatrizz[60][367] = 9'b111111111;
assign micromatrizz[60][368] = 9'b111111111;
assign micromatrizz[60][369] = 9'b111111111;
assign micromatrizz[60][370] = 9'b111111111;
assign micromatrizz[60][371] = 9'b111111111;
assign micromatrizz[60][372] = 9'b111110010;
assign micromatrizz[60][373] = 9'b111110010;
assign micromatrizz[60][374] = 9'b111110011;
assign micromatrizz[60][375] = 9'b111110011;
assign micromatrizz[60][376] = 9'b111110011;
assign micromatrizz[60][377] = 9'b111110011;
assign micromatrizz[60][378] = 9'b111110011;
assign micromatrizz[60][379] = 9'b111111111;
assign micromatrizz[60][380] = 9'b111111111;
assign micromatrizz[60][381] = 9'b111111111;
assign micromatrizz[60][382] = 9'b111111111;
assign micromatrizz[60][383] = 9'b111110111;
assign micromatrizz[60][384] = 9'b111110010;
assign micromatrizz[60][385] = 9'b111110010;
assign micromatrizz[60][386] = 9'b111110011;
assign micromatrizz[60][387] = 9'b111110011;
assign micromatrizz[60][388] = 9'b111110011;
assign micromatrizz[60][389] = 9'b111110011;
assign micromatrizz[60][390] = 9'b111110011;
assign micromatrizz[60][391] = 9'b111111111;
assign micromatrizz[60][392] = 9'b111111111;
assign micromatrizz[60][393] = 9'b111111111;
assign micromatrizz[60][394] = 9'b111111111;
assign micromatrizz[60][395] = 9'b111110110;
assign micromatrizz[60][396] = 9'b111110010;
assign micromatrizz[60][397] = 9'b111110010;
assign micromatrizz[60][398] = 9'b111110010;
assign micromatrizz[60][399] = 9'b111110010;
assign micromatrizz[60][400] = 9'b111110011;
assign micromatrizz[60][401] = 9'b111110010;
assign micromatrizz[60][402] = 9'b111110111;
assign micromatrizz[60][403] = 9'b111111111;
assign micromatrizz[60][404] = 9'b111111111;
assign micromatrizz[60][405] = 9'b111111111;
assign micromatrizz[60][406] = 9'b111111111;
assign micromatrizz[60][407] = 9'b111111111;
assign micromatrizz[60][408] = 9'b111111111;
assign micromatrizz[60][409] = 9'b111111111;
assign micromatrizz[60][410] = 9'b111111111;
assign micromatrizz[60][411] = 9'b111110010;
assign micromatrizz[60][412] = 9'b111110010;
assign micromatrizz[60][413] = 9'b111110011;
assign micromatrizz[60][414] = 9'b111110011;
assign micromatrizz[60][415] = 9'b111110011;
assign micromatrizz[60][416] = 9'b111110011;
assign micromatrizz[60][417] = 9'b111110111;
assign micromatrizz[60][418] = 9'b111111111;
assign micromatrizz[60][419] = 9'b111111111;
assign micromatrizz[60][420] = 9'b111111111;
assign micromatrizz[60][421] = 9'b111110111;
assign micromatrizz[60][422] = 9'b111110010;
assign micromatrizz[60][423] = 9'b111110010;
assign micromatrizz[60][424] = 9'b111110011;
assign micromatrizz[60][425] = 9'b111110011;
assign micromatrizz[60][426] = 9'b111110010;
assign micromatrizz[60][427] = 9'b111110111;
assign micromatrizz[60][428] = 9'b111111111;
assign micromatrizz[60][429] = 9'b111111111;
assign micromatrizz[60][430] = 9'b111110111;
assign micromatrizz[60][431] = 9'b111110010;
assign micromatrizz[60][432] = 9'b111110010;
assign micromatrizz[60][433] = 9'b111110010;
assign micromatrizz[60][434] = 9'b111110010;
assign micromatrizz[60][435] = 9'b111110011;
assign micromatrizz[60][436] = 9'b111110011;
assign micromatrizz[60][437] = 9'b111110011;
assign micromatrizz[60][438] = 9'b111111111;
assign micromatrizz[60][439] = 9'b111111111;
assign micromatrizz[60][440] = 9'b111111111;
assign micromatrizz[60][441] = 9'b111111111;
assign micromatrizz[60][442] = 9'b111111111;
assign micromatrizz[60][443] = 9'b111111111;
assign micromatrizz[60][444] = 9'b111111111;
assign micromatrizz[60][445] = 9'b111111111;
assign micromatrizz[60][446] = 9'b111110010;
assign micromatrizz[60][447] = 9'b111110010;
assign micromatrizz[60][448] = 9'b111110010;
assign micromatrizz[60][449] = 9'b111110010;
assign micromatrizz[60][450] = 9'b111110010;
assign micromatrizz[60][451] = 9'b111110011;
assign micromatrizz[60][452] = 9'b111110011;
assign micromatrizz[60][453] = 9'b111110011;
assign micromatrizz[60][454] = 9'b111111111;
assign micromatrizz[60][455] = 9'b111111111;
assign micromatrizz[60][456] = 9'b111111111;
assign micromatrizz[60][457] = 9'b111111111;
assign micromatrizz[60][458] = 9'b111111111;
assign micromatrizz[60][459] = 9'b111111111;
assign micromatrizz[60][460] = 9'b111111111;
assign micromatrizz[60][461] = 9'b111111111;
assign micromatrizz[60][462] = 9'b111110111;
assign micromatrizz[60][463] = 9'b111111111;
assign micromatrizz[60][464] = 9'b111111111;
assign micromatrizz[60][465] = 9'b111111111;
assign micromatrizz[60][466] = 9'b111110010;
assign micromatrizz[60][467] = 9'b111110010;
assign micromatrizz[60][468] = 9'b111110010;
assign micromatrizz[60][469] = 9'b111110010;
assign micromatrizz[60][470] = 9'b111110010;
assign micromatrizz[60][471] = 9'b111110010;
assign micromatrizz[60][472] = 9'b111110010;
assign micromatrizz[60][473] = 9'b111110011;
assign micromatrizz[60][474] = 9'b111110011;
assign micromatrizz[60][475] = 9'b111110011;
assign micromatrizz[60][476] = 9'b111111111;
assign micromatrizz[60][477] = 9'b111111111;
assign micromatrizz[60][478] = 9'b111111111;
assign micromatrizz[60][479] = 9'b111111111;
assign micromatrizz[60][480] = 9'b111111111;
assign micromatrizz[60][481] = 9'b111110010;
assign micromatrizz[60][482] = 9'b111110010;
assign micromatrizz[60][483] = 9'b111110010;
assign micromatrizz[60][484] = 9'b111110010;
assign micromatrizz[60][485] = 9'b111110011;
assign micromatrizz[60][486] = 9'b111110011;
assign micromatrizz[60][487] = 9'b111110011;
assign micromatrizz[60][488] = 9'b111110111;
assign micromatrizz[60][489] = 9'b111111111;
assign micromatrizz[60][490] = 9'b111111111;
assign micromatrizz[60][491] = 9'b111111111;
assign micromatrizz[60][492] = 9'b111111111;
assign micromatrizz[60][493] = 9'b111111111;
assign micromatrizz[60][494] = 9'b111111111;
assign micromatrizz[60][495] = 9'b111111111;
assign micromatrizz[60][496] = 9'b111111111;
assign micromatrizz[60][497] = 9'b111110010;
assign micromatrizz[60][498] = 9'b111110011;
assign micromatrizz[60][499] = 9'b111110011;
assign micromatrizz[60][500] = 9'b111110011;
assign micromatrizz[60][501] = 9'b111110010;
assign micromatrizz[60][502] = 9'b111110010;
assign micromatrizz[60][503] = 9'b111110111;
assign micromatrizz[60][504] = 9'b111111111;
assign micromatrizz[60][505] = 9'b111111111;
assign micromatrizz[60][506] = 9'b111111111;
assign micromatrizz[60][507] = 9'b111110010;
assign micromatrizz[60][508] = 9'b111110010;
assign micromatrizz[60][509] = 9'b111110010;
assign micromatrizz[60][510] = 9'b111110010;
assign micromatrizz[60][511] = 9'b111110010;
assign micromatrizz[60][512] = 9'b111110010;
assign micromatrizz[60][513] = 9'b111111111;
assign micromatrizz[60][514] = 9'b111111111;
assign micromatrizz[60][515] = 9'b111111111;
assign micromatrizz[60][516] = 9'b111110111;
assign micromatrizz[60][517] = 9'b111110011;
assign micromatrizz[60][518] = 9'b111110011;
assign micromatrizz[60][519] = 9'b111110011;
assign micromatrizz[60][520] = 9'b111110010;
assign micromatrizz[60][521] = 9'b111110010;
assign micromatrizz[60][522] = 9'b111110011;
assign micromatrizz[60][523] = 9'b111110111;
assign micromatrizz[60][524] = 9'b111111111;
assign micromatrizz[60][525] = 9'b111111111;
assign micromatrizz[60][526] = 9'b111111111;
assign micromatrizz[60][527] = 9'b111111111;
assign micromatrizz[60][528] = 9'b111110111;
assign micromatrizz[60][529] = 9'b111110010;
assign micromatrizz[60][530] = 9'b111110010;
assign micromatrizz[60][531] = 9'b111110010;
assign micromatrizz[60][532] = 9'b111110011;
assign micromatrizz[60][533] = 9'b111110011;
assign micromatrizz[60][534] = 9'b111110011;
assign micromatrizz[60][535] = 9'b111110011;
assign micromatrizz[60][536] = 9'b111111111;
assign micromatrizz[60][537] = 9'b111111111;
assign micromatrizz[60][538] = 9'b111110111;
assign micromatrizz[60][539] = 9'b111110010;
assign micromatrizz[60][540] = 9'b111110011;
assign micromatrizz[60][541] = 9'b111110011;
assign micromatrizz[60][542] = 9'b111110010;
assign micromatrizz[60][543] = 9'b111110011;
assign micromatrizz[60][544] = 9'b111110011;
assign micromatrizz[60][545] = 9'b111111111;
assign micromatrizz[60][546] = 9'b111111111;
assign micromatrizz[60][547] = 9'b111111111;
assign micromatrizz[60][548] = 9'b111111111;
assign micromatrizz[60][549] = 9'b111110010;
assign micromatrizz[60][550] = 9'b111110010;
assign micromatrizz[60][551] = 9'b111110010;
assign micromatrizz[60][552] = 9'b111110011;
assign micromatrizz[60][553] = 9'b111110010;
assign micromatrizz[60][554] = 9'b111110010;
assign micromatrizz[60][555] = 9'b111111111;
assign micromatrizz[60][556] = 9'b111111111;
assign micromatrizz[60][557] = 9'b111111111;
assign micromatrizz[60][558] = 9'b111110010;
assign micromatrizz[60][559] = 9'b111110010;
assign micromatrizz[60][560] = 9'b111110010;
assign micromatrizz[60][561] = 9'b111110010;
assign micromatrizz[60][562] = 9'b111110011;
assign micromatrizz[60][563] = 9'b111110011;
assign micromatrizz[60][564] = 9'b111110010;
assign micromatrizz[60][565] = 9'b111111111;
assign micromatrizz[60][566] = 9'b111111111;
assign micromatrizz[60][567] = 9'b111111111;
assign micromatrizz[60][568] = 9'b111110010;
assign micromatrizz[60][569] = 9'b111110010;
assign micromatrizz[60][570] = 9'b111110010;
assign micromatrizz[60][571] = 9'b111110010;
assign micromatrizz[60][572] = 9'b111110010;
assign micromatrizz[60][573] = 9'b111110011;
assign micromatrizz[60][574] = 9'b111110011;
assign micromatrizz[60][575] = 9'b111110011;
assign micromatrizz[60][576] = 9'b111111111;
assign micromatrizz[60][577] = 9'b111111111;
assign micromatrizz[60][578] = 9'b111111111;
assign micromatrizz[60][579] = 9'b111111111;
assign micromatrizz[60][580] = 9'b111111111;
assign micromatrizz[60][581] = 9'b111110010;
assign micromatrizz[60][582] = 9'b111110011;
assign micromatrizz[60][583] = 9'b111110010;
assign micromatrizz[60][584] = 9'b111110011;
assign micromatrizz[60][585] = 9'b111110011;
assign micromatrizz[60][586] = 9'b111110011;
assign micromatrizz[60][587] = 9'b111110010;
assign micromatrizz[60][588] = 9'b111111111;
assign micromatrizz[60][589] = 9'b111111111;
assign micromatrizz[60][590] = 9'b111111111;
assign micromatrizz[60][591] = 9'b111110111;
assign micromatrizz[60][592] = 9'b111110010;
assign micromatrizz[60][593] = 9'b111110010;
assign micromatrizz[60][594] = 9'b111110011;
assign micromatrizz[60][595] = 9'b111110011;
assign micromatrizz[60][596] = 9'b111110011;
assign micromatrizz[60][597] = 9'b111110011;
assign micromatrizz[60][598] = 9'b111111111;
assign micromatrizz[60][599] = 9'b111111111;
assign micromatrizz[60][600] = 9'b111111111;
assign micromatrizz[60][601] = 9'b111111111;
assign micromatrizz[60][602] = 9'b111110010;
assign micromatrizz[60][603] = 9'b111110011;
assign micromatrizz[60][604] = 9'b111110011;
assign micromatrizz[60][605] = 9'b111110011;
assign micromatrizz[60][606] = 9'b111110011;
assign micromatrizz[60][607] = 9'b111110111;
assign micromatrizz[60][608] = 9'b111111111;
assign micromatrizz[60][609] = 9'b111111111;
assign micromatrizz[60][610] = 9'b111111111;
assign micromatrizz[60][611] = 9'b111110010;
assign micromatrizz[60][612] = 9'b111110010;
assign micromatrizz[60][613] = 9'b111110010;
assign micromatrizz[60][614] = 9'b111110010;
assign micromatrizz[60][615] = 9'b111110011;
assign micromatrizz[60][616] = 9'b111110011;
assign micromatrizz[60][617] = 9'b111110011;
assign micromatrizz[60][618] = 9'b111110011;
assign micromatrizz[60][619] = 9'b111110011;
assign micromatrizz[60][620] = 9'b111110111;
assign micromatrizz[60][621] = 9'b111111111;
assign micromatrizz[60][622] = 9'b111111111;
assign micromatrizz[60][623] = 9'b111111111;
assign micromatrizz[60][624] = 9'b111111111;
assign micromatrizz[60][625] = 9'b111111111;
assign micromatrizz[60][626] = 9'b111111111;
assign micromatrizz[60][627] = 9'b111111111;
assign micromatrizz[60][628] = 9'b111111111;
assign micromatrizz[60][629] = 9'b111111111;
assign micromatrizz[60][630] = 9'b111111111;
assign micromatrizz[60][631] = 9'b111111111;
assign micromatrizz[60][632] = 9'b111111111;
assign micromatrizz[60][633] = 9'b111111111;
assign micromatrizz[60][634] = 9'b111111111;
assign micromatrizz[60][635] = 9'b111111111;
assign micromatrizz[60][636] = 9'b111111111;
assign micromatrizz[60][637] = 9'b111111111;
assign micromatrizz[60][638] = 9'b111111111;
assign micromatrizz[60][639] = 9'b111111111;
assign micromatrizz[61][0] = 9'b111111111;
assign micromatrizz[61][1] = 9'b111111111;
assign micromatrizz[61][2] = 9'b111111111;
assign micromatrizz[61][3] = 9'b111111111;
assign micromatrizz[61][4] = 9'b111111111;
assign micromatrizz[61][5] = 9'b111111111;
assign micromatrizz[61][6] = 9'b111111111;
assign micromatrizz[61][7] = 9'b111111111;
assign micromatrizz[61][8] = 9'b111111111;
assign micromatrizz[61][9] = 9'b111110111;
assign micromatrizz[61][10] = 9'b111110010;
assign micromatrizz[61][11] = 9'b111110010;
assign micromatrizz[61][12] = 9'b111110010;
assign micromatrizz[61][13] = 9'b111110010;
assign micromatrizz[61][14] = 9'b111110011;
assign micromatrizz[61][15] = 9'b111110010;
assign micromatrizz[61][16] = 9'b111110011;
assign micromatrizz[61][17] = 9'b111110011;
assign micromatrizz[61][18] = 9'b111110011;
assign micromatrizz[61][19] = 9'b111110111;
assign micromatrizz[61][20] = 9'b111111111;
assign micromatrizz[61][21] = 9'b111111111;
assign micromatrizz[61][22] = 9'b111111111;
assign micromatrizz[61][23] = 9'b111110111;
assign micromatrizz[61][24] = 9'b111110010;
assign micromatrizz[61][25] = 9'b111110010;
assign micromatrizz[61][26] = 9'b111110010;
assign micromatrizz[61][27] = 9'b111110011;
assign micromatrizz[61][28] = 9'b111110011;
assign micromatrizz[61][29] = 9'b111110011;
assign micromatrizz[61][30] = 9'b111110011;
assign micromatrizz[61][31] = 9'b111111111;
assign micromatrizz[61][32] = 9'b111111111;
assign micromatrizz[61][33] = 9'b111111111;
assign micromatrizz[61][34] = 9'b111111111;
assign micromatrizz[61][35] = 9'b111110111;
assign micromatrizz[61][36] = 9'b111110010;
assign micromatrizz[61][37] = 9'b111110010;
assign micromatrizz[61][38] = 9'b111110011;
assign micromatrizz[61][39] = 9'b111110011;
assign micromatrizz[61][40] = 9'b111110011;
assign micromatrizz[61][41] = 9'b111110011;
assign micromatrizz[61][42] = 9'b111110011;
assign micromatrizz[61][43] = 9'b111111111;
assign micromatrizz[61][44] = 9'b111111111;
assign micromatrizz[61][45] = 9'b111111111;
assign micromatrizz[61][46] = 9'b111111111;
assign micromatrizz[61][47] = 9'b111110010;
assign micromatrizz[61][48] = 9'b111110010;
assign micromatrizz[61][49] = 9'b111110010;
assign micromatrizz[61][50] = 9'b111110011;
assign micromatrizz[61][51] = 9'b111110011;
assign micromatrizz[61][52] = 9'b111110011;
assign micromatrizz[61][53] = 9'b111110011;
assign micromatrizz[61][54] = 9'b111111111;
assign micromatrizz[61][55] = 9'b111111111;
assign micromatrizz[61][56] = 9'b111111111;
assign micromatrizz[61][57] = 9'b111111111;
assign micromatrizz[61][58] = 9'b111111111;
assign micromatrizz[61][59] = 9'b111110010;
assign micromatrizz[61][60] = 9'b111110010;
assign micromatrizz[61][61] = 9'b111110010;
assign micromatrizz[61][62] = 9'b111110011;
assign micromatrizz[61][63] = 9'b111110011;
assign micromatrizz[61][64] = 9'b111110011;
assign micromatrizz[61][65] = 9'b111110011;
assign micromatrizz[61][66] = 9'b111111111;
assign micromatrizz[61][67] = 9'b111111111;
assign micromatrizz[61][68] = 9'b111110111;
assign micromatrizz[61][69] = 9'b111110010;
assign micromatrizz[61][70] = 9'b111110010;
assign micromatrizz[61][71] = 9'b111110010;
assign micromatrizz[61][72] = 9'b111110010;
assign micromatrizz[61][73] = 9'b111110011;
assign micromatrizz[61][74] = 9'b111110011;
assign micromatrizz[61][75] = 9'b111110111;
assign micromatrizz[61][76] = 9'b111110111;
assign micromatrizz[61][77] = 9'b111111111;
assign micromatrizz[61][78] = 9'b111110111;
assign micromatrizz[61][79] = 9'b111110110;
assign micromatrizz[61][80] = 9'b111110111;
assign micromatrizz[61][81] = 9'b111110111;
assign micromatrizz[61][82] = 9'b111110111;
assign micromatrizz[61][83] = 9'b111110111;
assign micromatrizz[61][84] = 9'b111110111;
assign micromatrizz[61][85] = 9'b111111111;
assign micromatrizz[61][86] = 9'b111111111;
assign micromatrizz[61][87] = 9'b111111111;
assign micromatrizz[61][88] = 9'b111110010;
assign micromatrizz[61][89] = 9'b111110010;
assign micromatrizz[61][90] = 9'b111110010;
assign micromatrizz[61][91] = 9'b111110010;
assign micromatrizz[61][92] = 9'b111110011;
assign micromatrizz[61][93] = 9'b111110011;
assign micromatrizz[61][94] = 9'b111110011;
assign micromatrizz[61][95] = 9'b111110111;
assign micromatrizz[61][96] = 9'b111111111;
assign micromatrizz[61][97] = 9'b111111111;
assign micromatrizz[61][98] = 9'b111111111;
assign micromatrizz[61][99] = 9'b111111111;
assign micromatrizz[61][100] = 9'b111111111;
assign micromatrizz[61][101] = 9'b111111111;
assign micromatrizz[61][102] = 9'b111111111;
assign micromatrizz[61][103] = 9'b111111111;
assign micromatrizz[61][104] = 9'b111111111;
assign micromatrizz[61][105] = 9'b111110111;
assign micromatrizz[61][106] = 9'b111110010;
assign micromatrizz[61][107] = 9'b111110010;
assign micromatrizz[61][108] = 9'b111110010;
assign micromatrizz[61][109] = 9'b111110010;
assign micromatrizz[61][110] = 9'b111110011;
assign micromatrizz[61][111] = 9'b111110011;
assign micromatrizz[61][112] = 9'b111110011;
assign micromatrizz[61][113] = 9'b111110011;
assign micromatrizz[61][114] = 9'b111110011;
assign micromatrizz[61][115] = 9'b111110111;
assign micromatrizz[61][116] = 9'b111111111;
assign micromatrizz[61][117] = 9'b111111111;
assign micromatrizz[61][118] = 9'b111111111;
assign micromatrizz[61][119] = 9'b111110010;
assign micromatrizz[61][120] = 9'b111110010;
assign micromatrizz[61][121] = 9'b111110010;
assign micromatrizz[61][122] = 9'b111110010;
assign micromatrizz[61][123] = 9'b111110010;
assign micromatrizz[61][124] = 9'b111110011;
assign micromatrizz[61][125] = 9'b111110011;
assign micromatrizz[61][126] = 9'b111110111;
assign micromatrizz[61][127] = 9'b111111111;
assign micromatrizz[61][128] = 9'b111111111;
assign micromatrizz[61][129] = 9'b111111111;
assign micromatrizz[61][130] = 9'b111111111;
assign micromatrizz[61][131] = 9'b111111111;
assign micromatrizz[61][132] = 9'b111111111;
assign micromatrizz[61][133] = 9'b111111111;
assign micromatrizz[61][134] = 9'b111110111;
assign micromatrizz[61][135] = 9'b111110111;
assign micromatrizz[61][136] = 9'b111111111;
assign micromatrizz[61][137] = 9'b111111111;
assign micromatrizz[61][138] = 9'b111110111;
assign micromatrizz[61][139] = 9'b111110010;
assign micromatrizz[61][140] = 9'b111110010;
assign micromatrizz[61][141] = 9'b111110010;
assign micromatrizz[61][142] = 9'b111110010;
assign micromatrizz[61][143] = 9'b111110011;
assign micromatrizz[61][144] = 9'b111110011;
assign micromatrizz[61][145] = 9'b111110011;
assign micromatrizz[61][146] = 9'b111111111;
assign micromatrizz[61][147] = 9'b111111111;
assign micromatrizz[61][148] = 9'b111111111;
assign micromatrizz[61][149] = 9'b111111111;
assign micromatrizz[61][150] = 9'b111110111;
assign micromatrizz[61][151] = 9'b111110010;
assign micromatrizz[61][152] = 9'b111110010;
assign micromatrizz[61][153] = 9'b111110010;
assign micromatrizz[61][154] = 9'b111110011;
assign micromatrizz[61][155] = 9'b111110011;
assign micromatrizz[61][156] = 9'b111110011;
assign micromatrizz[61][157] = 9'b111110011;
assign micromatrizz[61][158] = 9'b111111111;
assign micromatrizz[61][159] = 9'b111111111;
assign micromatrizz[61][160] = 9'b111111111;
assign micromatrizz[61][161] = 9'b111110111;
assign micromatrizz[61][162] = 9'b111110010;
assign micromatrizz[61][163] = 9'b111110010;
assign micromatrizz[61][164] = 9'b111110011;
assign micromatrizz[61][165] = 9'b111110011;
assign micromatrizz[61][166] = 9'b111110011;
assign micromatrizz[61][167] = 9'b111110011;
assign micromatrizz[61][168] = 9'b111111111;
assign micromatrizz[61][169] = 9'b111111111;
assign micromatrizz[61][170] = 9'b111111111;
assign micromatrizz[61][171] = 9'b111111111;
assign micromatrizz[61][172] = 9'b111110011;
assign micromatrizz[61][173] = 9'b111110010;
assign micromatrizz[61][174] = 9'b111110011;
assign micromatrizz[61][175] = 9'b111110011;
assign micromatrizz[61][176] = 9'b111110011;
assign micromatrizz[61][177] = 9'b111110011;
assign micromatrizz[61][178] = 9'b111110010;
assign micromatrizz[61][179] = 9'b111110111;
assign micromatrizz[61][180] = 9'b111111111;
assign micromatrizz[61][181] = 9'b111111111;
assign micromatrizz[61][182] = 9'b111110110;
assign micromatrizz[61][183] = 9'b111110010;
assign micromatrizz[61][184] = 9'b111110010;
assign micromatrizz[61][185] = 9'b111110011;
assign micromatrizz[61][186] = 9'b111110010;
assign micromatrizz[61][187] = 9'b111110010;
assign micromatrizz[61][188] = 9'b111110011;
assign micromatrizz[61][189] = 9'b111110011;
assign micromatrizz[61][190] = 9'b111110111;
assign micromatrizz[61][191] = 9'b111111111;
assign micromatrizz[61][192] = 9'b111111111;
assign micromatrizz[61][193] = 9'b111111111;
assign micromatrizz[61][194] = 9'b111111111;
assign micromatrizz[61][195] = 9'b111110010;
assign micromatrizz[61][196] = 9'b111110010;
assign micromatrizz[61][197] = 9'b111110011;
assign micromatrizz[61][198] = 9'b111110011;
assign micromatrizz[61][199] = 9'b111110010;
assign micromatrizz[61][200] = 9'b111110010;
assign micromatrizz[61][201] = 9'b111110011;
assign micromatrizz[61][202] = 9'b111110111;
assign micromatrizz[61][203] = 9'b111111111;
assign micromatrizz[61][204] = 9'b111111111;
assign micromatrizz[61][205] = 9'b111110111;
assign micromatrizz[61][206] = 9'b111110010;
assign micromatrizz[61][207] = 9'b111110010;
assign micromatrizz[61][208] = 9'b111110010;
assign micromatrizz[61][209] = 9'b111110010;
assign micromatrizz[61][210] = 9'b111110011;
assign micromatrizz[61][211] = 9'b111110011;
assign micromatrizz[61][212] = 9'b111110011;
assign micromatrizz[61][213] = 9'b111110111;
assign micromatrizz[61][214] = 9'b111111111;
assign micromatrizz[61][215] = 9'b111111111;
assign micromatrizz[61][216] = 9'b111111111;
assign micromatrizz[61][217] = 9'b111111111;
assign micromatrizz[61][218] = 9'b111111111;
assign micromatrizz[61][219] = 9'b111111111;
assign micromatrizz[61][220] = 9'b111111111;
assign micromatrizz[61][221] = 9'b111110111;
assign micromatrizz[61][222] = 9'b111111111;
assign micromatrizz[61][223] = 9'b111111111;
assign micromatrizz[61][224] = 9'b111111111;
assign micromatrizz[61][225] = 9'b111110010;
assign micromatrizz[61][226] = 9'b111110010;
assign micromatrizz[61][227] = 9'b111110010;
assign micromatrizz[61][228] = 9'b111110010;
assign micromatrizz[61][229] = 9'b111110011;
assign micromatrizz[61][230] = 9'b111110011;
assign micromatrizz[61][231] = 9'b111110011;
assign micromatrizz[61][232] = 9'b111110111;
assign micromatrizz[61][233] = 9'b111111111;
assign micromatrizz[61][234] = 9'b111111111;
assign micromatrizz[61][235] = 9'b111111111;
assign micromatrizz[61][236] = 9'b111111111;
assign micromatrizz[61][237] = 9'b111111111;
assign micromatrizz[61][238] = 9'b111111111;
assign micromatrizz[61][239] = 9'b111111111;
assign micromatrizz[61][240] = 9'b111111111;
assign micromatrizz[61][241] = 9'b111110010;
assign micromatrizz[61][242] = 9'b111110010;
assign micromatrizz[61][243] = 9'b111110010;
assign micromatrizz[61][244] = 9'b111110011;
assign micromatrizz[61][245] = 9'b111110011;
assign micromatrizz[61][246] = 9'b111110011;
assign micromatrizz[61][247] = 9'b111110011;
assign micromatrizz[61][248] = 9'b111110111;
assign micromatrizz[61][249] = 9'b111110111;
assign micromatrizz[61][250] = 9'b111110111;
assign micromatrizz[61][251] = 9'b111110111;
assign micromatrizz[61][252] = 9'b111110110;
assign micromatrizz[61][253] = 9'b111110110;
assign micromatrizz[61][254] = 9'b111110111;
assign micromatrizz[61][255] = 9'b111110011;
assign micromatrizz[61][256] = 9'b111110111;
assign micromatrizz[61][257] = 9'b111111111;
assign micromatrizz[61][258] = 9'b111111111;
assign micromatrizz[61][259] = 9'b111111111;
assign micromatrizz[61][260] = 9'b111111111;
assign micromatrizz[61][261] = 9'b111110110;
assign micromatrizz[61][262] = 9'b111110010;
assign micromatrizz[61][263] = 9'b111110010;
assign micromatrizz[61][264] = 9'b111110010;
assign micromatrizz[61][265] = 9'b111110010;
assign micromatrizz[61][266] = 9'b111110010;
assign micromatrizz[61][267] = 9'b111110011;
assign micromatrizz[61][268] = 9'b111110011;
assign micromatrizz[61][269] = 9'b111110011;
assign micromatrizz[61][270] = 9'b111110011;
assign micromatrizz[61][271] = 9'b111110111;
assign micromatrizz[61][272] = 9'b111111111;
assign micromatrizz[61][273] = 9'b111111111;
assign micromatrizz[61][274] = 9'b111111111;
assign micromatrizz[61][275] = 9'b111110111;
assign micromatrizz[61][276] = 9'b111110010;
assign micromatrizz[61][277] = 9'b111110010;
assign micromatrizz[61][278] = 9'b111110010;
assign micromatrizz[61][279] = 9'b111110011;
assign micromatrizz[61][280] = 9'b111110011;
assign micromatrizz[61][281] = 9'b111110011;
assign micromatrizz[61][282] = 9'b111111111;
assign micromatrizz[61][283] = 9'b111111111;
assign micromatrizz[61][284] = 9'b111111111;
assign micromatrizz[61][285] = 9'b111111111;
assign micromatrizz[61][286] = 9'b111110011;
assign micromatrizz[61][287] = 9'b111110010;
assign micromatrizz[61][288] = 9'b111110010;
assign micromatrizz[61][289] = 9'b111110011;
assign micromatrizz[61][290] = 9'b111110011;
assign micromatrizz[61][291] = 9'b111110011;
assign micromatrizz[61][292] = 9'b111110011;
assign micromatrizz[61][293] = 9'b111111111;
assign micromatrizz[61][294] = 9'b111111111;
assign micromatrizz[61][295] = 9'b111111111;
assign micromatrizz[61][296] = 9'b111111111;
assign micromatrizz[61][297] = 9'b111111111;
assign micromatrizz[61][298] = 9'b111111111;
assign micromatrizz[61][299] = 9'b111111111;
assign micromatrizz[61][300] = 9'b111110111;
assign micromatrizz[61][301] = 9'b111110010;
assign micromatrizz[61][302] = 9'b111110010;
assign micromatrizz[61][303] = 9'b111110010;
assign micromatrizz[61][304] = 9'b111110010;
assign micromatrizz[61][305] = 9'b111110010;
assign micromatrizz[61][306] = 9'b111110010;
assign micromatrizz[61][307] = 9'b111110011;
assign micromatrizz[61][308] = 9'b111110011;
assign micromatrizz[61][309] = 9'b111110011;
assign micromatrizz[61][310] = 9'b111111111;
assign micromatrizz[61][311] = 9'b111111111;
assign micromatrizz[61][312] = 9'b111111111;
assign micromatrizz[61][313] = 9'b111111111;
assign micromatrizz[61][314] = 9'b111111111;
assign micromatrizz[61][315] = 9'b111110111;
assign micromatrizz[61][316] = 9'b111110010;
assign micromatrizz[61][317] = 9'b111110011;
assign micromatrizz[61][318] = 9'b111110010;
assign micromatrizz[61][319] = 9'b111110011;
assign micromatrizz[61][320] = 9'b111110011;
assign micromatrizz[61][321] = 9'b111110011;
assign micromatrizz[61][322] = 9'b111110111;
assign micromatrizz[61][323] = 9'b111110111;
assign micromatrizz[61][324] = 9'b111110111;
assign micromatrizz[61][325] = 9'b111110111;
assign micromatrizz[61][326] = 9'b111110110;
assign micromatrizz[61][327] = 9'b111110111;
assign micromatrizz[61][328] = 9'b111110111;
assign micromatrizz[61][329] = 9'b111110111;
assign micromatrizz[61][330] = 9'b111110111;
assign micromatrizz[61][331] = 9'b111110111;
assign micromatrizz[61][332] = 9'b111111111;
assign micromatrizz[61][333] = 9'b111111111;
assign micromatrizz[61][334] = 9'b111111111;
assign micromatrizz[61][335] = 9'b111110010;
assign micromatrizz[61][336] = 9'b111110011;
assign micromatrizz[61][337] = 9'b111110011;
assign micromatrizz[61][338] = 9'b111110011;
assign micromatrizz[61][339] = 9'b111110010;
assign micromatrizz[61][340] = 9'b111110011;
assign micromatrizz[61][341] = 9'b111110011;
assign micromatrizz[61][342] = 9'b111111111;
assign micromatrizz[61][343] = 9'b111111111;
assign micromatrizz[61][344] = 9'b111111111;
assign micromatrizz[61][345] = 9'b111111111;
assign micromatrizz[61][346] = 9'b111111111;
assign micromatrizz[61][347] = 9'b111110010;
assign micromatrizz[61][348] = 9'b111110010;
assign micromatrizz[61][349] = 9'b111110010;
assign micromatrizz[61][350] = 9'b111110010;
assign micromatrizz[61][351] = 9'b111110011;
assign micromatrizz[61][352] = 9'b111110011;
assign micromatrizz[61][353] = 9'b111110011;
assign micromatrizz[61][354] = 9'b111111111;
assign micromatrizz[61][355] = 9'b111111111;
assign micromatrizz[61][356] = 9'b111111111;
assign micromatrizz[61][357] = 9'b111111111;
assign micromatrizz[61][358] = 9'b111111111;
assign micromatrizz[61][359] = 9'b111110010;
assign micromatrizz[61][360] = 9'b111110011;
assign micromatrizz[61][361] = 9'b111110010;
assign micromatrizz[61][362] = 9'b111110010;
assign micromatrizz[61][363] = 9'b111110011;
assign micromatrizz[61][364] = 9'b111110011;
assign micromatrizz[61][365] = 9'b111110011;
assign micromatrizz[61][366] = 9'b111111111;
assign micromatrizz[61][367] = 9'b111111111;
assign micromatrizz[61][368] = 9'b111111111;
assign micromatrizz[61][369] = 9'b111111111;
assign micromatrizz[61][370] = 9'b111111111;
assign micromatrizz[61][371] = 9'b111111111;
assign micromatrizz[61][372] = 9'b111110010;
assign micromatrizz[61][373] = 9'b111110010;
assign micromatrizz[61][374] = 9'b111110011;
assign micromatrizz[61][375] = 9'b111110011;
assign micromatrizz[61][376] = 9'b111110011;
assign micromatrizz[61][377] = 9'b111110011;
assign micromatrizz[61][378] = 9'b111110011;
assign micromatrizz[61][379] = 9'b111111111;
assign micromatrizz[61][380] = 9'b111111111;
assign micromatrizz[61][381] = 9'b111111111;
assign micromatrizz[61][382] = 9'b111111111;
assign micromatrizz[61][383] = 9'b111110111;
assign micromatrizz[61][384] = 9'b111110010;
assign micromatrizz[61][385] = 9'b111110010;
assign micromatrizz[61][386] = 9'b111110011;
assign micromatrizz[61][387] = 9'b111110011;
assign micromatrizz[61][388] = 9'b111110011;
assign micromatrizz[61][389] = 9'b111110011;
assign micromatrizz[61][390] = 9'b111110011;
assign micromatrizz[61][391] = 9'b111111111;
assign micromatrizz[61][392] = 9'b111111111;
assign micromatrizz[61][393] = 9'b111111111;
assign micromatrizz[61][394] = 9'b111111111;
assign micromatrizz[61][395] = 9'b111110110;
assign micromatrizz[61][396] = 9'b111110010;
assign micromatrizz[61][397] = 9'b111110010;
assign micromatrizz[61][398] = 9'b111110010;
assign micromatrizz[61][399] = 9'b111110010;
assign micromatrizz[61][400] = 9'b111110011;
assign micromatrizz[61][401] = 9'b111110011;
assign micromatrizz[61][402] = 9'b111110111;
assign micromatrizz[61][403] = 9'b111111111;
assign micromatrizz[61][404] = 9'b111111111;
assign micromatrizz[61][405] = 9'b111111111;
assign micromatrizz[61][406] = 9'b111111111;
assign micromatrizz[61][407] = 9'b111111111;
assign micromatrizz[61][408] = 9'b111111111;
assign micromatrizz[61][409] = 9'b111111111;
assign micromatrizz[61][410] = 9'b111111111;
assign micromatrizz[61][411] = 9'b111110010;
assign micromatrizz[61][412] = 9'b111110010;
assign micromatrizz[61][413] = 9'b111110010;
assign micromatrizz[61][414] = 9'b111110011;
assign micromatrizz[61][415] = 9'b111110011;
assign micromatrizz[61][416] = 9'b111110011;
assign micromatrizz[61][417] = 9'b111110011;
assign micromatrizz[61][418] = 9'b111110111;
assign micromatrizz[61][419] = 9'b111110111;
assign micromatrizz[61][420] = 9'b111110111;
assign micromatrizz[61][421] = 9'b111110111;
assign micromatrizz[61][422] = 9'b111110111;
assign micromatrizz[61][423] = 9'b111110110;
assign micromatrizz[61][424] = 9'b111110111;
assign micromatrizz[61][425] = 9'b111110111;
assign micromatrizz[61][426] = 9'b111110111;
assign micromatrizz[61][427] = 9'b111111111;
assign micromatrizz[61][428] = 9'b111111111;
assign micromatrizz[61][429] = 9'b111111111;
assign micromatrizz[61][430] = 9'b111110111;
assign micromatrizz[61][431] = 9'b111110010;
assign micromatrizz[61][432] = 9'b111110010;
assign micromatrizz[61][433] = 9'b111110010;
assign micromatrizz[61][434] = 9'b111110010;
assign micromatrizz[61][435] = 9'b111110011;
assign micromatrizz[61][436] = 9'b111110011;
assign micromatrizz[61][437] = 9'b111110011;
assign micromatrizz[61][438] = 9'b111111111;
assign micromatrizz[61][439] = 9'b111111111;
assign micromatrizz[61][440] = 9'b111111111;
assign micromatrizz[61][441] = 9'b111111111;
assign micromatrizz[61][442] = 9'b111111111;
assign micromatrizz[61][443] = 9'b111111111;
assign micromatrizz[61][444] = 9'b111111111;
assign micromatrizz[61][445] = 9'b111111111;
assign micromatrizz[61][446] = 9'b111110010;
assign micromatrizz[61][447] = 9'b111110011;
assign micromatrizz[61][448] = 9'b111110010;
assign micromatrizz[61][449] = 9'b111110010;
assign micromatrizz[61][450] = 9'b111110010;
assign micromatrizz[61][451] = 9'b111110011;
assign micromatrizz[61][452] = 9'b111110011;
assign micromatrizz[61][453] = 9'b111110011;
assign micromatrizz[61][454] = 9'b111111111;
assign micromatrizz[61][455] = 9'b111111111;
assign micromatrizz[61][456] = 9'b111111111;
assign micromatrizz[61][457] = 9'b111111111;
assign micromatrizz[61][458] = 9'b111111111;
assign micromatrizz[61][459] = 9'b111111111;
assign micromatrizz[61][460] = 9'b111111111;
assign micromatrizz[61][461] = 9'b111111111;
assign micromatrizz[61][462] = 9'b111110111;
assign micromatrizz[61][463] = 9'b111111111;
assign micromatrizz[61][464] = 9'b111111111;
assign micromatrizz[61][465] = 9'b111111111;
assign micromatrizz[61][466] = 9'b111110111;
assign micromatrizz[61][467] = 9'b111110010;
assign micromatrizz[61][468] = 9'b111110010;
assign micromatrizz[61][469] = 9'b111110010;
assign micromatrizz[61][470] = 9'b111110010;
assign micromatrizz[61][471] = 9'b111110010;
assign micromatrizz[61][472] = 9'b111110011;
assign micromatrizz[61][473] = 9'b111110011;
assign micromatrizz[61][474] = 9'b111110011;
assign micromatrizz[61][475] = 9'b111110011;
assign micromatrizz[61][476] = 9'b111110111;
assign micromatrizz[61][477] = 9'b111111111;
assign micromatrizz[61][478] = 9'b111111111;
assign micromatrizz[61][479] = 9'b111111111;
assign micromatrizz[61][480] = 9'b111111111;
assign micromatrizz[61][481] = 9'b111110010;
assign micromatrizz[61][482] = 9'b111110010;
assign micromatrizz[61][483] = 9'b111110010;
assign micromatrizz[61][484] = 9'b111110010;
assign micromatrizz[61][485] = 9'b111110011;
assign micromatrizz[61][486] = 9'b111110011;
assign micromatrizz[61][487] = 9'b111110011;
assign micromatrizz[61][488] = 9'b111110111;
assign micromatrizz[61][489] = 9'b111111111;
assign micromatrizz[61][490] = 9'b111111111;
assign micromatrizz[61][491] = 9'b111111111;
assign micromatrizz[61][492] = 9'b111111111;
assign micromatrizz[61][493] = 9'b111111111;
assign micromatrizz[61][494] = 9'b111111111;
assign micromatrizz[61][495] = 9'b111111111;
assign micromatrizz[61][496] = 9'b111111111;
assign micromatrizz[61][497] = 9'b111110010;
assign micromatrizz[61][498] = 9'b111110010;
assign micromatrizz[61][499] = 9'b111110011;
assign micromatrizz[61][500] = 9'b111110011;
assign micromatrizz[61][501] = 9'b111110011;
assign micromatrizz[61][502] = 9'b111110011;
assign micromatrizz[61][503] = 9'b111110011;
assign micromatrizz[61][504] = 9'b111110111;
assign micromatrizz[61][505] = 9'b111110111;
assign micromatrizz[61][506] = 9'b111110111;
assign micromatrizz[61][507] = 9'b111110111;
assign micromatrizz[61][508] = 9'b111110110;
assign micromatrizz[61][509] = 9'b111110110;
assign micromatrizz[61][510] = 9'b111110111;
assign micromatrizz[61][511] = 9'b111110111;
assign micromatrizz[61][512] = 9'b111110111;
assign micromatrizz[61][513] = 9'b111111111;
assign micromatrizz[61][514] = 9'b111111111;
assign micromatrizz[61][515] = 9'b111111111;
assign micromatrizz[61][516] = 9'b111110111;
assign micromatrizz[61][517] = 9'b111110010;
assign micromatrizz[61][518] = 9'b111110011;
assign micromatrizz[61][519] = 9'b111110011;
assign micromatrizz[61][520] = 9'b111110010;
assign micromatrizz[61][521] = 9'b111110010;
assign micromatrizz[61][522] = 9'b111110011;
assign micromatrizz[61][523] = 9'b111110111;
assign micromatrizz[61][524] = 9'b111111111;
assign micromatrizz[61][525] = 9'b111111111;
assign micromatrizz[61][526] = 9'b111111111;
assign micromatrizz[61][527] = 9'b111111111;
assign micromatrizz[61][528] = 9'b111110111;
assign micromatrizz[61][529] = 9'b111110010;
assign micromatrizz[61][530] = 9'b111110010;
assign micromatrizz[61][531] = 9'b111110010;
assign micromatrizz[61][532] = 9'b111110011;
assign micromatrizz[61][533] = 9'b111110011;
assign micromatrizz[61][534] = 9'b111110011;
assign micromatrizz[61][535] = 9'b111110011;
assign micromatrizz[61][536] = 9'b111110111;
assign micromatrizz[61][537] = 9'b111111111;
assign micromatrizz[61][538] = 9'b111110111;
assign micromatrizz[61][539] = 9'b111110010;
assign micromatrizz[61][540] = 9'b111110010;
assign micromatrizz[61][541] = 9'b111110011;
assign micromatrizz[61][542] = 9'b111110011;
assign micromatrizz[61][543] = 9'b111110010;
assign micromatrizz[61][544] = 9'b111110011;
assign micromatrizz[61][545] = 9'b111110111;
assign micromatrizz[61][546] = 9'b111110111;
assign micromatrizz[61][547] = 9'b111111111;
assign micromatrizz[61][548] = 9'b111110111;
assign micromatrizz[61][549] = 9'b111110111;
assign micromatrizz[61][550] = 9'b111110111;
assign micromatrizz[61][551] = 9'b111110111;
assign micromatrizz[61][552] = 9'b111110111;
assign micromatrizz[61][553] = 9'b111110111;
assign micromatrizz[61][554] = 9'b111110111;
assign micromatrizz[61][555] = 9'b111111111;
assign micromatrizz[61][556] = 9'b111111111;
assign micromatrizz[61][557] = 9'b111111111;
assign micromatrizz[61][558] = 9'b111110010;
assign micromatrizz[61][559] = 9'b111110010;
assign micromatrizz[61][560] = 9'b111110010;
assign micromatrizz[61][561] = 9'b111110010;
assign micromatrizz[61][562] = 9'b111110011;
assign micromatrizz[61][563] = 9'b111110011;
assign micromatrizz[61][564] = 9'b111110010;
assign micromatrizz[61][565] = 9'b111111111;
assign micromatrizz[61][566] = 9'b111111111;
assign micromatrizz[61][567] = 9'b111111111;
assign micromatrizz[61][568] = 9'b111110010;
assign micromatrizz[61][569] = 9'b111110010;
assign micromatrizz[61][570] = 9'b111110010;
assign micromatrizz[61][571] = 9'b111110010;
assign micromatrizz[61][572] = 9'b111110010;
assign micromatrizz[61][573] = 9'b111110011;
assign micromatrizz[61][574] = 9'b111110011;
assign micromatrizz[61][575] = 9'b111110011;
assign micromatrizz[61][576] = 9'b111111111;
assign micromatrizz[61][577] = 9'b111111111;
assign micromatrizz[61][578] = 9'b111111111;
assign micromatrizz[61][579] = 9'b111111111;
assign micromatrizz[61][580] = 9'b111111111;
assign micromatrizz[61][581] = 9'b111110010;
assign micromatrizz[61][582] = 9'b111110011;
assign micromatrizz[61][583] = 9'b111110010;
assign micromatrizz[61][584] = 9'b111110011;
assign micromatrizz[61][585] = 9'b111110011;
assign micromatrizz[61][586] = 9'b111110011;
assign micromatrizz[61][587] = 9'b111110010;
assign micromatrizz[61][588] = 9'b111111111;
assign micromatrizz[61][589] = 9'b111111111;
assign micromatrizz[61][590] = 9'b111111111;
assign micromatrizz[61][591] = 9'b111110111;
assign micromatrizz[61][592] = 9'b111110010;
assign micromatrizz[61][593] = 9'b111110010;
assign micromatrizz[61][594] = 9'b111110010;
assign micromatrizz[61][595] = 9'b111110011;
assign micromatrizz[61][596] = 9'b111110011;
assign micromatrizz[61][597] = 9'b111110011;
assign micromatrizz[61][598] = 9'b111110111;
assign micromatrizz[61][599] = 9'b111111111;
assign micromatrizz[61][600] = 9'b111110111;
assign micromatrizz[61][601] = 9'b111110111;
assign micromatrizz[61][602] = 9'b111110111;
assign micromatrizz[61][603] = 9'b111110111;
assign micromatrizz[61][604] = 9'b111110111;
assign micromatrizz[61][605] = 9'b111110111;
assign micromatrizz[61][606] = 9'b111110111;
assign micromatrizz[61][607] = 9'b111110111;
assign micromatrizz[61][608] = 9'b111111111;
assign micromatrizz[61][609] = 9'b111111111;
assign micromatrizz[61][610] = 9'b111111111;
assign micromatrizz[61][611] = 9'b111111111;
assign micromatrizz[61][612] = 9'b111110010;
assign micromatrizz[61][613] = 9'b111110010;
assign micromatrizz[61][614] = 9'b111110010;
assign micromatrizz[61][615] = 9'b111110010;
assign micromatrizz[61][616] = 9'b111110011;
assign micromatrizz[61][617] = 9'b111110011;
assign micromatrizz[61][618] = 9'b111110011;
assign micromatrizz[61][619] = 9'b111110011;
assign micromatrizz[61][620] = 9'b111110011;
assign micromatrizz[61][621] = 9'b111110011;
assign micromatrizz[61][622] = 9'b111111111;
assign micromatrizz[61][623] = 9'b111111111;
assign micromatrizz[61][624] = 9'b111111111;
assign micromatrizz[61][625] = 9'b111111111;
assign micromatrizz[61][626] = 9'b111111111;
assign micromatrizz[61][627] = 9'b111111111;
assign micromatrizz[61][628] = 9'b111111111;
assign micromatrizz[61][629] = 9'b111111111;
assign micromatrizz[61][630] = 9'b111111111;
assign micromatrizz[61][631] = 9'b111111111;
assign micromatrizz[61][632] = 9'b111111111;
assign micromatrizz[61][633] = 9'b111111111;
assign micromatrizz[61][634] = 9'b111111111;
assign micromatrizz[61][635] = 9'b111111111;
assign micromatrizz[61][636] = 9'b111111111;
assign micromatrizz[61][637] = 9'b111111111;
assign micromatrizz[61][638] = 9'b111111111;
assign micromatrizz[61][639] = 9'b111111111;
assign micromatrizz[62][0] = 9'b111111111;
assign micromatrizz[62][1] = 9'b111111111;
assign micromatrizz[62][2] = 9'b111111111;
assign micromatrizz[62][3] = 9'b111111111;
assign micromatrizz[62][4] = 9'b111111111;
assign micromatrizz[62][5] = 9'b111111111;
assign micromatrizz[62][6] = 9'b111111111;
assign micromatrizz[62][7] = 9'b111111111;
assign micromatrizz[62][8] = 9'b111111111;
assign micromatrizz[62][9] = 9'b111111111;
assign micromatrizz[62][10] = 9'b111110111;
assign micromatrizz[62][11] = 9'b111110010;
assign micromatrizz[62][12] = 9'b111110010;
assign micromatrizz[62][13] = 9'b111110010;
assign micromatrizz[62][14] = 9'b111110011;
assign micromatrizz[62][15] = 9'b111110011;
assign micromatrizz[62][16] = 9'b111110011;
assign micromatrizz[62][17] = 9'b111110011;
assign micromatrizz[62][18] = 9'b111110011;
assign micromatrizz[62][19] = 9'b111110011;
assign micromatrizz[62][20] = 9'b111111111;
assign micromatrizz[62][21] = 9'b111111111;
assign micromatrizz[62][22] = 9'b111111111;
assign micromatrizz[62][23] = 9'b111110111;
assign micromatrizz[62][24] = 9'b111110010;
assign micromatrizz[62][25] = 9'b111110010;
assign micromatrizz[62][26] = 9'b111110010;
assign micromatrizz[62][27] = 9'b111110011;
assign micromatrizz[62][28] = 9'b111110011;
assign micromatrizz[62][29] = 9'b111110011;
assign micromatrizz[62][30] = 9'b111110011;
assign micromatrizz[62][31] = 9'b111111111;
assign micromatrizz[62][32] = 9'b111111111;
assign micromatrizz[62][33] = 9'b111111111;
assign micromatrizz[62][34] = 9'b111111111;
assign micromatrizz[62][35] = 9'b111110111;
assign micromatrizz[62][36] = 9'b111110010;
assign micromatrizz[62][37] = 9'b111110010;
assign micromatrizz[62][38] = 9'b111110011;
assign micromatrizz[62][39] = 9'b111110011;
assign micromatrizz[62][40] = 9'b111110011;
assign micromatrizz[62][41] = 9'b111110011;
assign micromatrizz[62][42] = 9'b111110011;
assign micromatrizz[62][43] = 9'b111111111;
assign micromatrizz[62][44] = 9'b111111111;
assign micromatrizz[62][45] = 9'b111111111;
assign micromatrizz[62][46] = 9'b111111111;
assign micromatrizz[62][47] = 9'b111110010;
assign micromatrizz[62][48] = 9'b111110010;
assign micromatrizz[62][49] = 9'b111110010;
assign micromatrizz[62][50] = 9'b111110011;
assign micromatrizz[62][51] = 9'b111110011;
assign micromatrizz[62][52] = 9'b111110011;
assign micromatrizz[62][53] = 9'b111110010;
assign micromatrizz[62][54] = 9'b111111111;
assign micromatrizz[62][55] = 9'b111111111;
assign micromatrizz[62][56] = 9'b111111111;
assign micromatrizz[62][57] = 9'b111111111;
assign micromatrizz[62][58] = 9'b111111111;
assign micromatrizz[62][59] = 9'b111110010;
assign micromatrizz[62][60] = 9'b111110010;
assign micromatrizz[62][61] = 9'b111110010;
assign micromatrizz[62][62] = 9'b111110011;
assign micromatrizz[62][63] = 9'b111110011;
assign micromatrizz[62][64] = 9'b111110011;
assign micromatrizz[62][65] = 9'b111110010;
assign micromatrizz[62][66] = 9'b111111111;
assign micromatrizz[62][67] = 9'b111111111;
assign micromatrizz[62][68] = 9'b111110111;
assign micromatrizz[62][69] = 9'b111110010;
assign micromatrizz[62][70] = 9'b111110010;
assign micromatrizz[62][71] = 9'b111110010;
assign micromatrizz[62][72] = 9'b111110010;
assign micromatrizz[62][73] = 9'b111110011;
assign micromatrizz[62][74] = 9'b111110011;
assign micromatrizz[62][75] = 9'b111111111;
assign micromatrizz[62][76] = 9'b111111111;
assign micromatrizz[62][77] = 9'b111111111;
assign micromatrizz[62][78] = 9'b111111111;
assign micromatrizz[62][79] = 9'b111111111;
assign micromatrizz[62][80] = 9'b111111111;
assign micromatrizz[62][81] = 9'b111111111;
assign micromatrizz[62][82] = 9'b111111111;
assign micromatrizz[62][83] = 9'b111111111;
assign micromatrizz[62][84] = 9'b111111111;
assign micromatrizz[62][85] = 9'b111111111;
assign micromatrizz[62][86] = 9'b111111111;
assign micromatrizz[62][87] = 9'b111111111;
assign micromatrizz[62][88] = 9'b111110011;
assign micromatrizz[62][89] = 9'b111110010;
assign micromatrizz[62][90] = 9'b111110010;
assign micromatrizz[62][91] = 9'b111110010;
assign micromatrizz[62][92] = 9'b111110011;
assign micromatrizz[62][93] = 9'b111110011;
assign micromatrizz[62][94] = 9'b111110011;
assign micromatrizz[62][95] = 9'b111110111;
assign micromatrizz[62][96] = 9'b111111111;
assign micromatrizz[62][97] = 9'b111111111;
assign micromatrizz[62][98] = 9'b111111111;
assign micromatrizz[62][99] = 9'b111111111;
assign micromatrizz[62][100] = 9'b111111111;
assign micromatrizz[62][101] = 9'b111111111;
assign micromatrizz[62][102] = 9'b111111111;
assign micromatrizz[62][103] = 9'b111111111;
assign micromatrizz[62][104] = 9'b111111111;
assign micromatrizz[62][105] = 9'b111111111;
assign micromatrizz[62][106] = 9'b111110111;
assign micromatrizz[62][107] = 9'b111110010;
assign micromatrizz[62][108] = 9'b111110010;
assign micromatrizz[62][109] = 9'b111110010;
assign micromatrizz[62][110] = 9'b111110011;
assign micromatrizz[62][111] = 9'b111110011;
assign micromatrizz[62][112] = 9'b111110010;
assign micromatrizz[62][113] = 9'b111110011;
assign micromatrizz[62][114] = 9'b111110011;
assign micromatrizz[62][115] = 9'b111110011;
assign micromatrizz[62][116] = 9'b111110111;
assign micromatrizz[62][117] = 9'b111111111;
assign micromatrizz[62][118] = 9'b111111111;
assign micromatrizz[62][119] = 9'b111110010;
assign micromatrizz[62][120] = 9'b111110010;
assign micromatrizz[62][121] = 9'b111110011;
assign micromatrizz[62][122] = 9'b111110010;
assign micromatrizz[62][123] = 9'b111110010;
assign micromatrizz[62][124] = 9'b111110011;
assign micromatrizz[62][125] = 9'b111110011;
assign micromatrizz[62][126] = 9'b111110111;
assign micromatrizz[62][127] = 9'b111111111;
assign micromatrizz[62][128] = 9'b111111111;
assign micromatrizz[62][129] = 9'b111111111;
assign micromatrizz[62][130] = 9'b111111111;
assign micromatrizz[62][131] = 9'b111111111;
assign micromatrizz[62][132] = 9'b111111111;
assign micromatrizz[62][133] = 9'b111111111;
assign micromatrizz[62][134] = 9'b111110111;
assign micromatrizz[62][135] = 9'b111110111;
assign micromatrizz[62][136] = 9'b111111111;
assign micromatrizz[62][137] = 9'b111111111;
assign micromatrizz[62][138] = 9'b111110111;
assign micromatrizz[62][139] = 9'b111110010;
assign micromatrizz[62][140] = 9'b111110010;
assign micromatrizz[62][141] = 9'b111110010;
assign micromatrizz[62][142] = 9'b111110010;
assign micromatrizz[62][143] = 9'b111110011;
assign micromatrizz[62][144] = 9'b111110011;
assign micromatrizz[62][145] = 9'b111110011;
assign micromatrizz[62][146] = 9'b111111111;
assign micromatrizz[62][147] = 9'b111111111;
assign micromatrizz[62][148] = 9'b111111111;
assign micromatrizz[62][149] = 9'b111111111;
assign micromatrizz[62][150] = 9'b111110111;
assign micromatrizz[62][151] = 9'b111110010;
assign micromatrizz[62][152] = 9'b111110010;
assign micromatrizz[62][153] = 9'b111110010;
assign micromatrizz[62][154] = 9'b111110011;
assign micromatrizz[62][155] = 9'b111110011;
assign micromatrizz[62][156] = 9'b111110011;
assign micromatrizz[62][157] = 9'b111110011;
assign micromatrizz[62][158] = 9'b111111111;
assign micromatrizz[62][159] = 9'b111111111;
assign micromatrizz[62][160] = 9'b111111111;
assign micromatrizz[62][161] = 9'b111110010;
assign micromatrizz[62][162] = 9'b111110010;
assign micromatrizz[62][163] = 9'b111110010;
assign micromatrizz[62][164] = 9'b111110011;
assign micromatrizz[62][165] = 9'b111110011;
assign micromatrizz[62][166] = 9'b111110011;
assign micromatrizz[62][167] = 9'b111110011;
assign micromatrizz[62][168] = 9'b111111111;
assign micromatrizz[62][169] = 9'b111111111;
assign micromatrizz[62][170] = 9'b111111111;
assign micromatrizz[62][171] = 9'b111111111;
assign micromatrizz[62][172] = 9'b111110010;
assign micromatrizz[62][173] = 9'b111110010;
assign micromatrizz[62][174] = 9'b111110011;
assign micromatrizz[62][175] = 9'b111110011;
assign micromatrizz[62][176] = 9'b111110011;
assign micromatrizz[62][177] = 9'b111110011;
assign micromatrizz[62][178] = 9'b111110010;
assign micromatrizz[62][179] = 9'b111110111;
assign micromatrizz[62][180] = 9'b111111111;
assign micromatrizz[62][181] = 9'b111111111;
assign micromatrizz[62][182] = 9'b111110111;
assign micromatrizz[62][183] = 9'b111110010;
assign micromatrizz[62][184] = 9'b111110011;
assign micromatrizz[62][185] = 9'b111110011;
assign micromatrizz[62][186] = 9'b111110010;
assign micromatrizz[62][187] = 9'b111110010;
assign micromatrizz[62][188] = 9'b111110011;
assign micromatrizz[62][189] = 9'b111110011;
assign micromatrizz[62][190] = 9'b111110111;
assign micromatrizz[62][191] = 9'b111111111;
assign micromatrizz[62][192] = 9'b111111111;
assign micromatrizz[62][193] = 9'b111111111;
assign micromatrizz[62][194] = 9'b111111111;
assign micromatrizz[62][195] = 9'b111110010;
assign micromatrizz[62][196] = 9'b111110011;
assign micromatrizz[62][197] = 9'b111110011;
assign micromatrizz[62][198] = 9'b111110011;
assign micromatrizz[62][199] = 9'b111110010;
assign micromatrizz[62][200] = 9'b111110010;
assign micromatrizz[62][201] = 9'b111110011;
assign micromatrizz[62][202] = 9'b111110111;
assign micromatrizz[62][203] = 9'b111111111;
assign micromatrizz[62][204] = 9'b111111111;
assign micromatrizz[62][205] = 9'b111111111;
assign micromatrizz[62][206] = 9'b111110010;
assign micromatrizz[62][207] = 9'b111110010;
assign micromatrizz[62][208] = 9'b111110010;
assign micromatrizz[62][209] = 9'b111110010;
assign micromatrizz[62][210] = 9'b111110011;
assign micromatrizz[62][211] = 9'b111110011;
assign micromatrizz[62][212] = 9'b111110011;
assign micromatrizz[62][213] = 9'b111110111;
assign micromatrizz[62][214] = 9'b111111111;
assign micromatrizz[62][215] = 9'b111111111;
assign micromatrizz[62][216] = 9'b111111111;
assign micromatrizz[62][217] = 9'b111111111;
assign micromatrizz[62][218] = 9'b111111111;
assign micromatrizz[62][219] = 9'b111111111;
assign micromatrizz[62][220] = 9'b111111111;
assign micromatrizz[62][221] = 9'b111110111;
assign micromatrizz[62][222] = 9'b111111111;
assign micromatrizz[62][223] = 9'b111111111;
assign micromatrizz[62][224] = 9'b111111111;
assign micromatrizz[62][225] = 9'b111110010;
assign micromatrizz[62][226] = 9'b111110010;
assign micromatrizz[62][227] = 9'b111110010;
assign micromatrizz[62][228] = 9'b111110010;
assign micromatrizz[62][229] = 9'b111110011;
assign micromatrizz[62][230] = 9'b111110011;
assign micromatrizz[62][231] = 9'b111110010;
assign micromatrizz[62][232] = 9'b111110111;
assign micromatrizz[62][233] = 9'b111111111;
assign micromatrizz[62][234] = 9'b111111111;
assign micromatrizz[62][235] = 9'b111111111;
assign micromatrizz[62][236] = 9'b111111111;
assign micromatrizz[62][237] = 9'b111111111;
assign micromatrizz[62][238] = 9'b111111111;
assign micromatrizz[62][239] = 9'b111111111;
assign micromatrizz[62][240] = 9'b111111111;
assign micromatrizz[62][241] = 9'b111110010;
assign micromatrizz[62][242] = 9'b111110010;
assign micromatrizz[62][243] = 9'b111110011;
assign micromatrizz[62][244] = 9'b111110010;
assign micromatrizz[62][245] = 9'b111110010;
assign micromatrizz[62][246] = 9'b111110011;
assign micromatrizz[62][247] = 9'b111110111;
assign micromatrizz[62][248] = 9'b111111111;
assign micromatrizz[62][249] = 9'b111111111;
assign micromatrizz[62][250] = 9'b111111111;
assign micromatrizz[62][251] = 9'b111111111;
assign micromatrizz[62][252] = 9'b111111111;
assign micromatrizz[62][253] = 9'b111111111;
assign micromatrizz[62][254] = 9'b111111111;
assign micromatrizz[62][255] = 9'b111111111;
assign micromatrizz[62][256] = 9'b111111111;
assign micromatrizz[62][257] = 9'b111111111;
assign micromatrizz[62][258] = 9'b111111111;
assign micromatrizz[62][259] = 9'b111111111;
assign micromatrizz[62][260] = 9'b111111111;
assign micromatrizz[62][261] = 9'b111111111;
assign micromatrizz[62][262] = 9'b111110010;
assign micromatrizz[62][263] = 9'b111110010;
assign micromatrizz[62][264] = 9'b111110010;
assign micromatrizz[62][265] = 9'b111110010;
assign micromatrizz[62][266] = 9'b111110010;
assign micromatrizz[62][267] = 9'b111110011;
assign micromatrizz[62][268] = 9'b111110011;
assign micromatrizz[62][269] = 9'b111110011;
assign micromatrizz[62][270] = 9'b111110011;
assign micromatrizz[62][271] = 9'b111110011;
assign micromatrizz[62][272] = 9'b111111111;
assign micromatrizz[62][273] = 9'b111111111;
assign micromatrizz[62][274] = 9'b111111111;
assign micromatrizz[62][275] = 9'b111110010;
assign micromatrizz[62][276] = 9'b111110010;
assign micromatrizz[62][277] = 9'b111110010;
assign micromatrizz[62][278] = 9'b111110010;
assign micromatrizz[62][279] = 9'b111110011;
assign micromatrizz[62][280] = 9'b111110011;
assign micromatrizz[62][281] = 9'b111110011;
assign micromatrizz[62][282] = 9'b111111111;
assign micromatrizz[62][283] = 9'b111111111;
assign micromatrizz[62][284] = 9'b111111111;
assign micromatrizz[62][285] = 9'b111111111;
assign micromatrizz[62][286] = 9'b111110010;
assign micromatrizz[62][287] = 9'b111110010;
assign micromatrizz[62][288] = 9'b111110011;
assign micromatrizz[62][289] = 9'b111110011;
assign micromatrizz[62][290] = 9'b111110011;
assign micromatrizz[62][291] = 9'b111110011;
assign micromatrizz[62][292] = 9'b111110011;
assign micromatrizz[62][293] = 9'b111111111;
assign micromatrizz[62][294] = 9'b111111111;
assign micromatrizz[62][295] = 9'b111111111;
assign micromatrizz[62][296] = 9'b111111111;
assign micromatrizz[62][297] = 9'b111111111;
assign micromatrizz[62][298] = 9'b111111111;
assign micromatrizz[62][299] = 9'b111111111;
assign micromatrizz[62][300] = 9'b111111111;
assign micromatrizz[62][301] = 9'b111110010;
assign micromatrizz[62][302] = 9'b111110010;
assign micromatrizz[62][303] = 9'b111110010;
assign micromatrizz[62][304] = 9'b111110011;
assign micromatrizz[62][305] = 9'b111110010;
assign micromatrizz[62][306] = 9'b111110010;
assign micromatrizz[62][307] = 9'b111110011;
assign micromatrizz[62][308] = 9'b111110011;
assign micromatrizz[62][309] = 9'b111110111;
assign micromatrizz[62][310] = 9'b111111111;
assign micromatrizz[62][311] = 9'b111111111;
assign micromatrizz[62][312] = 9'b111111111;
assign micromatrizz[62][313] = 9'b111111111;
assign micromatrizz[62][314] = 9'b111111111;
assign micromatrizz[62][315] = 9'b111110111;
assign micromatrizz[62][316] = 9'b111110010;
assign micromatrizz[62][317] = 9'b111110010;
assign micromatrizz[62][318] = 9'b111110011;
assign micromatrizz[62][319] = 9'b111110010;
assign micromatrizz[62][320] = 9'b111110011;
assign micromatrizz[62][321] = 9'b111110011;
assign micromatrizz[62][322] = 9'b111110111;
assign micromatrizz[62][323] = 9'b111111111;
assign micromatrizz[62][324] = 9'b111111111;
assign micromatrizz[62][325] = 9'b111111111;
assign micromatrizz[62][326] = 9'b111111111;
assign micromatrizz[62][327] = 9'b111111111;
assign micromatrizz[62][328] = 9'b111111111;
assign micromatrizz[62][329] = 9'b111111111;
assign micromatrizz[62][330] = 9'b111111111;
assign micromatrizz[62][331] = 9'b111111111;
assign micromatrizz[62][332] = 9'b111111111;
assign micromatrizz[62][333] = 9'b111111111;
assign micromatrizz[62][334] = 9'b111111111;
assign micromatrizz[62][335] = 9'b111110010;
assign micromatrizz[62][336] = 9'b111110010;
assign micromatrizz[62][337] = 9'b111110011;
assign micromatrizz[62][338] = 9'b111110011;
assign micromatrizz[62][339] = 9'b111110010;
assign micromatrizz[62][340] = 9'b111110011;
assign micromatrizz[62][341] = 9'b111110011;
assign micromatrizz[62][342] = 9'b111111111;
assign micromatrizz[62][343] = 9'b111111111;
assign micromatrizz[62][344] = 9'b111111111;
assign micromatrizz[62][345] = 9'b111111111;
assign micromatrizz[62][346] = 9'b111111111;
assign micromatrizz[62][347] = 9'b111110010;
assign micromatrizz[62][348] = 9'b111110010;
assign micromatrizz[62][349] = 9'b111110010;
assign micromatrizz[62][350] = 9'b111110010;
assign micromatrizz[62][351] = 9'b111110011;
assign micromatrizz[62][352] = 9'b111110011;
assign micromatrizz[62][353] = 9'b111110011;
assign micromatrizz[62][354] = 9'b111111111;
assign micromatrizz[62][355] = 9'b111111111;
assign micromatrizz[62][356] = 9'b111111111;
assign micromatrizz[62][357] = 9'b111111111;
assign micromatrizz[62][358] = 9'b111111111;
assign micromatrizz[62][359] = 9'b111110010;
assign micromatrizz[62][360] = 9'b111110011;
assign micromatrizz[62][361] = 9'b111110010;
assign micromatrizz[62][362] = 9'b111110010;
assign micromatrizz[62][363] = 9'b111110011;
assign micromatrizz[62][364] = 9'b111110011;
assign micromatrizz[62][365] = 9'b111110011;
assign micromatrizz[62][366] = 9'b111111111;
assign micromatrizz[62][367] = 9'b111111111;
assign micromatrizz[62][368] = 9'b111111111;
assign micromatrizz[62][369] = 9'b111111111;
assign micromatrizz[62][370] = 9'b111111111;
assign micromatrizz[62][371] = 9'b111111111;
assign micromatrizz[62][372] = 9'b111110010;
assign micromatrizz[62][373] = 9'b111110011;
assign micromatrizz[62][374] = 9'b111110011;
assign micromatrizz[62][375] = 9'b111110011;
assign micromatrizz[62][376] = 9'b111110011;
assign micromatrizz[62][377] = 9'b111110011;
assign micromatrizz[62][378] = 9'b111110011;
assign micromatrizz[62][379] = 9'b111111111;
assign micromatrizz[62][380] = 9'b111111111;
assign micromatrizz[62][381] = 9'b111111111;
assign micromatrizz[62][382] = 9'b111111111;
assign micromatrizz[62][383] = 9'b111111111;
assign micromatrizz[62][384] = 9'b111110010;
assign micromatrizz[62][385] = 9'b111110010;
assign micromatrizz[62][386] = 9'b111110011;
assign micromatrizz[62][387] = 9'b111110011;
assign micromatrizz[62][388] = 9'b111110011;
assign micromatrizz[62][389] = 9'b111110011;
assign micromatrizz[62][390] = 9'b111110011;
assign micromatrizz[62][391] = 9'b111111111;
assign micromatrizz[62][392] = 9'b111111111;
assign micromatrizz[62][393] = 9'b111111111;
assign micromatrizz[62][394] = 9'b111111111;
assign micromatrizz[62][395] = 9'b111110110;
assign micromatrizz[62][396] = 9'b111110010;
assign micromatrizz[62][397] = 9'b111110010;
assign micromatrizz[62][398] = 9'b111110010;
assign micromatrizz[62][399] = 9'b111110010;
assign micromatrizz[62][400] = 9'b111110011;
assign micromatrizz[62][401] = 9'b111110011;
assign micromatrizz[62][402] = 9'b111110111;
assign micromatrizz[62][403] = 9'b111111111;
assign micromatrizz[62][404] = 9'b111111111;
assign micromatrizz[62][405] = 9'b111111111;
assign micromatrizz[62][406] = 9'b111111111;
assign micromatrizz[62][407] = 9'b111111111;
assign micromatrizz[62][408] = 9'b111111111;
assign micromatrizz[62][409] = 9'b111111111;
assign micromatrizz[62][410] = 9'b111111111;
assign micromatrizz[62][411] = 9'b111110010;
assign micromatrizz[62][412] = 9'b111110010;
assign micromatrizz[62][413] = 9'b111110010;
assign micromatrizz[62][414] = 9'b111110010;
assign micromatrizz[62][415] = 9'b111110011;
assign micromatrizz[62][416] = 9'b111110010;
assign micromatrizz[62][417] = 9'b111110111;
assign micromatrizz[62][418] = 9'b111111111;
assign micromatrizz[62][419] = 9'b111111111;
assign micromatrizz[62][420] = 9'b111111111;
assign micromatrizz[62][421] = 9'b111111111;
assign micromatrizz[62][422] = 9'b111111111;
assign micromatrizz[62][423] = 9'b111111111;
assign micromatrizz[62][424] = 9'b111111111;
assign micromatrizz[62][425] = 9'b111111111;
assign micromatrizz[62][426] = 9'b111111111;
assign micromatrizz[62][427] = 9'b111111111;
assign micromatrizz[62][428] = 9'b111111111;
assign micromatrizz[62][429] = 9'b111111111;
assign micromatrizz[62][430] = 9'b111110111;
assign micromatrizz[62][431] = 9'b111110010;
assign micromatrizz[62][432] = 9'b111110010;
assign micromatrizz[62][433] = 9'b111110010;
assign micromatrizz[62][434] = 9'b111110010;
assign micromatrizz[62][435] = 9'b111110011;
assign micromatrizz[62][436] = 9'b111110011;
assign micromatrizz[62][437] = 9'b111110011;
assign micromatrizz[62][438] = 9'b111111111;
assign micromatrizz[62][439] = 9'b111111111;
assign micromatrizz[62][440] = 9'b111111111;
assign micromatrizz[62][441] = 9'b111111111;
assign micromatrizz[62][442] = 9'b111111111;
assign micromatrizz[62][443] = 9'b111111111;
assign micromatrizz[62][444] = 9'b111111111;
assign micromatrizz[62][445] = 9'b111111111;
assign micromatrizz[62][446] = 9'b111110110;
assign micromatrizz[62][447] = 9'b111110010;
assign micromatrizz[62][448] = 9'b111110010;
assign micromatrizz[62][449] = 9'b111110010;
assign micromatrizz[62][450] = 9'b111110010;
assign micromatrizz[62][451] = 9'b111110011;
assign micromatrizz[62][452] = 9'b111110011;
assign micromatrizz[62][453] = 9'b111110011;
assign micromatrizz[62][454] = 9'b111111111;
assign micromatrizz[62][455] = 9'b111111111;
assign micromatrizz[62][456] = 9'b111111111;
assign micromatrizz[62][457] = 9'b111111111;
assign micromatrizz[62][458] = 9'b111111111;
assign micromatrizz[62][459] = 9'b111111111;
assign micromatrizz[62][460] = 9'b111111111;
assign micromatrizz[62][461] = 9'b111111111;
assign micromatrizz[62][462] = 9'b111110111;
assign micromatrizz[62][463] = 9'b111111111;
assign micromatrizz[62][464] = 9'b111111111;
assign micromatrizz[62][465] = 9'b111111111;
assign micromatrizz[62][466] = 9'b111111111;
assign micromatrizz[62][467] = 9'b111110110;
assign micromatrizz[62][468] = 9'b111110010;
assign micromatrizz[62][469] = 9'b111110010;
assign micromatrizz[62][470] = 9'b111110010;
assign micromatrizz[62][471] = 9'b111110011;
assign micromatrizz[62][472] = 9'b111110011;
assign micromatrizz[62][473] = 9'b111110011;
assign micromatrizz[62][474] = 9'b111110011;
assign micromatrizz[62][475] = 9'b111110011;
assign micromatrizz[62][476] = 9'b111110011;
assign micromatrizz[62][477] = 9'b111111111;
assign micromatrizz[62][478] = 9'b111111111;
assign micromatrizz[62][479] = 9'b111111111;
assign micromatrizz[62][480] = 9'b111111111;
assign micromatrizz[62][481] = 9'b111110010;
assign micromatrizz[62][482] = 9'b111110010;
assign micromatrizz[62][483] = 9'b111110010;
assign micromatrizz[62][484] = 9'b111110010;
assign micromatrizz[62][485] = 9'b111110011;
assign micromatrizz[62][486] = 9'b111110011;
assign micromatrizz[62][487] = 9'b111110011;
assign micromatrizz[62][488] = 9'b111110111;
assign micromatrizz[62][489] = 9'b111111111;
assign micromatrizz[62][490] = 9'b111111111;
assign micromatrizz[62][491] = 9'b111111111;
assign micromatrizz[62][492] = 9'b111111111;
assign micromatrizz[62][493] = 9'b111111111;
assign micromatrizz[62][494] = 9'b111111111;
assign micromatrizz[62][495] = 9'b111111111;
assign micromatrizz[62][496] = 9'b111111111;
assign micromatrizz[62][497] = 9'b111110010;
assign micromatrizz[62][498] = 9'b111110010;
assign micromatrizz[62][499] = 9'b111110010;
assign micromatrizz[62][500] = 9'b111110011;
assign micromatrizz[62][501] = 9'b111110010;
assign micromatrizz[62][502] = 9'b111110010;
assign micromatrizz[62][503] = 9'b111110111;
assign micromatrizz[62][504] = 9'b111111111;
assign micromatrizz[62][505] = 9'b111111111;
assign micromatrizz[62][506] = 9'b111111111;
assign micromatrizz[62][507] = 9'b111111111;
assign micromatrizz[62][508] = 9'b111111111;
assign micromatrizz[62][509] = 9'b111111111;
assign micromatrizz[62][510] = 9'b111111111;
assign micromatrizz[62][511] = 9'b111111111;
assign micromatrizz[62][512] = 9'b111111111;
assign micromatrizz[62][513] = 9'b111111111;
assign micromatrizz[62][514] = 9'b111111111;
assign micromatrizz[62][515] = 9'b111111111;
assign micromatrizz[62][516] = 9'b111110111;
assign micromatrizz[62][517] = 9'b111110011;
assign micromatrizz[62][518] = 9'b111110011;
assign micromatrizz[62][519] = 9'b111110011;
assign micromatrizz[62][520] = 9'b111110010;
assign micromatrizz[62][521] = 9'b111110010;
assign micromatrizz[62][522] = 9'b111110011;
assign micromatrizz[62][523] = 9'b111110111;
assign micromatrizz[62][524] = 9'b111111111;
assign micromatrizz[62][525] = 9'b111111111;
assign micromatrizz[62][526] = 9'b111111111;
assign micromatrizz[62][527] = 9'b111111111;
assign micromatrizz[62][528] = 9'b111111111;
assign micromatrizz[62][529] = 9'b111110010;
assign micromatrizz[62][530] = 9'b111110010;
assign micromatrizz[62][531] = 9'b111110010;
assign micromatrizz[62][532] = 9'b111110011;
assign micromatrizz[62][533] = 9'b111110011;
assign micromatrizz[62][534] = 9'b111110011;
assign micromatrizz[62][535] = 9'b111110011;
assign micromatrizz[62][536] = 9'b111111111;
assign micromatrizz[62][537] = 9'b111111111;
assign micromatrizz[62][538] = 9'b111110111;
assign micromatrizz[62][539] = 9'b111110010;
assign micromatrizz[62][540] = 9'b111110010;
assign micromatrizz[62][541] = 9'b111110010;
assign micromatrizz[62][542] = 9'b111110011;
assign micromatrizz[62][543] = 9'b111110011;
assign micromatrizz[62][544] = 9'b111110010;
assign micromatrizz[62][545] = 9'b111111111;
assign micromatrizz[62][546] = 9'b111111111;
assign micromatrizz[62][547] = 9'b111111111;
assign micromatrizz[62][548] = 9'b111111111;
assign micromatrizz[62][549] = 9'b111111111;
assign micromatrizz[62][550] = 9'b111111111;
assign micromatrizz[62][551] = 9'b111111111;
assign micromatrizz[62][552] = 9'b111111111;
assign micromatrizz[62][553] = 9'b111111111;
assign micromatrizz[62][554] = 9'b111111111;
assign micromatrizz[62][555] = 9'b111111111;
assign micromatrizz[62][556] = 9'b111111111;
assign micromatrizz[62][557] = 9'b111111111;
assign micromatrizz[62][558] = 9'b111110010;
assign micromatrizz[62][559] = 9'b111110010;
assign micromatrizz[62][560] = 9'b111110010;
assign micromatrizz[62][561] = 9'b111110010;
assign micromatrizz[62][562] = 9'b111110011;
assign micromatrizz[62][563] = 9'b111110010;
assign micromatrizz[62][564] = 9'b111110010;
assign micromatrizz[62][565] = 9'b111111111;
assign micromatrizz[62][566] = 9'b111111111;
assign micromatrizz[62][567] = 9'b111111111;
assign micromatrizz[62][568] = 9'b111110111;
assign micromatrizz[62][569] = 9'b111110010;
assign micromatrizz[62][570] = 9'b111110010;
assign micromatrizz[62][571] = 9'b111110010;
assign micromatrizz[62][572] = 9'b111110010;
assign micromatrizz[62][573] = 9'b111110011;
assign micromatrizz[62][574] = 9'b111110011;
assign micromatrizz[62][575] = 9'b111110011;
assign micromatrizz[62][576] = 9'b111111111;
assign micromatrizz[62][577] = 9'b111111111;
assign micromatrizz[62][578] = 9'b111111111;
assign micromatrizz[62][579] = 9'b111111111;
assign micromatrizz[62][580] = 9'b111111111;
assign micromatrizz[62][581] = 9'b111110010;
assign micromatrizz[62][582] = 9'b111110011;
assign micromatrizz[62][583] = 9'b111110011;
assign micromatrizz[62][584] = 9'b111110011;
assign micromatrizz[62][585] = 9'b111110011;
assign micromatrizz[62][586] = 9'b111110011;
assign micromatrizz[62][587] = 9'b111110010;
assign micromatrizz[62][588] = 9'b111111111;
assign micromatrizz[62][589] = 9'b111111111;
assign micromatrizz[62][590] = 9'b111111111;
assign micromatrizz[62][591] = 9'b111110111;
assign micromatrizz[62][592] = 9'b111110010;
assign micromatrizz[62][593] = 9'b111110010;
assign micromatrizz[62][594] = 9'b111110010;
assign micromatrizz[62][595] = 9'b111110011;
assign micromatrizz[62][596] = 9'b111110011;
assign micromatrizz[62][597] = 9'b111110011;
assign micromatrizz[62][598] = 9'b111111111;
assign micromatrizz[62][599] = 9'b111111111;
assign micromatrizz[62][600] = 9'b111111111;
assign micromatrizz[62][601] = 9'b111111111;
assign micromatrizz[62][602] = 9'b111111111;
assign micromatrizz[62][603] = 9'b111111111;
assign micromatrizz[62][604] = 9'b111111111;
assign micromatrizz[62][605] = 9'b111111111;
assign micromatrizz[62][606] = 9'b111111111;
assign micromatrizz[62][607] = 9'b111111111;
assign micromatrizz[62][608] = 9'b111111111;
assign micromatrizz[62][609] = 9'b111111111;
assign micromatrizz[62][610] = 9'b111111111;
assign micromatrizz[62][611] = 9'b111111111;
assign micromatrizz[62][612] = 9'b111110111;
assign micromatrizz[62][613] = 9'b111110010;
assign micromatrizz[62][614] = 9'b111110010;
assign micromatrizz[62][615] = 9'b111110010;
assign micromatrizz[62][616] = 9'b111110011;
assign micromatrizz[62][617] = 9'b111110011;
assign micromatrizz[62][618] = 9'b111110011;
assign micromatrizz[62][619] = 9'b111110011;
assign micromatrizz[62][620] = 9'b111110011;
assign micromatrizz[62][621] = 9'b111110011;
assign micromatrizz[62][622] = 9'b111110111;
assign micromatrizz[62][623] = 9'b111111111;
assign micromatrizz[62][624] = 9'b111111111;
assign micromatrizz[62][625] = 9'b111111111;
assign micromatrizz[62][626] = 9'b111111111;
assign micromatrizz[62][627] = 9'b111111111;
assign micromatrizz[62][628] = 9'b111111111;
assign micromatrizz[62][629] = 9'b111111111;
assign micromatrizz[62][630] = 9'b111111111;
assign micromatrizz[62][631] = 9'b111111111;
assign micromatrizz[62][632] = 9'b111111111;
assign micromatrizz[62][633] = 9'b111111111;
assign micromatrizz[62][634] = 9'b111111111;
assign micromatrizz[62][635] = 9'b111111111;
assign micromatrizz[62][636] = 9'b111111111;
assign micromatrizz[62][637] = 9'b111111111;
assign micromatrizz[62][638] = 9'b111111111;
assign micromatrizz[62][639] = 9'b111111111;
assign micromatrizz[63][0] = 9'b111111111;
assign micromatrizz[63][1] = 9'b111111111;
assign micromatrizz[63][2] = 9'b111111111;
assign micromatrizz[63][3] = 9'b111111111;
assign micromatrizz[63][4] = 9'b111111111;
assign micromatrizz[63][5] = 9'b111111111;
assign micromatrizz[63][6] = 9'b111111111;
assign micromatrizz[63][7] = 9'b111111111;
assign micromatrizz[63][8] = 9'b111111111;
assign micromatrizz[63][9] = 9'b111111111;
assign micromatrizz[63][10] = 9'b111111111;
assign micromatrizz[63][11] = 9'b111110010;
assign micromatrizz[63][12] = 9'b111110010;
assign micromatrizz[63][13] = 9'b111110010;
assign micromatrizz[63][14] = 9'b111110010;
assign micromatrizz[63][15] = 9'b111110011;
assign micromatrizz[63][16] = 9'b111110011;
assign micromatrizz[63][17] = 9'b111110011;
assign micromatrizz[63][18] = 9'b111110011;
assign micromatrizz[63][19] = 9'b111110010;
assign micromatrizz[63][20] = 9'b111110111;
assign micromatrizz[63][21] = 9'b111111111;
assign micromatrizz[63][22] = 9'b111111111;
assign micromatrizz[63][23] = 9'b111110111;
assign micromatrizz[63][24] = 9'b111110010;
assign micromatrizz[63][25] = 9'b111110010;
assign micromatrizz[63][26] = 9'b111110010;
assign micromatrizz[63][27] = 9'b111110011;
assign micromatrizz[63][28] = 9'b111110011;
assign micromatrizz[63][29] = 9'b111110011;
assign micromatrizz[63][30] = 9'b111110011;
assign micromatrizz[63][31] = 9'b111111111;
assign micromatrizz[63][32] = 9'b111111111;
assign micromatrizz[63][33] = 9'b111111111;
assign micromatrizz[63][34] = 9'b111111111;
assign micromatrizz[63][35] = 9'b111110111;
assign micromatrizz[63][36] = 9'b111110010;
assign micromatrizz[63][37] = 9'b111110011;
assign micromatrizz[63][38] = 9'b111110011;
assign micromatrizz[63][39] = 9'b111110011;
assign micromatrizz[63][40] = 9'b111110011;
assign micromatrizz[63][41] = 9'b111110011;
assign micromatrizz[63][42] = 9'b111110011;
assign micromatrizz[63][43] = 9'b111111111;
assign micromatrizz[63][44] = 9'b111111111;
assign micromatrizz[63][45] = 9'b111111111;
assign micromatrizz[63][46] = 9'b111111111;
assign micromatrizz[63][47] = 9'b111110010;
assign micromatrizz[63][48] = 9'b111110010;
assign micromatrizz[63][49] = 9'b111110010;
assign micromatrizz[63][50] = 9'b111110011;
assign micromatrizz[63][51] = 9'b111110011;
assign micromatrizz[63][52] = 9'b111110011;
assign micromatrizz[63][53] = 9'b111110011;
assign micromatrizz[63][54] = 9'b111111111;
assign micromatrizz[63][55] = 9'b111111111;
assign micromatrizz[63][56] = 9'b111111111;
assign micromatrizz[63][57] = 9'b111111111;
assign micromatrizz[63][58] = 9'b111111111;
assign micromatrizz[63][59] = 9'b111110010;
assign micromatrizz[63][60] = 9'b111110010;
assign micromatrizz[63][61] = 9'b111110010;
assign micromatrizz[63][62] = 9'b111110011;
assign micromatrizz[63][63] = 9'b111110011;
assign micromatrizz[63][64] = 9'b111110011;
assign micromatrizz[63][65] = 9'b111110011;
assign micromatrizz[63][66] = 9'b111111111;
assign micromatrizz[63][67] = 9'b111111111;
assign micromatrizz[63][68] = 9'b111110111;
assign micromatrizz[63][69] = 9'b111110010;
assign micromatrizz[63][70] = 9'b111110010;
assign micromatrizz[63][71] = 9'b111110010;
assign micromatrizz[63][72] = 9'b111110011;
assign micromatrizz[63][73] = 9'b111110011;
assign micromatrizz[63][74] = 9'b111110011;
assign micromatrizz[63][75] = 9'b111111111;
assign micromatrizz[63][76] = 9'b111111111;
assign micromatrizz[63][77] = 9'b111111111;
assign micromatrizz[63][78] = 9'b111111111;
assign micromatrizz[63][79] = 9'b111111111;
assign micromatrizz[63][80] = 9'b111111111;
assign micromatrizz[63][81] = 9'b111111111;
assign micromatrizz[63][82] = 9'b111111111;
assign micromatrizz[63][83] = 9'b111111111;
assign micromatrizz[63][84] = 9'b111111111;
assign micromatrizz[63][85] = 9'b111111111;
assign micromatrizz[63][86] = 9'b111111111;
assign micromatrizz[63][87] = 9'b111111111;
assign micromatrizz[63][88] = 9'b111110110;
assign micromatrizz[63][89] = 9'b111110010;
assign micromatrizz[63][90] = 9'b111110010;
assign micromatrizz[63][91] = 9'b111110011;
assign micromatrizz[63][92] = 9'b111110011;
assign micromatrizz[63][93] = 9'b111110011;
assign micromatrizz[63][94] = 9'b111110011;
assign micromatrizz[63][95] = 9'b111110111;
assign micromatrizz[63][96] = 9'b111111111;
assign micromatrizz[63][97] = 9'b111111111;
assign micromatrizz[63][98] = 9'b111111111;
assign micromatrizz[63][99] = 9'b111111111;
assign micromatrizz[63][100] = 9'b111111111;
assign micromatrizz[63][101] = 9'b111111111;
assign micromatrizz[63][102] = 9'b111111111;
assign micromatrizz[63][103] = 9'b111111111;
assign micromatrizz[63][104] = 9'b111111111;
assign micromatrizz[63][105] = 9'b111111111;
assign micromatrizz[63][106] = 9'b111111111;
assign micromatrizz[63][107] = 9'b111110111;
assign micromatrizz[63][108] = 9'b111110010;
assign micromatrizz[63][109] = 9'b111110011;
assign micromatrizz[63][110] = 9'b111110010;
assign micromatrizz[63][111] = 9'b111110011;
assign micromatrizz[63][112] = 9'b111110011;
assign micromatrizz[63][113] = 9'b111110011;
assign micromatrizz[63][114] = 9'b111110011;
assign micromatrizz[63][115] = 9'b111110011;
assign micromatrizz[63][116] = 9'b111110011;
assign micromatrizz[63][117] = 9'b111111111;
assign micromatrizz[63][118] = 9'b111111111;
assign micromatrizz[63][119] = 9'b111110111;
assign micromatrizz[63][120] = 9'b111110010;
assign micromatrizz[63][121] = 9'b111110010;
assign micromatrizz[63][122] = 9'b111110010;
assign micromatrizz[63][123] = 9'b111110010;
assign micromatrizz[63][124] = 9'b111110011;
assign micromatrizz[63][125] = 9'b111110011;
assign micromatrizz[63][126] = 9'b111110111;
assign micromatrizz[63][127] = 9'b111111111;
assign micromatrizz[63][128] = 9'b111111111;
assign micromatrizz[63][129] = 9'b111111111;
assign micromatrizz[63][130] = 9'b111111111;
assign micromatrizz[63][131] = 9'b111111111;
assign micromatrizz[63][132] = 9'b111111111;
assign micromatrizz[63][133] = 9'b111111111;
assign micromatrizz[63][134] = 9'b111110111;
assign micromatrizz[63][135] = 9'b111111111;
assign micromatrizz[63][136] = 9'b111111111;
assign micromatrizz[63][137] = 9'b111111111;
assign micromatrizz[63][138] = 9'b111110111;
assign micromatrizz[63][139] = 9'b111110010;
assign micromatrizz[63][140] = 9'b111110010;
assign micromatrizz[63][141] = 9'b111110010;
assign micromatrizz[63][142] = 9'b111110010;
assign micromatrizz[63][143] = 9'b111110011;
assign micromatrizz[63][144] = 9'b111110011;
assign micromatrizz[63][145] = 9'b111110011;
assign micromatrizz[63][146] = 9'b111111111;
assign micromatrizz[63][147] = 9'b111111111;
assign micromatrizz[63][148] = 9'b111111111;
assign micromatrizz[63][149] = 9'b111111111;
assign micromatrizz[63][150] = 9'b111110111;
assign micromatrizz[63][151] = 9'b111110010;
assign micromatrizz[63][152] = 9'b111110010;
assign micromatrizz[63][153] = 9'b111110011;
assign micromatrizz[63][154] = 9'b111110011;
assign micromatrizz[63][155] = 9'b111110011;
assign micromatrizz[63][156] = 9'b111110011;
assign micromatrizz[63][157] = 9'b111110111;
assign micromatrizz[63][158] = 9'b111111111;
assign micromatrizz[63][159] = 9'b111111111;
assign micromatrizz[63][160] = 9'b111111111;
assign micromatrizz[63][161] = 9'b111110010;
assign micromatrizz[63][162] = 9'b111110010;
assign micromatrizz[63][163] = 9'b111110010;
assign micromatrizz[63][164] = 9'b111110011;
assign micromatrizz[63][165] = 9'b111110010;
assign micromatrizz[63][166] = 9'b111110011;
assign micromatrizz[63][167] = 9'b111110011;
assign micromatrizz[63][168] = 9'b111111111;
assign micromatrizz[63][169] = 9'b111111111;
assign micromatrizz[63][170] = 9'b111111111;
assign micromatrizz[63][171] = 9'b111111111;
assign micromatrizz[63][172] = 9'b111110010;
assign micromatrizz[63][173] = 9'b111110011;
assign micromatrizz[63][174] = 9'b111110011;
assign micromatrizz[63][175] = 9'b111110011;
assign micromatrizz[63][176] = 9'b111110011;
assign micromatrizz[63][177] = 9'b111110011;
assign micromatrizz[63][178] = 9'b111110010;
assign micromatrizz[63][179] = 9'b111110111;
assign micromatrizz[63][180] = 9'b111111111;
assign micromatrizz[63][181] = 9'b111111111;
assign micromatrizz[63][182] = 9'b111111111;
assign micromatrizz[63][183] = 9'b111110010;
assign micromatrizz[63][184] = 9'b111110011;
assign micromatrizz[63][185] = 9'b111110011;
assign micromatrizz[63][186] = 9'b111110010;
assign micromatrizz[63][187] = 9'b111110010;
assign micromatrizz[63][188] = 9'b111110011;
assign micromatrizz[63][189] = 9'b111110011;
assign micromatrizz[63][190] = 9'b111111111;
assign micromatrizz[63][191] = 9'b111111111;
assign micromatrizz[63][192] = 9'b111111111;
assign micromatrizz[63][193] = 9'b111111111;
assign micromatrizz[63][194] = 9'b111111111;
assign micromatrizz[63][195] = 9'b111110010;
assign micromatrizz[63][196] = 9'b111110010;
assign micromatrizz[63][197] = 9'b111110011;
assign micromatrizz[63][198] = 9'b111110011;
assign micromatrizz[63][199] = 9'b111110010;
assign micromatrizz[63][200] = 9'b111110010;
assign micromatrizz[63][201] = 9'b111110011;
assign micromatrizz[63][202] = 9'b111110111;
assign micromatrizz[63][203] = 9'b111111111;
assign micromatrizz[63][204] = 9'b111111111;
assign micromatrizz[63][205] = 9'b111111111;
assign micromatrizz[63][206] = 9'b111110010;
assign micromatrizz[63][207] = 9'b111110010;
assign micromatrizz[63][208] = 9'b111110010;
assign micromatrizz[63][209] = 9'b111110010;
assign micromatrizz[63][210] = 9'b111110011;
assign micromatrizz[63][211] = 9'b111110011;
assign micromatrizz[63][212] = 9'b111110011;
assign micromatrizz[63][213] = 9'b111110111;
assign micromatrizz[63][214] = 9'b111111111;
assign micromatrizz[63][215] = 9'b111111111;
assign micromatrizz[63][216] = 9'b111111111;
assign micromatrizz[63][217] = 9'b111111111;
assign micromatrizz[63][218] = 9'b111111111;
assign micromatrizz[63][219] = 9'b111111111;
assign micromatrizz[63][220] = 9'b111111111;
assign micromatrizz[63][221] = 9'b111110110;
assign micromatrizz[63][222] = 9'b111111111;
assign micromatrizz[63][223] = 9'b111111111;
assign micromatrizz[63][224] = 9'b111111111;
assign micromatrizz[63][225] = 9'b111110010;
assign micromatrizz[63][226] = 9'b111110010;
assign micromatrizz[63][227] = 9'b111110010;
assign micromatrizz[63][228] = 9'b111110010;
assign micromatrizz[63][229] = 9'b111110011;
assign micromatrizz[63][230] = 9'b111110011;
assign micromatrizz[63][231] = 9'b111110011;
assign micromatrizz[63][232] = 9'b111110111;
assign micromatrizz[63][233] = 9'b111111111;
assign micromatrizz[63][234] = 9'b111111111;
assign micromatrizz[63][235] = 9'b111111111;
assign micromatrizz[63][236] = 9'b111111111;
assign micromatrizz[63][237] = 9'b111111111;
assign micromatrizz[63][238] = 9'b111111111;
assign micromatrizz[63][239] = 9'b111111111;
assign micromatrizz[63][240] = 9'b111111111;
assign micromatrizz[63][241] = 9'b111110010;
assign micromatrizz[63][242] = 9'b111110010;
assign micromatrizz[63][243] = 9'b111110010;
assign micromatrizz[63][244] = 9'b111110010;
assign micromatrizz[63][245] = 9'b111110011;
assign micromatrizz[63][246] = 9'b111110011;
assign micromatrizz[63][247] = 9'b111110111;
assign micromatrizz[63][248] = 9'b111111111;
assign micromatrizz[63][249] = 9'b111111111;
assign micromatrizz[63][250] = 9'b111111111;
assign micromatrizz[63][251] = 9'b111111111;
assign micromatrizz[63][252] = 9'b111111111;
assign micromatrizz[63][253] = 9'b111111111;
assign micromatrizz[63][254] = 9'b111111111;
assign micromatrizz[63][255] = 9'b111111111;
assign micromatrizz[63][256] = 9'b111111111;
assign micromatrizz[63][257] = 9'b111111111;
assign micromatrizz[63][258] = 9'b111111111;
assign micromatrizz[63][259] = 9'b111111111;
assign micromatrizz[63][260] = 9'b111111111;
assign micromatrizz[63][261] = 9'b111111111;
assign micromatrizz[63][262] = 9'b111111111;
assign micromatrizz[63][263] = 9'b111110010;
assign micromatrizz[63][264] = 9'b111110010;
assign micromatrizz[63][265] = 9'b111110010;
assign micromatrizz[63][266] = 9'b111110010;
assign micromatrizz[63][267] = 9'b111110011;
assign micromatrizz[63][268] = 9'b111110011;
assign micromatrizz[63][269] = 9'b111110011;
assign micromatrizz[63][270] = 9'b111110011;
assign micromatrizz[63][271] = 9'b111110011;
assign micromatrizz[63][272] = 9'b111110111;
assign micromatrizz[63][273] = 9'b111111111;
assign micromatrizz[63][274] = 9'b111110111;
assign micromatrizz[63][275] = 9'b111110010;
assign micromatrizz[63][276] = 9'b111110010;
assign micromatrizz[63][277] = 9'b111110010;
assign micromatrizz[63][278] = 9'b111110011;
assign micromatrizz[63][279] = 9'b111110011;
assign micromatrizz[63][280] = 9'b111110011;
assign micromatrizz[63][281] = 9'b111110011;
assign micromatrizz[63][282] = 9'b111111111;
assign micromatrizz[63][283] = 9'b111111111;
assign micromatrizz[63][284] = 9'b111111111;
assign micromatrizz[63][285] = 9'b111111111;
assign micromatrizz[63][286] = 9'b111110010;
assign micromatrizz[63][287] = 9'b111110010;
assign micromatrizz[63][288] = 9'b111110010;
assign micromatrizz[63][289] = 9'b111110011;
assign micromatrizz[63][290] = 9'b111110011;
assign micromatrizz[63][291] = 9'b111110011;
assign micromatrizz[63][292] = 9'b111110011;
assign micromatrizz[63][293] = 9'b111110111;
assign micromatrizz[63][294] = 9'b111111111;
assign micromatrizz[63][295] = 9'b111111111;
assign micromatrizz[63][296] = 9'b111111111;
assign micromatrizz[63][297] = 9'b111111111;
assign micromatrizz[63][298] = 9'b111111111;
assign micromatrizz[63][299] = 9'b111111111;
assign micromatrizz[63][300] = 9'b111111111;
assign micromatrizz[63][301] = 9'b111111111;
assign micromatrizz[63][302] = 9'b111110010;
assign micromatrizz[63][303] = 9'b111110010;
assign micromatrizz[63][304] = 9'b111110010;
assign micromatrizz[63][305] = 9'b111110011;
assign micromatrizz[63][306] = 9'b111110011;
assign micromatrizz[63][307] = 9'b111110010;
assign micromatrizz[63][308] = 9'b111110010;
assign micromatrizz[63][309] = 9'b111111111;
assign micromatrizz[63][310] = 9'b111111111;
assign micromatrizz[63][311] = 9'b111111111;
assign micromatrizz[63][312] = 9'b111111111;
assign micromatrizz[63][313] = 9'b111111111;
assign micromatrizz[63][314] = 9'b111111111;
assign micromatrizz[63][315] = 9'b111111111;
assign micromatrizz[63][316] = 9'b111110010;
assign micromatrizz[63][317] = 9'b111110010;
assign micromatrizz[63][318] = 9'b111110011;
assign micromatrizz[63][319] = 9'b111110011;
assign micromatrizz[63][320] = 9'b111110011;
assign micromatrizz[63][321] = 9'b111110011;
assign micromatrizz[63][322] = 9'b111111111;
assign micromatrizz[63][323] = 9'b111111111;
assign micromatrizz[63][324] = 9'b111111111;
assign micromatrizz[63][325] = 9'b111111111;
assign micromatrizz[63][326] = 9'b111111111;
assign micromatrizz[63][327] = 9'b111111111;
assign micromatrizz[63][328] = 9'b111111111;
assign micromatrizz[63][329] = 9'b111111111;
assign micromatrizz[63][330] = 9'b111111111;
assign micromatrizz[63][331] = 9'b111111111;
assign micromatrizz[63][332] = 9'b111111111;
assign micromatrizz[63][333] = 9'b111111111;
assign micromatrizz[63][334] = 9'b111111111;
assign micromatrizz[63][335] = 9'b111110010;
assign micromatrizz[63][336] = 9'b111110010;
assign micromatrizz[63][337] = 9'b111110011;
assign micromatrizz[63][338] = 9'b111110011;
assign micromatrizz[63][339] = 9'b111110010;
assign micromatrizz[63][340] = 9'b111110010;
assign micromatrizz[63][341] = 9'b111110011;
assign micromatrizz[63][342] = 9'b111111111;
assign micromatrizz[63][343] = 9'b111111111;
assign micromatrizz[63][344] = 9'b111111111;
assign micromatrizz[63][345] = 9'b111111111;
assign micromatrizz[63][346] = 9'b111111111;
assign micromatrizz[63][347] = 9'b111110010;
assign micromatrizz[63][348] = 9'b111110010;
assign micromatrizz[63][349] = 9'b111110010;
assign micromatrizz[63][350] = 9'b111110010;
assign micromatrizz[63][351] = 9'b111110011;
assign micromatrizz[63][352] = 9'b111110011;
assign micromatrizz[63][353] = 9'b111110011;
assign micromatrizz[63][354] = 9'b111111111;
assign micromatrizz[63][355] = 9'b111111111;
assign micromatrizz[63][356] = 9'b111111111;
assign micromatrizz[63][357] = 9'b111111111;
assign micromatrizz[63][358] = 9'b111111111;
assign micromatrizz[63][359] = 9'b111110010;
assign micromatrizz[63][360] = 9'b111110011;
assign micromatrizz[63][361] = 9'b111110010;
assign micromatrizz[63][362] = 9'b111110010;
assign micromatrizz[63][363] = 9'b111110011;
assign micromatrizz[63][364] = 9'b111110011;
assign micromatrizz[63][365] = 9'b111110010;
assign micromatrizz[63][366] = 9'b111111111;
assign micromatrizz[63][367] = 9'b111111111;
assign micromatrizz[63][368] = 9'b111111111;
assign micromatrizz[63][369] = 9'b111111111;
assign micromatrizz[63][370] = 9'b111111111;
assign micromatrizz[63][371] = 9'b111111111;
assign micromatrizz[63][372] = 9'b111110010;
assign micromatrizz[63][373] = 9'b111110010;
assign micromatrizz[63][374] = 9'b111110011;
assign micromatrizz[63][375] = 9'b111110011;
assign micromatrizz[63][376] = 9'b111110011;
assign micromatrizz[63][377] = 9'b111110011;
assign micromatrizz[63][378] = 9'b111110011;
assign micromatrizz[63][379] = 9'b111111111;
assign micromatrizz[63][380] = 9'b111111111;
assign micromatrizz[63][381] = 9'b111111111;
assign micromatrizz[63][382] = 9'b111111111;
assign micromatrizz[63][383] = 9'b111111111;
assign micromatrizz[63][384] = 9'b111110010;
assign micromatrizz[63][385] = 9'b111110010;
assign micromatrizz[63][386] = 9'b111110011;
assign micromatrizz[63][387] = 9'b111110011;
assign micromatrizz[63][388] = 9'b111110011;
assign micromatrizz[63][389] = 9'b111110011;
assign micromatrizz[63][390] = 9'b111110011;
assign micromatrizz[63][391] = 9'b111111111;
assign micromatrizz[63][392] = 9'b111111111;
assign micromatrizz[63][393] = 9'b111111111;
assign micromatrizz[63][394] = 9'b111111111;
assign micromatrizz[63][395] = 9'b111110110;
assign micromatrizz[63][396] = 9'b111110010;
assign micromatrizz[63][397] = 9'b111110010;
assign micromatrizz[63][398] = 9'b111110010;
assign micromatrizz[63][399] = 9'b111110011;
assign micromatrizz[63][400] = 9'b111110011;
assign micromatrizz[63][401] = 9'b111110011;
assign micromatrizz[63][402] = 9'b111110111;
assign micromatrizz[63][403] = 9'b111111111;
assign micromatrizz[63][404] = 9'b111111111;
assign micromatrizz[63][405] = 9'b111111111;
assign micromatrizz[63][406] = 9'b111111111;
assign micromatrizz[63][407] = 9'b111111111;
assign micromatrizz[63][408] = 9'b111111111;
assign micromatrizz[63][409] = 9'b111111111;
assign micromatrizz[63][410] = 9'b111111111;
assign micromatrizz[63][411] = 9'b111110110;
assign micromatrizz[63][412] = 9'b111110010;
assign micromatrizz[63][413] = 9'b111110010;
assign micromatrizz[63][414] = 9'b111110011;
assign micromatrizz[63][415] = 9'b111110011;
assign micromatrizz[63][416] = 9'b111110011;
assign micromatrizz[63][417] = 9'b111110111;
assign micromatrizz[63][418] = 9'b111111111;
assign micromatrizz[63][419] = 9'b111111111;
assign micromatrizz[63][420] = 9'b111111111;
assign micromatrizz[63][421] = 9'b111111111;
assign micromatrizz[63][422] = 9'b111111111;
assign micromatrizz[63][423] = 9'b111111111;
assign micromatrizz[63][424] = 9'b111111111;
assign micromatrizz[63][425] = 9'b111111111;
assign micromatrizz[63][426] = 9'b111111111;
assign micromatrizz[63][427] = 9'b111111111;
assign micromatrizz[63][428] = 9'b111111111;
assign micromatrizz[63][429] = 9'b111111111;
assign micromatrizz[63][430] = 9'b111110111;
assign micromatrizz[63][431] = 9'b111110010;
assign micromatrizz[63][432] = 9'b111110010;
assign micromatrizz[63][433] = 9'b111110010;
assign micromatrizz[63][434] = 9'b111110010;
assign micromatrizz[63][435] = 9'b111110011;
assign micromatrizz[63][436] = 9'b111110011;
assign micromatrizz[63][437] = 9'b111110011;
assign micromatrizz[63][438] = 9'b111111111;
assign micromatrizz[63][439] = 9'b111111111;
assign micromatrizz[63][440] = 9'b111111111;
assign micromatrizz[63][441] = 9'b111111111;
assign micromatrizz[63][442] = 9'b111111111;
assign micromatrizz[63][443] = 9'b111111111;
assign micromatrizz[63][444] = 9'b111111111;
assign micromatrizz[63][445] = 9'b111111111;
assign micromatrizz[63][446] = 9'b111110111;
assign micromatrizz[63][447] = 9'b111110010;
assign micromatrizz[63][448] = 9'b111110010;
assign micromatrizz[63][449] = 9'b111110010;
assign micromatrizz[63][450] = 9'b111110010;
assign micromatrizz[63][451] = 9'b111110011;
assign micromatrizz[63][452] = 9'b111110011;
assign micromatrizz[63][453] = 9'b111110011;
assign micromatrizz[63][454] = 9'b111111111;
assign micromatrizz[63][455] = 9'b111111111;
assign micromatrizz[63][456] = 9'b111111111;
assign micromatrizz[63][457] = 9'b111111111;
assign micromatrizz[63][458] = 9'b111111111;
assign micromatrizz[63][459] = 9'b111111111;
assign micromatrizz[63][460] = 9'b111111111;
assign micromatrizz[63][461] = 9'b111110111;
assign micromatrizz[63][462] = 9'b111110111;
assign micromatrizz[63][463] = 9'b111111111;
assign micromatrizz[63][464] = 9'b111111111;
assign micromatrizz[63][465] = 9'b111111111;
assign micromatrizz[63][466] = 9'b111111111;
assign micromatrizz[63][467] = 9'b111111111;
assign micromatrizz[63][468] = 9'b111110110;
assign micromatrizz[63][469] = 9'b111110010;
assign micromatrizz[63][470] = 9'b111110010;
assign micromatrizz[63][471] = 9'b111110010;
assign micromatrizz[63][472] = 9'b111110010;
assign micromatrizz[63][473] = 9'b111110011;
assign micromatrizz[63][474] = 9'b111110011;
assign micromatrizz[63][475] = 9'b111110011;
assign micromatrizz[63][476] = 9'b111110011;
assign micromatrizz[63][477] = 9'b111110011;
assign micromatrizz[63][478] = 9'b111111111;
assign micromatrizz[63][479] = 9'b111111111;
assign micromatrizz[63][480] = 9'b111111111;
assign micromatrizz[63][481] = 9'b111110010;
assign micromatrizz[63][482] = 9'b111110010;
assign micromatrizz[63][483] = 9'b111110010;
assign micromatrizz[63][484] = 9'b111110010;
assign micromatrizz[63][485] = 9'b111110011;
assign micromatrizz[63][486] = 9'b111110011;
assign micromatrizz[63][487] = 9'b111110011;
assign micromatrizz[63][488] = 9'b111110111;
assign micromatrizz[63][489] = 9'b111111111;
assign micromatrizz[63][490] = 9'b111111111;
assign micromatrizz[63][491] = 9'b111111111;
assign micromatrizz[63][492] = 9'b111111111;
assign micromatrizz[63][493] = 9'b111111111;
assign micromatrizz[63][494] = 9'b111111111;
assign micromatrizz[63][495] = 9'b111111111;
assign micromatrizz[63][496] = 9'b111111111;
assign micromatrizz[63][497] = 9'b111110010;
assign micromatrizz[63][498] = 9'b111110010;
assign micromatrizz[63][499] = 9'b111110010;
assign micromatrizz[63][500] = 9'b111110011;
assign micromatrizz[63][501] = 9'b111110011;
assign micromatrizz[63][502] = 9'b111110011;
assign micromatrizz[63][503] = 9'b111110111;
assign micromatrizz[63][504] = 9'b111111111;
assign micromatrizz[63][505] = 9'b111111111;
assign micromatrizz[63][506] = 9'b111111111;
assign micromatrizz[63][507] = 9'b111111111;
assign micromatrizz[63][508] = 9'b111111111;
assign micromatrizz[63][509] = 9'b111111111;
assign micromatrizz[63][510] = 9'b111111111;
assign micromatrizz[63][511] = 9'b111111111;
assign micromatrizz[63][512] = 9'b111111111;
assign micromatrizz[63][513] = 9'b111111111;
assign micromatrizz[63][514] = 9'b111111111;
assign micromatrizz[63][515] = 9'b111111111;
assign micromatrizz[63][516] = 9'b111110111;
assign micromatrizz[63][517] = 9'b111110011;
assign micromatrizz[63][518] = 9'b111110011;
assign micromatrizz[63][519] = 9'b111110010;
assign micromatrizz[63][520] = 9'b111110010;
assign micromatrizz[63][521] = 9'b111110010;
assign micromatrizz[63][522] = 9'b111110011;
assign micromatrizz[63][523] = 9'b111110111;
assign micromatrizz[63][524] = 9'b111111111;
assign micromatrizz[63][525] = 9'b111111111;
assign micromatrizz[63][526] = 9'b111111111;
assign micromatrizz[63][527] = 9'b111111111;
assign micromatrizz[63][528] = 9'b111111111;
assign micromatrizz[63][529] = 9'b111110010;
assign micromatrizz[63][530] = 9'b111110010;
assign micromatrizz[63][531] = 9'b111110010;
assign micromatrizz[63][532] = 9'b111110011;
assign micromatrizz[63][533] = 9'b111110011;
assign micromatrizz[63][534] = 9'b111110011;
assign micromatrizz[63][535] = 9'b111110011;
assign micromatrizz[63][536] = 9'b111111111;
assign micromatrizz[63][537] = 9'b111111111;
assign micromatrizz[63][538] = 9'b111111111;
assign micromatrizz[63][539] = 9'b111110010;
assign micromatrizz[63][540] = 9'b111110011;
assign micromatrizz[63][541] = 9'b111110011;
assign micromatrizz[63][542] = 9'b111110010;
assign micromatrizz[63][543] = 9'b111110011;
assign micromatrizz[63][544] = 9'b111110010;
assign micromatrizz[63][545] = 9'b111111111;
assign micromatrizz[63][546] = 9'b111111111;
assign micromatrizz[63][547] = 9'b111111111;
assign micromatrizz[63][548] = 9'b111111111;
assign micromatrizz[63][549] = 9'b111111111;
assign micromatrizz[63][550] = 9'b111111111;
assign micromatrizz[63][551] = 9'b111111111;
assign micromatrizz[63][552] = 9'b111111111;
assign micromatrizz[63][553] = 9'b111111111;
assign micromatrizz[63][554] = 9'b111111111;
assign micromatrizz[63][555] = 9'b111111111;
assign micromatrizz[63][556] = 9'b111111111;
assign micromatrizz[63][557] = 9'b111111111;
assign micromatrizz[63][558] = 9'b111110010;
assign micromatrizz[63][559] = 9'b111110010;
assign micromatrizz[63][560] = 9'b111110010;
assign micromatrizz[63][561] = 9'b111110010;
assign micromatrizz[63][562] = 9'b111110011;
assign micromatrizz[63][563] = 9'b111110011;
assign micromatrizz[63][564] = 9'b111110010;
assign micromatrizz[63][565] = 9'b111111111;
assign micromatrizz[63][566] = 9'b111111111;
assign micromatrizz[63][567] = 9'b111111111;
assign micromatrizz[63][568] = 9'b111110111;
assign micromatrizz[63][569] = 9'b111110010;
assign micromatrizz[63][570] = 9'b111110010;
assign micromatrizz[63][571] = 9'b111110010;
assign micromatrizz[63][572] = 9'b111110010;
assign micromatrizz[63][573] = 9'b111110011;
assign micromatrizz[63][574] = 9'b111110011;
assign micromatrizz[63][575] = 9'b111110011;
assign micromatrizz[63][576] = 9'b111111111;
assign micromatrizz[63][577] = 9'b111111111;
assign micromatrizz[63][578] = 9'b111111111;
assign micromatrizz[63][579] = 9'b111111111;
assign micromatrizz[63][580] = 9'b111111111;
assign micromatrizz[63][581] = 9'b111110010;
assign micromatrizz[63][582] = 9'b111110010;
assign micromatrizz[63][583] = 9'b111110011;
assign micromatrizz[63][584] = 9'b111110011;
assign micromatrizz[63][585] = 9'b111110011;
assign micromatrizz[63][586] = 9'b111110011;
assign micromatrizz[63][587] = 9'b111110011;
assign micromatrizz[63][588] = 9'b111111111;
assign micromatrizz[63][589] = 9'b111111111;
assign micromatrizz[63][590] = 9'b111111111;
assign micromatrizz[63][591] = 9'b111111111;
assign micromatrizz[63][592] = 9'b111110010;
assign micromatrizz[63][593] = 9'b111110010;
assign micromatrizz[63][594] = 9'b111110011;
assign micromatrizz[63][595] = 9'b111110011;
assign micromatrizz[63][596] = 9'b111110011;
assign micromatrizz[63][597] = 9'b111110011;
assign micromatrizz[63][598] = 9'b111111111;
assign micromatrizz[63][599] = 9'b111111111;
assign micromatrizz[63][600] = 9'b111111111;
assign micromatrizz[63][601] = 9'b111111111;
assign micromatrizz[63][602] = 9'b111111111;
assign micromatrizz[63][603] = 9'b111111111;
assign micromatrizz[63][604] = 9'b111111111;
assign micromatrizz[63][605] = 9'b111111111;
assign micromatrizz[63][606] = 9'b111111111;
assign micromatrizz[63][607] = 9'b111111111;
assign micromatrizz[63][608] = 9'b111111111;
assign micromatrizz[63][609] = 9'b111111111;
assign micromatrizz[63][610] = 9'b111111111;
assign micromatrizz[63][611] = 9'b111111111;
assign micromatrizz[63][612] = 9'b111111111;
assign micromatrizz[63][613] = 9'b111110111;
assign micromatrizz[63][614] = 9'b111110010;
assign micromatrizz[63][615] = 9'b111110011;
assign micromatrizz[63][616] = 9'b111110011;
assign micromatrizz[63][617] = 9'b111110011;
assign micromatrizz[63][618] = 9'b111110010;
assign micromatrizz[63][619] = 9'b111110011;
assign micromatrizz[63][620] = 9'b111110011;
assign micromatrizz[63][621] = 9'b111110011;
assign micromatrizz[63][622] = 9'b111110111;
assign micromatrizz[63][623] = 9'b111111111;
assign micromatrizz[63][624] = 9'b111111111;
assign micromatrizz[63][625] = 9'b111111111;
assign micromatrizz[63][626] = 9'b111111111;
assign micromatrizz[63][627] = 9'b111111111;
assign micromatrizz[63][628] = 9'b111111111;
assign micromatrizz[63][629] = 9'b111111111;
assign micromatrizz[63][630] = 9'b111111111;
assign micromatrizz[63][631] = 9'b111111111;
assign micromatrizz[63][632] = 9'b111111111;
assign micromatrizz[63][633] = 9'b111111111;
assign micromatrizz[63][634] = 9'b111111111;
assign micromatrizz[63][635] = 9'b111111111;
assign micromatrizz[63][636] = 9'b111111111;
assign micromatrizz[63][637] = 9'b111111111;
assign micromatrizz[63][638] = 9'b111111111;
assign micromatrizz[63][639] = 9'b111111111;
assign micromatrizz[64][0] = 9'b111111111;
assign micromatrizz[64][1] = 9'b111111111;
assign micromatrizz[64][2] = 9'b111111111;
assign micromatrizz[64][3] = 9'b111111111;
assign micromatrizz[64][4] = 9'b111111111;
assign micromatrizz[64][5] = 9'b111111111;
assign micromatrizz[64][6] = 9'b111111111;
assign micromatrizz[64][7] = 9'b111111111;
assign micromatrizz[64][8] = 9'b111111111;
assign micromatrizz[64][9] = 9'b111111111;
assign micromatrizz[64][10] = 9'b111111111;
assign micromatrizz[64][11] = 9'b111111111;
assign micromatrizz[64][12] = 9'b111110010;
assign micromatrizz[64][13] = 9'b111110010;
assign micromatrizz[64][14] = 9'b111110011;
assign micromatrizz[64][15] = 9'b111110011;
assign micromatrizz[64][16] = 9'b111110011;
assign micromatrizz[64][17] = 9'b111110011;
assign micromatrizz[64][18] = 9'b111110011;
assign micromatrizz[64][19] = 9'b111110011;
assign micromatrizz[64][20] = 9'b111110011;
assign micromatrizz[64][21] = 9'b111111111;
assign micromatrizz[64][22] = 9'b111111111;
assign micromatrizz[64][23] = 9'b111111111;
assign micromatrizz[64][24] = 9'b111110010;
assign micromatrizz[64][25] = 9'b111110010;
assign micromatrizz[64][26] = 9'b111110010;
assign micromatrizz[64][27] = 9'b111110011;
assign micromatrizz[64][28] = 9'b111110011;
assign micromatrizz[64][29] = 9'b111110011;
assign micromatrizz[64][30] = 9'b111110011;
assign micromatrizz[64][31] = 9'b111111111;
assign micromatrizz[64][32] = 9'b111111111;
assign micromatrizz[64][33] = 9'b111111111;
assign micromatrizz[64][34] = 9'b111111111;
assign micromatrizz[64][35] = 9'b111110111;
assign micromatrizz[64][36] = 9'b111110010;
assign micromatrizz[64][37] = 9'b111110011;
assign micromatrizz[64][38] = 9'b111110011;
assign micromatrizz[64][39] = 9'b111110011;
assign micromatrizz[64][40] = 9'b111110011;
assign micromatrizz[64][41] = 9'b111110011;
assign micromatrizz[64][42] = 9'b111110011;
assign micromatrizz[64][43] = 9'b111111111;
assign micromatrizz[64][44] = 9'b111111111;
assign micromatrizz[64][45] = 9'b111111111;
assign micromatrizz[64][46] = 9'b111111111;
assign micromatrizz[64][47] = 9'b111110010;
assign micromatrizz[64][48] = 9'b111110010;
assign micromatrizz[64][49] = 9'b111110010;
assign micromatrizz[64][50] = 9'b111110011;
assign micromatrizz[64][51] = 9'b111110011;
assign micromatrizz[64][52] = 9'b111110011;
assign micromatrizz[64][53] = 9'b111110011;
assign micromatrizz[64][54] = 9'b111110111;
assign micromatrizz[64][55] = 9'b111111111;
assign micromatrizz[64][56] = 9'b111111111;
assign micromatrizz[64][57] = 9'b111111111;
assign micromatrizz[64][58] = 9'b111111111;
assign micromatrizz[64][59] = 9'b111110010;
assign micromatrizz[64][60] = 9'b111110010;
assign micromatrizz[64][61] = 9'b111110010;
assign micromatrizz[64][62] = 9'b111110011;
assign micromatrizz[64][63] = 9'b111110011;
assign micromatrizz[64][64] = 9'b111110011;
assign micromatrizz[64][65] = 9'b111110111;
assign micromatrizz[64][66] = 9'b111111111;
assign micromatrizz[64][67] = 9'b111111111;
assign micromatrizz[64][68] = 9'b111111111;
assign micromatrizz[64][69] = 9'b111110010;
assign micromatrizz[64][70] = 9'b111110010;
assign micromatrizz[64][71] = 9'b111110010;
assign micromatrizz[64][72] = 9'b111110010;
assign micromatrizz[64][73] = 9'b111110010;
assign micromatrizz[64][74] = 9'b111110011;
assign micromatrizz[64][75] = 9'b111111111;
assign micromatrizz[64][76] = 9'b111111111;
assign micromatrizz[64][77] = 9'b111111111;
assign micromatrizz[64][78] = 9'b111111111;
assign micromatrizz[64][79] = 9'b111111111;
assign micromatrizz[64][80] = 9'b111111111;
assign micromatrizz[64][81] = 9'b111111111;
assign micromatrizz[64][82] = 9'b111111111;
assign micromatrizz[64][83] = 9'b111111111;
assign micromatrizz[64][84] = 9'b111111111;
assign micromatrizz[64][85] = 9'b111111111;
assign micromatrizz[64][86] = 9'b111111111;
assign micromatrizz[64][87] = 9'b111111111;
assign micromatrizz[64][88] = 9'b111110110;
assign micromatrizz[64][89] = 9'b111110010;
assign micromatrizz[64][90] = 9'b111110010;
assign micromatrizz[64][91] = 9'b111110011;
assign micromatrizz[64][92] = 9'b111110011;
assign micromatrizz[64][93] = 9'b111110011;
assign micromatrizz[64][94] = 9'b111110011;
assign micromatrizz[64][95] = 9'b111110111;
assign micromatrizz[64][96] = 9'b111111111;
assign micromatrizz[64][97] = 9'b111111111;
assign micromatrizz[64][98] = 9'b111111111;
assign micromatrizz[64][99] = 9'b111111111;
assign micromatrizz[64][100] = 9'b111111111;
assign micromatrizz[64][101] = 9'b111111111;
assign micromatrizz[64][102] = 9'b111111111;
assign micromatrizz[64][103] = 9'b111111111;
assign micromatrizz[64][104] = 9'b111111111;
assign micromatrizz[64][105] = 9'b111111111;
assign micromatrizz[64][106] = 9'b111111111;
assign micromatrizz[64][107] = 9'b111111111;
assign micromatrizz[64][108] = 9'b111110010;
assign micromatrizz[64][109] = 9'b111110010;
assign micromatrizz[64][110] = 9'b111110010;
assign micromatrizz[64][111] = 9'b111110011;
assign micromatrizz[64][112] = 9'b111110011;
assign micromatrizz[64][113] = 9'b111110011;
assign micromatrizz[64][114] = 9'b111110011;
assign micromatrizz[64][115] = 9'b111110011;
assign micromatrizz[64][116] = 9'b111110011;
assign micromatrizz[64][117] = 9'b111111111;
assign micromatrizz[64][118] = 9'b111111111;
assign micromatrizz[64][119] = 9'b111110111;
assign micromatrizz[64][120] = 9'b111110010;
assign micromatrizz[64][121] = 9'b111110010;
assign micromatrizz[64][122] = 9'b111110010;
assign micromatrizz[64][123] = 9'b111110010;
assign micromatrizz[64][124] = 9'b111110011;
assign micromatrizz[64][125] = 9'b111110011;
assign micromatrizz[64][126] = 9'b111110011;
assign micromatrizz[64][127] = 9'b111111111;
assign micromatrizz[64][128] = 9'b111111111;
assign micromatrizz[64][129] = 9'b111111111;
assign micromatrizz[64][130] = 9'b111111111;
assign micromatrizz[64][131] = 9'b111111111;
assign micromatrizz[64][132] = 9'b111111111;
assign micromatrizz[64][133] = 9'b111111111;
assign micromatrizz[64][134] = 9'b111110110;
assign micromatrizz[64][135] = 9'b111111111;
assign micromatrizz[64][136] = 9'b111111111;
assign micromatrizz[64][137] = 9'b111111111;
assign micromatrizz[64][138] = 9'b111110111;
assign micromatrizz[64][139] = 9'b111110010;
assign micromatrizz[64][140] = 9'b111110010;
assign micromatrizz[64][141] = 9'b111110010;
assign micromatrizz[64][142] = 9'b111110010;
assign micromatrizz[64][143] = 9'b111110011;
assign micromatrizz[64][144] = 9'b111110011;
assign micromatrizz[64][145] = 9'b111110011;
assign micromatrizz[64][146] = 9'b111111111;
assign micromatrizz[64][147] = 9'b111111111;
assign micromatrizz[64][148] = 9'b111111111;
assign micromatrizz[64][149] = 9'b111111111;
assign micromatrizz[64][150] = 9'b111110111;
assign micromatrizz[64][151] = 9'b111110010;
assign micromatrizz[64][152] = 9'b111110010;
assign micromatrizz[64][153] = 9'b111110011;
assign micromatrizz[64][154] = 9'b111110011;
assign micromatrizz[64][155] = 9'b111110011;
assign micromatrizz[64][156] = 9'b111110011;
assign micromatrizz[64][157] = 9'b111110111;
assign micromatrizz[64][158] = 9'b111111111;
assign micromatrizz[64][159] = 9'b111111111;
assign micromatrizz[64][160] = 9'b111111111;
assign micromatrizz[64][161] = 9'b111110010;
assign micromatrizz[64][162] = 9'b111110010;
assign micromatrizz[64][163] = 9'b111110010;
assign micromatrizz[64][164] = 9'b111110011;
assign micromatrizz[64][165] = 9'b111110011;
assign micromatrizz[64][166] = 9'b111110011;
assign micromatrizz[64][167] = 9'b111110010;
assign micromatrizz[64][168] = 9'b111111111;
assign micromatrizz[64][169] = 9'b111111111;
assign micromatrizz[64][170] = 9'b111111111;
assign micromatrizz[64][171] = 9'b111111111;
assign micromatrizz[64][172] = 9'b111110010;
assign micromatrizz[64][173] = 9'b111110011;
assign micromatrizz[64][174] = 9'b111110011;
assign micromatrizz[64][175] = 9'b111110011;
assign micromatrizz[64][176] = 9'b111110011;
assign micromatrizz[64][177] = 9'b111110011;
assign micromatrizz[64][178] = 9'b111110010;
assign micromatrizz[64][179] = 9'b111110111;
assign micromatrizz[64][180] = 9'b111111111;
assign micromatrizz[64][181] = 9'b111111111;
assign micromatrizz[64][182] = 9'b111111111;
assign micromatrizz[64][183] = 9'b111110010;
assign micromatrizz[64][184] = 9'b111110011;
assign micromatrizz[64][185] = 9'b111110011;
assign micromatrizz[64][186] = 9'b111110010;
assign micromatrizz[64][187] = 9'b111110010;
assign micromatrizz[64][188] = 9'b111110011;
assign micromatrizz[64][189] = 9'b111110011;
assign micromatrizz[64][190] = 9'b111111111;
assign micromatrizz[64][191] = 9'b111111111;
assign micromatrizz[64][192] = 9'b111111111;
assign micromatrizz[64][193] = 9'b111111111;
assign micromatrizz[64][194] = 9'b111111111;
assign micromatrizz[64][195] = 9'b111110110;
assign micromatrizz[64][196] = 9'b111110010;
assign micromatrizz[64][197] = 9'b111110011;
assign micromatrizz[64][198] = 9'b111110011;
assign micromatrizz[64][199] = 9'b111110010;
assign micromatrizz[64][200] = 9'b111110010;
assign micromatrizz[64][201] = 9'b111110011;
assign micromatrizz[64][202] = 9'b111110111;
assign micromatrizz[64][203] = 9'b111111111;
assign micromatrizz[64][204] = 9'b111111111;
assign micromatrizz[64][205] = 9'b111111111;
assign micromatrizz[64][206] = 9'b111110110;
assign micromatrizz[64][207] = 9'b111110010;
assign micromatrizz[64][208] = 9'b111110010;
assign micromatrizz[64][209] = 9'b111110010;
assign micromatrizz[64][210] = 9'b111110010;
assign micromatrizz[64][211] = 9'b111110011;
assign micromatrizz[64][212] = 9'b111110011;
assign micromatrizz[64][213] = 9'b111110111;
assign micromatrizz[64][214] = 9'b111111111;
assign micromatrizz[64][215] = 9'b111111111;
assign micromatrizz[64][216] = 9'b111111111;
assign micromatrizz[64][217] = 9'b111111111;
assign micromatrizz[64][218] = 9'b111111111;
assign micromatrizz[64][219] = 9'b111111111;
assign micromatrizz[64][220] = 9'b111111111;
assign micromatrizz[64][221] = 9'b111110111;
assign micromatrizz[64][222] = 9'b111111111;
assign micromatrizz[64][223] = 9'b111111111;
assign micromatrizz[64][224] = 9'b111111111;
assign micromatrizz[64][225] = 9'b111110010;
assign micromatrizz[64][226] = 9'b111110010;
assign micromatrizz[64][227] = 9'b111110010;
assign micromatrizz[64][228] = 9'b111110010;
assign micromatrizz[64][229] = 9'b111110011;
assign micromatrizz[64][230] = 9'b111110011;
assign micromatrizz[64][231] = 9'b111110011;
assign micromatrizz[64][232] = 9'b111110111;
assign micromatrizz[64][233] = 9'b111111111;
assign micromatrizz[64][234] = 9'b111111111;
assign micromatrizz[64][235] = 9'b111111111;
assign micromatrizz[64][236] = 9'b111111111;
assign micromatrizz[64][237] = 9'b111111111;
assign micromatrizz[64][238] = 9'b111111111;
assign micromatrizz[64][239] = 9'b111111111;
assign micromatrizz[64][240] = 9'b111111111;
assign micromatrizz[64][241] = 9'b111110111;
assign micromatrizz[64][242] = 9'b111110010;
assign micromatrizz[64][243] = 9'b111110010;
assign micromatrizz[64][244] = 9'b111110010;
assign micromatrizz[64][245] = 9'b111110011;
assign micromatrizz[64][246] = 9'b111110010;
assign micromatrizz[64][247] = 9'b111110111;
assign micromatrizz[64][248] = 9'b111111111;
assign micromatrizz[64][249] = 9'b111111111;
assign micromatrizz[64][250] = 9'b111111111;
assign micromatrizz[64][251] = 9'b111111111;
assign micromatrizz[64][252] = 9'b111111111;
assign micromatrizz[64][253] = 9'b111111111;
assign micromatrizz[64][254] = 9'b111111111;
assign micromatrizz[64][255] = 9'b111111111;
assign micromatrizz[64][256] = 9'b111111111;
assign micromatrizz[64][257] = 9'b111111111;
assign micromatrizz[64][258] = 9'b111111111;
assign micromatrizz[64][259] = 9'b111111111;
assign micromatrizz[64][260] = 9'b111111111;
assign micromatrizz[64][261] = 9'b111111111;
assign micromatrizz[64][262] = 9'b111111111;
assign micromatrizz[64][263] = 9'b111111111;
assign micromatrizz[64][264] = 9'b111110010;
assign micromatrizz[64][265] = 9'b111110010;
assign micromatrizz[64][266] = 9'b111110011;
assign micromatrizz[64][267] = 9'b111110011;
assign micromatrizz[64][268] = 9'b111110011;
assign micromatrizz[64][269] = 9'b111110011;
assign micromatrizz[64][270] = 9'b111110011;
assign micromatrizz[64][271] = 9'b111110010;
assign micromatrizz[64][272] = 9'b111110111;
assign micromatrizz[64][273] = 9'b111111111;
assign micromatrizz[64][274] = 9'b111110111;
assign micromatrizz[64][275] = 9'b111110010;
assign micromatrizz[64][276] = 9'b111110010;
assign micromatrizz[64][277] = 9'b111110010;
assign micromatrizz[64][278] = 9'b111110011;
assign micromatrizz[64][279] = 9'b111110011;
assign micromatrizz[64][280] = 9'b111110011;
assign micromatrizz[64][281] = 9'b111110011;
assign micromatrizz[64][282] = 9'b111111111;
assign micromatrizz[64][283] = 9'b111111111;
assign micromatrizz[64][284] = 9'b111111111;
assign micromatrizz[64][285] = 9'b111111111;
assign micromatrizz[64][286] = 9'b111110010;
assign micromatrizz[64][287] = 9'b111110011;
assign micromatrizz[64][288] = 9'b111110011;
assign micromatrizz[64][289] = 9'b111110011;
assign micromatrizz[64][290] = 9'b111110011;
assign micromatrizz[64][291] = 9'b111110011;
assign micromatrizz[64][292] = 9'b111110011;
assign micromatrizz[64][293] = 9'b111110111;
assign micromatrizz[64][294] = 9'b111111111;
assign micromatrizz[64][295] = 9'b111111111;
assign micromatrizz[64][296] = 9'b111111111;
assign micromatrizz[64][297] = 9'b111111111;
assign micromatrizz[64][298] = 9'b111111111;
assign micromatrizz[64][299] = 9'b111111111;
assign micromatrizz[64][300] = 9'b111111111;
assign micromatrizz[64][301] = 9'b111111111;
assign micromatrizz[64][302] = 9'b111110111;
assign micromatrizz[64][303] = 9'b111110010;
assign micromatrizz[64][304] = 9'b111110011;
assign micromatrizz[64][305] = 9'b111110011;
assign micromatrizz[64][306] = 9'b111110011;
assign micromatrizz[64][307] = 9'b111110010;
assign micromatrizz[64][308] = 9'b111110111;
assign micromatrizz[64][309] = 9'b111111111;
assign micromatrizz[64][310] = 9'b111111111;
assign micromatrizz[64][311] = 9'b111111111;
assign micromatrizz[64][312] = 9'b111111111;
assign micromatrizz[64][313] = 9'b111111111;
assign micromatrizz[64][314] = 9'b111111111;
assign micromatrizz[64][315] = 9'b111111111;
assign micromatrizz[64][316] = 9'b111110010;
assign micromatrizz[64][317] = 9'b111110011;
assign micromatrizz[64][318] = 9'b111110010;
assign micromatrizz[64][319] = 9'b111110011;
assign micromatrizz[64][320] = 9'b111110011;
assign micromatrizz[64][321] = 9'b111110011;
assign micromatrizz[64][322] = 9'b111111111;
assign micromatrizz[64][323] = 9'b111111111;
assign micromatrizz[64][324] = 9'b111111111;
assign micromatrizz[64][325] = 9'b111111111;
assign micromatrizz[64][326] = 9'b111111111;
assign micromatrizz[64][327] = 9'b111111111;
assign micromatrizz[64][328] = 9'b111111111;
assign micromatrizz[64][329] = 9'b111111111;
assign micromatrizz[64][330] = 9'b111111111;
assign micromatrizz[64][331] = 9'b111111111;
assign micromatrizz[64][332] = 9'b111111111;
assign micromatrizz[64][333] = 9'b111111111;
assign micromatrizz[64][334] = 9'b111111111;
assign micromatrizz[64][335] = 9'b111110010;
assign micromatrizz[64][336] = 9'b111110011;
assign micromatrizz[64][337] = 9'b111110011;
assign micromatrizz[64][338] = 9'b111110011;
assign micromatrizz[64][339] = 9'b111110010;
assign micromatrizz[64][340] = 9'b111110010;
assign micromatrizz[64][341] = 9'b111110011;
assign micromatrizz[64][342] = 9'b111111111;
assign micromatrizz[64][343] = 9'b111111111;
assign micromatrizz[64][344] = 9'b111111111;
assign micromatrizz[64][345] = 9'b111111111;
assign micromatrizz[64][346] = 9'b111111111;
assign micromatrizz[64][347] = 9'b111110010;
assign micromatrizz[64][348] = 9'b111110010;
assign micromatrizz[64][349] = 9'b111110010;
assign micromatrizz[64][350] = 9'b111110010;
assign micromatrizz[64][351] = 9'b111110011;
assign micromatrizz[64][352] = 9'b111110011;
assign micromatrizz[64][353] = 9'b111110011;
assign micromatrizz[64][354] = 9'b111111111;
assign micromatrizz[64][355] = 9'b111111111;
assign micromatrizz[64][356] = 9'b111111111;
assign micromatrizz[64][357] = 9'b111111111;
assign micromatrizz[64][358] = 9'b111111111;
assign micromatrizz[64][359] = 9'b111110010;
assign micromatrizz[64][360] = 9'b111110011;
assign micromatrizz[64][361] = 9'b111110010;
assign micromatrizz[64][362] = 9'b111110010;
assign micromatrizz[64][363] = 9'b111110011;
assign micromatrizz[64][364] = 9'b111110011;
assign micromatrizz[64][365] = 9'b111110010;
assign micromatrizz[64][366] = 9'b111111111;
assign micromatrizz[64][367] = 9'b111111111;
assign micromatrizz[64][368] = 9'b111111111;
assign micromatrizz[64][369] = 9'b111111111;
assign micromatrizz[64][370] = 9'b111111111;
assign micromatrizz[64][371] = 9'b111110111;
assign micromatrizz[64][372] = 9'b111110010;
assign micromatrizz[64][373] = 9'b111110011;
assign micromatrizz[64][374] = 9'b111110011;
assign micromatrizz[64][375] = 9'b111110011;
assign micromatrizz[64][376] = 9'b111110011;
assign micromatrizz[64][377] = 9'b111110011;
assign micromatrizz[64][378] = 9'b111110011;
assign micromatrizz[64][379] = 9'b111111111;
assign micromatrizz[64][380] = 9'b111111111;
assign micromatrizz[64][381] = 9'b111111111;
assign micromatrizz[64][382] = 9'b111111111;
assign micromatrizz[64][383] = 9'b111111111;
assign micromatrizz[64][384] = 9'b111110010;
assign micromatrizz[64][385] = 9'b111110010;
assign micromatrizz[64][386] = 9'b111110011;
assign micromatrizz[64][387] = 9'b111110011;
assign micromatrizz[64][388] = 9'b111110011;
assign micromatrizz[64][389] = 9'b111110011;
assign micromatrizz[64][390] = 9'b111110011;
assign micromatrizz[64][391] = 9'b111111111;
assign micromatrizz[64][392] = 9'b111111111;
assign micromatrizz[64][393] = 9'b111111111;
assign micromatrizz[64][394] = 9'b111111111;
assign micromatrizz[64][395] = 9'b111110010;
assign micromatrizz[64][396] = 9'b111110010;
assign micromatrizz[64][397] = 9'b111110010;
assign micromatrizz[64][398] = 9'b111110010;
assign micromatrizz[64][399] = 9'b111110011;
assign micromatrizz[64][400] = 9'b111110011;
assign micromatrizz[64][401] = 9'b111110011;
assign micromatrizz[64][402] = 9'b111110111;
assign micromatrizz[64][403] = 9'b111111111;
assign micromatrizz[64][404] = 9'b111111111;
assign micromatrizz[64][405] = 9'b111111111;
assign micromatrizz[64][406] = 9'b111111111;
assign micromatrizz[64][407] = 9'b111111111;
assign micromatrizz[64][408] = 9'b111111111;
assign micromatrizz[64][409] = 9'b111111111;
assign micromatrizz[64][410] = 9'b111111111;
assign micromatrizz[64][411] = 9'b111110111;
assign micromatrizz[64][412] = 9'b111110010;
assign micromatrizz[64][413] = 9'b111110011;
assign micromatrizz[64][414] = 9'b111110011;
assign micromatrizz[64][415] = 9'b111110010;
assign micromatrizz[64][416] = 9'b111110011;
assign micromatrizz[64][417] = 9'b111110111;
assign micromatrizz[64][418] = 9'b111111111;
assign micromatrizz[64][419] = 9'b111111111;
assign micromatrizz[64][420] = 9'b111111111;
assign micromatrizz[64][421] = 9'b111111111;
assign micromatrizz[64][422] = 9'b111111111;
assign micromatrizz[64][423] = 9'b111111111;
assign micromatrizz[64][424] = 9'b111111111;
assign micromatrizz[64][425] = 9'b111111111;
assign micromatrizz[64][426] = 9'b111111111;
assign micromatrizz[64][427] = 9'b111111111;
assign micromatrizz[64][428] = 9'b111111111;
assign micromatrizz[64][429] = 9'b111111111;
assign micromatrizz[64][430] = 9'b111110111;
assign micromatrizz[64][431] = 9'b111110010;
assign micromatrizz[64][432] = 9'b111110010;
assign micromatrizz[64][433] = 9'b111110010;
assign micromatrizz[64][434] = 9'b111110010;
assign micromatrizz[64][435] = 9'b111110011;
assign micromatrizz[64][436] = 9'b111110011;
assign micromatrizz[64][437] = 9'b111110011;
assign micromatrizz[64][438] = 9'b111111111;
assign micromatrizz[64][439] = 9'b111111111;
assign micromatrizz[64][440] = 9'b111111111;
assign micromatrizz[64][441] = 9'b111111111;
assign micromatrizz[64][442] = 9'b111111111;
assign micromatrizz[64][443] = 9'b111111111;
assign micromatrizz[64][444] = 9'b111111111;
assign micromatrizz[64][445] = 9'b111111111;
assign micromatrizz[64][446] = 9'b111111111;
assign micromatrizz[64][447] = 9'b111110010;
assign micromatrizz[64][448] = 9'b111110010;
assign micromatrizz[64][449] = 9'b111110010;
assign micromatrizz[64][450] = 9'b111110010;
assign micromatrizz[64][451] = 9'b111110011;
assign micromatrizz[64][452] = 9'b111110011;
assign micromatrizz[64][453] = 9'b111110011;
assign micromatrizz[64][454] = 9'b111111111;
assign micromatrizz[64][455] = 9'b111111111;
assign micromatrizz[64][456] = 9'b111111111;
assign micromatrizz[64][457] = 9'b111111111;
assign micromatrizz[64][458] = 9'b111111111;
assign micromatrizz[64][459] = 9'b111111111;
assign micromatrizz[64][460] = 9'b111111111;
assign micromatrizz[64][461] = 9'b111110111;
assign micromatrizz[64][462] = 9'b111111111;
assign micromatrizz[64][463] = 9'b111111111;
assign micromatrizz[64][464] = 9'b111111111;
assign micromatrizz[64][465] = 9'b111111111;
assign micromatrizz[64][466] = 9'b111111111;
assign micromatrizz[64][467] = 9'b111111111;
assign micromatrizz[64][468] = 9'b111111111;
assign micromatrizz[64][469] = 9'b111110110;
assign micromatrizz[64][470] = 9'b111110010;
assign micromatrizz[64][471] = 9'b111110011;
assign micromatrizz[64][472] = 9'b111110011;
assign micromatrizz[64][473] = 9'b111110010;
assign micromatrizz[64][474] = 9'b111110011;
assign micromatrizz[64][475] = 9'b111110011;
assign micromatrizz[64][476] = 9'b111110011;
assign micromatrizz[64][477] = 9'b111110011;
assign micromatrizz[64][478] = 9'b111111111;
assign micromatrizz[64][479] = 9'b111111111;
assign micromatrizz[64][480] = 9'b111111111;
assign micromatrizz[64][481] = 9'b111110010;
assign micromatrizz[64][482] = 9'b111110010;
assign micromatrizz[64][483] = 9'b111110010;
assign micromatrizz[64][484] = 9'b111110010;
assign micromatrizz[64][485] = 9'b111110011;
assign micromatrizz[64][486] = 9'b111110011;
assign micromatrizz[64][487] = 9'b111110011;
assign micromatrizz[64][488] = 9'b111110111;
assign micromatrizz[64][489] = 9'b111111111;
assign micromatrizz[64][490] = 9'b111111111;
assign micromatrizz[64][491] = 9'b111111111;
assign micromatrizz[64][492] = 9'b111111111;
assign micromatrizz[64][493] = 9'b111111111;
assign micromatrizz[64][494] = 9'b111111111;
assign micromatrizz[64][495] = 9'b111111111;
assign micromatrizz[64][496] = 9'b111111111;
assign micromatrizz[64][497] = 9'b111110111;
assign micromatrizz[64][498] = 9'b111110010;
assign micromatrizz[64][499] = 9'b111110010;
assign micromatrizz[64][500] = 9'b111110011;
assign micromatrizz[64][501] = 9'b111110010;
assign micromatrizz[64][502] = 9'b111110010;
assign micromatrizz[64][503] = 9'b111110111;
assign micromatrizz[64][504] = 9'b111111111;
assign micromatrizz[64][505] = 9'b111111111;
assign micromatrizz[64][506] = 9'b111111111;
assign micromatrizz[64][507] = 9'b111111111;
assign micromatrizz[64][508] = 9'b111111111;
assign micromatrizz[64][509] = 9'b111111111;
assign micromatrizz[64][510] = 9'b111111111;
assign micromatrizz[64][511] = 9'b111111111;
assign micromatrizz[64][512] = 9'b111111111;
assign micromatrizz[64][513] = 9'b111111111;
assign micromatrizz[64][514] = 9'b111111111;
assign micromatrizz[64][515] = 9'b111111111;
assign micromatrizz[64][516] = 9'b111110111;
assign micromatrizz[64][517] = 9'b111110010;
assign micromatrizz[64][518] = 9'b111110011;
assign micromatrizz[64][519] = 9'b111110011;
assign micromatrizz[64][520] = 9'b111110010;
assign micromatrizz[64][521] = 9'b111110010;
assign micromatrizz[64][522] = 9'b111110011;
assign micromatrizz[64][523] = 9'b111110111;
assign micromatrizz[64][524] = 9'b111111111;
assign micromatrizz[64][525] = 9'b111111111;
assign micromatrizz[64][526] = 9'b111111111;
assign micromatrizz[64][527] = 9'b111111111;
assign micromatrizz[64][528] = 9'b111111111;
assign micromatrizz[64][529] = 9'b111110010;
assign micromatrizz[64][530] = 9'b111110010;
assign micromatrizz[64][531] = 9'b111110010;
assign micromatrizz[64][532] = 9'b111110011;
assign micromatrizz[64][533] = 9'b111110011;
assign micromatrizz[64][534] = 9'b111110011;
assign micromatrizz[64][535] = 9'b111110011;
assign micromatrizz[64][536] = 9'b111111111;
assign micromatrizz[64][537] = 9'b111111111;
assign micromatrizz[64][538] = 9'b111111111;
assign micromatrizz[64][539] = 9'b111110010;
assign micromatrizz[64][540] = 9'b111110010;
assign micromatrizz[64][541] = 9'b111110011;
assign micromatrizz[64][542] = 9'b111110010;
assign micromatrizz[64][543] = 9'b111110011;
assign micromatrizz[64][544] = 9'b111110010;
assign micromatrizz[64][545] = 9'b111111111;
assign micromatrizz[64][546] = 9'b111111111;
assign micromatrizz[64][547] = 9'b111111111;
assign micromatrizz[64][548] = 9'b111111111;
assign micromatrizz[64][549] = 9'b111111111;
assign micromatrizz[64][550] = 9'b111111111;
assign micromatrizz[64][551] = 9'b111111111;
assign micromatrizz[64][552] = 9'b111111111;
assign micromatrizz[64][553] = 9'b111111111;
assign micromatrizz[64][554] = 9'b111111111;
assign micromatrizz[64][555] = 9'b111111111;
assign micromatrizz[64][556] = 9'b111111111;
assign micromatrizz[64][557] = 9'b111111111;
assign micromatrizz[64][558] = 9'b111110010;
assign micromatrizz[64][559] = 9'b111110010;
assign micromatrizz[64][560] = 9'b111110010;
assign micromatrizz[64][561] = 9'b111110010;
assign micromatrizz[64][562] = 9'b111110011;
assign micromatrizz[64][563] = 9'b111110011;
assign micromatrizz[64][564] = 9'b111110010;
assign micromatrizz[64][565] = 9'b111111111;
assign micromatrizz[64][566] = 9'b111111111;
assign micromatrizz[64][567] = 9'b111111111;
assign micromatrizz[64][568] = 9'b111111111;
assign micromatrizz[64][569] = 9'b111110010;
assign micromatrizz[64][570] = 9'b111110010;
assign micromatrizz[64][571] = 9'b111110010;
assign micromatrizz[64][572] = 9'b111110010;
assign micromatrizz[64][573] = 9'b111110011;
assign micromatrizz[64][574] = 9'b111110011;
assign micromatrizz[64][575] = 9'b111110011;
assign micromatrizz[64][576] = 9'b111111111;
assign micromatrizz[64][577] = 9'b111111111;
assign micromatrizz[64][578] = 9'b111111111;
assign micromatrizz[64][579] = 9'b111111111;
assign micromatrizz[64][580] = 9'b111111111;
assign micromatrizz[64][581] = 9'b111110010;
assign micromatrizz[64][582] = 9'b111110011;
assign micromatrizz[64][583] = 9'b111110011;
assign micromatrizz[64][584] = 9'b111110011;
assign micromatrizz[64][585] = 9'b111110011;
assign micromatrizz[64][586] = 9'b111110011;
assign micromatrizz[64][587] = 9'b111110011;
assign micromatrizz[64][588] = 9'b111111111;
assign micromatrizz[64][589] = 9'b111111111;
assign micromatrizz[64][590] = 9'b111111111;
assign micromatrizz[64][591] = 9'b111111111;
assign micromatrizz[64][592] = 9'b111110010;
assign micromatrizz[64][593] = 9'b111110011;
assign micromatrizz[64][594] = 9'b111110010;
assign micromatrizz[64][595] = 9'b111110011;
assign micromatrizz[64][596] = 9'b111110011;
assign micromatrizz[64][597] = 9'b111110010;
assign micromatrizz[64][598] = 9'b111111111;
assign micromatrizz[64][599] = 9'b111111111;
assign micromatrizz[64][600] = 9'b111111111;
assign micromatrizz[64][601] = 9'b111111111;
assign micromatrizz[64][602] = 9'b111111111;
assign micromatrizz[64][603] = 9'b111111111;
assign micromatrizz[64][604] = 9'b111111111;
assign micromatrizz[64][605] = 9'b111111111;
assign micromatrizz[64][606] = 9'b111111111;
assign micromatrizz[64][607] = 9'b111111111;
assign micromatrizz[64][608] = 9'b111111111;
assign micromatrizz[64][609] = 9'b111111111;
assign micromatrizz[64][610] = 9'b111111111;
assign micromatrizz[64][611] = 9'b111111111;
assign micromatrizz[64][612] = 9'b111111111;
assign micromatrizz[64][613] = 9'b111111111;
assign micromatrizz[64][614] = 9'b111110111;
assign micromatrizz[64][615] = 9'b111110010;
assign micromatrizz[64][616] = 9'b111110010;
assign micromatrizz[64][617] = 9'b111110011;
assign micromatrizz[64][618] = 9'b111110011;
assign micromatrizz[64][619] = 9'b111110011;
assign micromatrizz[64][620] = 9'b111110011;
assign micromatrizz[64][621] = 9'b111110011;
assign micromatrizz[64][622] = 9'b111110011;
assign micromatrizz[64][623] = 9'b111111111;
assign micromatrizz[64][624] = 9'b111111111;
assign micromatrizz[64][625] = 9'b111111111;
assign micromatrizz[64][626] = 9'b111111111;
assign micromatrizz[64][627] = 9'b111111111;
assign micromatrizz[64][628] = 9'b111111111;
assign micromatrizz[64][629] = 9'b111111111;
assign micromatrizz[64][630] = 9'b111111111;
assign micromatrizz[64][631] = 9'b111111111;
assign micromatrizz[64][632] = 9'b111111111;
assign micromatrizz[64][633] = 9'b111111111;
assign micromatrizz[64][634] = 9'b111111111;
assign micromatrizz[64][635] = 9'b111111111;
assign micromatrizz[64][636] = 9'b111111111;
assign micromatrizz[64][637] = 9'b111111111;
assign micromatrizz[64][638] = 9'b111111111;
assign micromatrizz[64][639] = 9'b111111111;
assign micromatrizz[65][0] = 9'b111111111;
assign micromatrizz[65][1] = 9'b111111111;
assign micromatrizz[65][2] = 9'b111111111;
assign micromatrizz[65][3] = 9'b111111111;
assign micromatrizz[65][4] = 9'b111111111;
assign micromatrizz[65][5] = 9'b111111111;
assign micromatrizz[65][6] = 9'b111111111;
assign micromatrizz[65][7] = 9'b111111111;
assign micromatrizz[65][8] = 9'b111111111;
assign micromatrizz[65][9] = 9'b111111111;
assign micromatrizz[65][10] = 9'b111111111;
assign micromatrizz[65][11] = 9'b111111111;
assign micromatrizz[65][12] = 9'b111111111;
assign micromatrizz[65][13] = 9'b111110010;
assign micromatrizz[65][14] = 9'b111110010;
assign micromatrizz[65][15] = 9'b111110011;
assign micromatrizz[65][16] = 9'b111110011;
assign micromatrizz[65][17] = 9'b111110011;
assign micromatrizz[65][18] = 9'b111110011;
assign micromatrizz[65][19] = 9'b111110011;
assign micromatrizz[65][20] = 9'b111110011;
assign micromatrizz[65][21] = 9'b111111111;
assign micromatrizz[65][22] = 9'b111111111;
assign micromatrizz[65][23] = 9'b111111111;
assign micromatrizz[65][24] = 9'b111110010;
assign micromatrizz[65][25] = 9'b111110010;
assign micromatrizz[65][26] = 9'b111110010;
assign micromatrizz[65][27] = 9'b111110011;
assign micromatrizz[65][28] = 9'b111110011;
assign micromatrizz[65][29] = 9'b111110011;
assign micromatrizz[65][30] = 9'b111110011;
assign micromatrizz[65][31] = 9'b111111111;
assign micromatrizz[65][32] = 9'b111111111;
assign micromatrizz[65][33] = 9'b111111111;
assign micromatrizz[65][34] = 9'b111111111;
assign micromatrizz[65][35] = 9'b111110111;
assign micromatrizz[65][36] = 9'b111110010;
assign micromatrizz[65][37] = 9'b111110011;
assign micromatrizz[65][38] = 9'b111110011;
assign micromatrizz[65][39] = 9'b111110011;
assign micromatrizz[65][40] = 9'b111110011;
assign micromatrizz[65][41] = 9'b111110011;
assign micromatrizz[65][42] = 9'b111110011;
assign micromatrizz[65][43] = 9'b111111111;
assign micromatrizz[65][44] = 9'b111111111;
assign micromatrizz[65][45] = 9'b111111111;
assign micromatrizz[65][46] = 9'b111111111;
assign micromatrizz[65][47] = 9'b111110010;
assign micromatrizz[65][48] = 9'b111110010;
assign micromatrizz[65][49] = 9'b111110010;
assign micromatrizz[65][50] = 9'b111110011;
assign micromatrizz[65][51] = 9'b111110011;
assign micromatrizz[65][52] = 9'b111110011;
assign micromatrizz[65][53] = 9'b111110011;
assign micromatrizz[65][54] = 9'b111110010;
assign micromatrizz[65][55] = 9'b111110111;
assign micromatrizz[65][56] = 9'b111111111;
assign micromatrizz[65][57] = 9'b111111111;
assign micromatrizz[65][58] = 9'b111111111;
assign micromatrizz[65][59] = 9'b111110010;
assign micromatrizz[65][60] = 9'b111110010;
assign micromatrizz[65][61] = 9'b111110010;
assign micromatrizz[65][62] = 9'b111110011;
assign micromatrizz[65][63] = 9'b111110011;
assign micromatrizz[65][64] = 9'b111110010;
assign micromatrizz[65][65] = 9'b111111111;
assign micromatrizz[65][66] = 9'b111111111;
assign micromatrizz[65][67] = 9'b111111111;
assign micromatrizz[65][68] = 9'b111111111;
assign micromatrizz[65][69] = 9'b111110111;
assign micromatrizz[65][70] = 9'b111110010;
assign micromatrizz[65][71] = 9'b111110010;
assign micromatrizz[65][72] = 9'b111110011;
assign micromatrizz[65][73] = 9'b111110011;
assign micromatrizz[65][74] = 9'b111110011;
assign micromatrizz[65][75] = 9'b111111111;
assign micromatrizz[65][76] = 9'b111111111;
assign micromatrizz[65][77] = 9'b111111111;
assign micromatrizz[65][78] = 9'b111111111;
assign micromatrizz[65][79] = 9'b111111111;
assign micromatrizz[65][80] = 9'b111111111;
assign micromatrizz[65][81] = 9'b111111111;
assign micromatrizz[65][82] = 9'b111111111;
assign micromatrizz[65][83] = 9'b111110111;
assign micromatrizz[65][84] = 9'b111110111;
assign micromatrizz[65][85] = 9'b111111111;
assign micromatrizz[65][86] = 9'b111111111;
assign micromatrizz[65][87] = 9'b111111111;
assign micromatrizz[65][88] = 9'b111110110;
assign micromatrizz[65][89] = 9'b111110010;
assign micromatrizz[65][90] = 9'b111110010;
assign micromatrizz[65][91] = 9'b111110011;
assign micromatrizz[65][92] = 9'b111110011;
assign micromatrizz[65][93] = 9'b111110011;
assign micromatrizz[65][94] = 9'b111110011;
assign micromatrizz[65][95] = 9'b111110111;
assign micromatrizz[65][96] = 9'b111111111;
assign micromatrizz[65][97] = 9'b111111111;
assign micromatrizz[65][98] = 9'b111111111;
assign micromatrizz[65][99] = 9'b111111111;
assign micromatrizz[65][100] = 9'b111111111;
assign micromatrizz[65][101] = 9'b111111111;
assign micromatrizz[65][102] = 9'b111111111;
assign micromatrizz[65][103] = 9'b111111111;
assign micromatrizz[65][104] = 9'b111111111;
assign micromatrizz[65][105] = 9'b111111111;
assign micromatrizz[65][106] = 9'b111111111;
assign micromatrizz[65][107] = 9'b111111111;
assign micromatrizz[65][108] = 9'b111111111;
assign micromatrizz[65][109] = 9'b111110010;
assign micromatrizz[65][110] = 9'b111110010;
assign micromatrizz[65][111] = 9'b111110011;
assign micromatrizz[65][112] = 9'b111110010;
assign micromatrizz[65][113] = 9'b111110010;
assign micromatrizz[65][114] = 9'b111110011;
assign micromatrizz[65][115] = 9'b111110011;
assign micromatrizz[65][116] = 9'b111110011;
assign micromatrizz[65][117] = 9'b111111111;
assign micromatrizz[65][118] = 9'b111111111;
assign micromatrizz[65][119] = 9'b111111111;
assign micromatrizz[65][120] = 9'b111110010;
assign micromatrizz[65][121] = 9'b111110010;
assign micromatrizz[65][122] = 9'b111110010;
assign micromatrizz[65][123] = 9'b111110010;
assign micromatrizz[65][124] = 9'b111110011;
assign micromatrizz[65][125] = 9'b111110011;
assign micromatrizz[65][126] = 9'b111110011;
assign micromatrizz[65][127] = 9'b111111111;
assign micromatrizz[65][128] = 9'b111111111;
assign micromatrizz[65][129] = 9'b111111111;
assign micromatrizz[65][130] = 9'b111111111;
assign micromatrizz[65][131] = 9'b111111111;
assign micromatrizz[65][132] = 9'b111111111;
assign micromatrizz[65][133] = 9'b111111111;
assign micromatrizz[65][134] = 9'b111110111;
assign micromatrizz[65][135] = 9'b111111111;
assign micromatrizz[65][136] = 9'b111111111;
assign micromatrizz[65][137] = 9'b111111111;
assign micromatrizz[65][138] = 9'b111110111;
assign micromatrizz[65][139] = 9'b111110010;
assign micromatrizz[65][140] = 9'b111110010;
assign micromatrizz[65][141] = 9'b111110010;
assign micromatrizz[65][142] = 9'b111110010;
assign micromatrizz[65][143] = 9'b111110011;
assign micromatrizz[65][144] = 9'b111110011;
assign micromatrizz[65][145] = 9'b111110011;
assign micromatrizz[65][146] = 9'b111111111;
assign micromatrizz[65][147] = 9'b111111111;
assign micromatrizz[65][148] = 9'b111111111;
assign micromatrizz[65][149] = 9'b111111111;
assign micromatrizz[65][150] = 9'b111110111;
assign micromatrizz[65][151] = 9'b111110010;
assign micromatrizz[65][152] = 9'b111110010;
assign micromatrizz[65][153] = 9'b111110011;
assign micromatrizz[65][154] = 9'b111110011;
assign micromatrizz[65][155] = 9'b111110011;
assign micromatrizz[65][156] = 9'b111110011;
assign micromatrizz[65][157] = 9'b111110111;
assign micromatrizz[65][158] = 9'b111111111;
assign micromatrizz[65][159] = 9'b111111111;
assign micromatrizz[65][160] = 9'b111111111;
assign micromatrizz[65][161] = 9'b111110010;
assign micromatrizz[65][162] = 9'b111110010;
assign micromatrizz[65][163] = 9'b111110010;
assign micromatrizz[65][164] = 9'b111110011;
assign micromatrizz[65][165] = 9'b111110011;
assign micromatrizz[65][166] = 9'b111110011;
assign micromatrizz[65][167] = 9'b111110011;
assign micromatrizz[65][168] = 9'b111111111;
assign micromatrizz[65][169] = 9'b111111111;
assign micromatrizz[65][170] = 9'b111111111;
assign micromatrizz[65][171] = 9'b111111111;
assign micromatrizz[65][172] = 9'b111110010;
assign micromatrizz[65][173] = 9'b111110010;
assign micromatrizz[65][174] = 9'b111110011;
assign micromatrizz[65][175] = 9'b111110011;
assign micromatrizz[65][176] = 9'b111110011;
assign micromatrizz[65][177] = 9'b111110011;
assign micromatrizz[65][178] = 9'b111110010;
assign micromatrizz[65][179] = 9'b111110111;
assign micromatrizz[65][180] = 9'b111111111;
assign micromatrizz[65][181] = 9'b111111111;
assign micromatrizz[65][182] = 9'b111111111;
assign micromatrizz[65][183] = 9'b111110111;
assign micromatrizz[65][184] = 9'b111110010;
assign micromatrizz[65][185] = 9'b111110011;
assign micromatrizz[65][186] = 9'b111110010;
assign micromatrizz[65][187] = 9'b111110010;
assign micromatrizz[65][188] = 9'b111110011;
assign micromatrizz[65][189] = 9'b111110011;
assign micromatrizz[65][190] = 9'b111111111;
assign micromatrizz[65][191] = 9'b111111111;
assign micromatrizz[65][192] = 9'b111111111;
assign micromatrizz[65][193] = 9'b111111111;
assign micromatrizz[65][194] = 9'b111111111;
assign micromatrizz[65][195] = 9'b111110110;
assign micromatrizz[65][196] = 9'b111110010;
assign micromatrizz[65][197] = 9'b111110011;
assign micromatrizz[65][198] = 9'b111110011;
assign micromatrizz[65][199] = 9'b111110010;
assign micromatrizz[65][200] = 9'b111110010;
assign micromatrizz[65][201] = 9'b111110011;
assign micromatrizz[65][202] = 9'b111110111;
assign micromatrizz[65][203] = 9'b111111111;
assign micromatrizz[65][204] = 9'b111111111;
assign micromatrizz[65][205] = 9'b111111111;
assign micromatrizz[65][206] = 9'b111111111;
assign micromatrizz[65][207] = 9'b111110010;
assign micromatrizz[65][208] = 9'b111110010;
assign micromatrizz[65][209] = 9'b111110010;
assign micromatrizz[65][210] = 9'b111110010;
assign micromatrizz[65][211] = 9'b111110011;
assign micromatrizz[65][212] = 9'b111110011;
assign micromatrizz[65][213] = 9'b111110111;
assign micromatrizz[65][214] = 9'b111111111;
assign micromatrizz[65][215] = 9'b111111111;
assign micromatrizz[65][216] = 9'b111111111;
assign micromatrizz[65][217] = 9'b111111111;
assign micromatrizz[65][218] = 9'b111111111;
assign micromatrizz[65][219] = 9'b111111111;
assign micromatrizz[65][220] = 9'b111110111;
assign micromatrizz[65][221] = 9'b111111111;
assign micromatrizz[65][222] = 9'b111111111;
assign micromatrizz[65][223] = 9'b111111111;
assign micromatrizz[65][224] = 9'b111111111;
assign micromatrizz[65][225] = 9'b111110110;
assign micromatrizz[65][226] = 9'b111110010;
assign micromatrizz[65][227] = 9'b111110010;
assign micromatrizz[65][228] = 9'b111110010;
assign micromatrizz[65][229] = 9'b111110011;
assign micromatrizz[65][230] = 9'b111110011;
assign micromatrizz[65][231] = 9'b111110011;
assign micromatrizz[65][232] = 9'b111110111;
assign micromatrizz[65][233] = 9'b111111111;
assign micromatrizz[65][234] = 9'b111111111;
assign micromatrizz[65][235] = 9'b111111111;
assign micromatrizz[65][236] = 9'b111111111;
assign micromatrizz[65][237] = 9'b111111111;
assign micromatrizz[65][238] = 9'b111111111;
assign micromatrizz[65][239] = 9'b111111111;
assign micromatrizz[65][240] = 9'b111111111;
assign micromatrizz[65][241] = 9'b111111111;
assign micromatrizz[65][242] = 9'b111110010;
assign micromatrizz[65][243] = 9'b111110010;
assign micromatrizz[65][244] = 9'b111110010;
assign micromatrizz[65][245] = 9'b111110010;
assign micromatrizz[65][246] = 9'b111110010;
assign micromatrizz[65][247] = 9'b111110111;
assign micromatrizz[65][248] = 9'b111111111;
assign micromatrizz[65][249] = 9'b111111111;
assign micromatrizz[65][250] = 9'b111111111;
assign micromatrizz[65][251] = 9'b111111111;
assign micromatrizz[65][252] = 9'b111111111;
assign micromatrizz[65][253] = 9'b111111111;
assign micromatrizz[65][254] = 9'b111111111;
assign micromatrizz[65][255] = 9'b111111111;
assign micromatrizz[65][256] = 9'b111110110;
assign micromatrizz[65][257] = 9'b111111111;
assign micromatrizz[65][258] = 9'b111111111;
assign micromatrizz[65][259] = 9'b111111111;
assign micromatrizz[65][260] = 9'b111111111;
assign micromatrizz[65][261] = 9'b111111111;
assign micromatrizz[65][262] = 9'b111111111;
assign micromatrizz[65][263] = 9'b111111111;
assign micromatrizz[65][264] = 9'b111111111;
assign micromatrizz[65][265] = 9'b111110010;
assign micromatrizz[65][266] = 9'b111110011;
assign micromatrizz[65][267] = 9'b111110011;
assign micromatrizz[65][268] = 9'b111110010;
assign micromatrizz[65][269] = 9'b111110011;
assign micromatrizz[65][270] = 9'b111110011;
assign micromatrizz[65][271] = 9'b111110010;
assign micromatrizz[65][272] = 9'b111110111;
assign micromatrizz[65][273] = 9'b111111111;
assign micromatrizz[65][274] = 9'b111111111;
assign micromatrizz[65][275] = 9'b111110010;
assign micromatrizz[65][276] = 9'b111110010;
assign micromatrizz[65][277] = 9'b111110010;
assign micromatrizz[65][278] = 9'b111110011;
assign micromatrizz[65][279] = 9'b111110011;
assign micromatrizz[65][280] = 9'b111110011;
assign micromatrizz[65][281] = 9'b111110011;
assign micromatrizz[65][282] = 9'b111111111;
assign micromatrizz[65][283] = 9'b111111111;
assign micromatrizz[65][284] = 9'b111111111;
assign micromatrizz[65][285] = 9'b111111111;
assign micromatrizz[65][286] = 9'b111110010;
assign micromatrizz[65][287] = 9'b111110010;
assign micromatrizz[65][288] = 9'b111110010;
assign micromatrizz[65][289] = 9'b111110011;
assign micromatrizz[65][290] = 9'b111110011;
assign micromatrizz[65][291] = 9'b111110011;
assign micromatrizz[65][292] = 9'b111110011;
assign micromatrizz[65][293] = 9'b111110111;
assign micromatrizz[65][294] = 9'b111111111;
assign micromatrizz[65][295] = 9'b111111111;
assign micromatrizz[65][296] = 9'b111111111;
assign micromatrizz[65][297] = 9'b111111111;
assign micromatrizz[65][298] = 9'b111111111;
assign micromatrizz[65][299] = 9'b111111111;
assign micromatrizz[65][300] = 9'b111111111;
assign micromatrizz[65][301] = 9'b111111111;
assign micromatrizz[65][302] = 9'b111111111;
assign micromatrizz[65][303] = 9'b111110010;
assign micromatrizz[65][304] = 9'b111110011;
assign micromatrizz[65][305] = 9'b111110011;
assign micromatrizz[65][306] = 9'b111110010;
assign micromatrizz[65][307] = 9'b111110011;
assign micromatrizz[65][308] = 9'b111111111;
assign micromatrizz[65][309] = 9'b111111111;
assign micromatrizz[65][310] = 9'b111111111;
assign micromatrizz[65][311] = 9'b111111111;
assign micromatrizz[65][312] = 9'b111111111;
assign micromatrizz[65][313] = 9'b111111111;
assign micromatrizz[65][314] = 9'b111111111;
assign micromatrizz[65][315] = 9'b111111111;
assign micromatrizz[65][316] = 9'b111110111;
assign micromatrizz[65][317] = 9'b111110010;
assign micromatrizz[65][318] = 9'b111110010;
assign micromatrizz[65][319] = 9'b111110011;
assign micromatrizz[65][320] = 9'b111110011;
assign micromatrizz[65][321] = 9'b111110011;
assign micromatrizz[65][322] = 9'b111111111;
assign micromatrizz[65][323] = 9'b111111111;
assign micromatrizz[65][324] = 9'b111111111;
assign micromatrizz[65][325] = 9'b111111111;
assign micromatrizz[65][326] = 9'b111111111;
assign micromatrizz[65][327] = 9'b111111111;
assign micromatrizz[65][328] = 9'b111111111;
assign micromatrizz[65][329] = 9'b111111111;
assign micromatrizz[65][330] = 9'b111110111;
assign micromatrizz[65][331] = 9'b111110111;
assign micromatrizz[65][332] = 9'b111111111;
assign micromatrizz[65][333] = 9'b111111111;
assign micromatrizz[65][334] = 9'b111111111;
assign micromatrizz[65][335] = 9'b111110010;
assign micromatrizz[65][336] = 9'b111110011;
assign micromatrizz[65][337] = 9'b111110011;
assign micromatrizz[65][338] = 9'b111110011;
assign micromatrizz[65][339] = 9'b111110010;
assign micromatrizz[65][340] = 9'b111110010;
assign micromatrizz[65][341] = 9'b111110010;
assign micromatrizz[65][342] = 9'b111111111;
assign micromatrizz[65][343] = 9'b111111111;
assign micromatrizz[65][344] = 9'b111111111;
assign micromatrizz[65][345] = 9'b111111111;
assign micromatrizz[65][346] = 9'b111111111;
assign micromatrizz[65][347] = 9'b111110010;
assign micromatrizz[65][348] = 9'b111110010;
assign micromatrizz[65][349] = 9'b111110010;
assign micromatrizz[65][350] = 9'b111110010;
assign micromatrizz[65][351] = 9'b111110011;
assign micromatrizz[65][352] = 9'b111110011;
assign micromatrizz[65][353] = 9'b111110011;
assign micromatrizz[65][354] = 9'b111111111;
assign micromatrizz[65][355] = 9'b111111111;
assign micromatrizz[65][356] = 9'b111111111;
assign micromatrizz[65][357] = 9'b111111111;
assign micromatrizz[65][358] = 9'b111111111;
assign micromatrizz[65][359] = 9'b111110010;
assign micromatrizz[65][360] = 9'b111110011;
assign micromatrizz[65][361] = 9'b111110010;
assign micromatrizz[65][362] = 9'b111110010;
assign micromatrizz[65][363] = 9'b111110010;
assign micromatrizz[65][364] = 9'b111110011;
assign micromatrizz[65][365] = 9'b111110010;
assign micromatrizz[65][366] = 9'b111111111;
assign micromatrizz[65][367] = 9'b111111111;
assign micromatrizz[65][368] = 9'b111111111;
assign micromatrizz[65][369] = 9'b111110010;
assign micromatrizz[65][370] = 9'b111111111;
assign micromatrizz[65][371] = 9'b111110111;
assign micromatrizz[65][372] = 9'b111110010;
assign micromatrizz[65][373] = 9'b111110011;
assign micromatrizz[65][374] = 9'b111110011;
assign micromatrizz[65][375] = 9'b111110011;
assign micromatrizz[65][376] = 9'b111110011;
assign micromatrizz[65][377] = 9'b111110010;
assign micromatrizz[65][378] = 9'b111110010;
assign micromatrizz[65][379] = 9'b111111111;
assign micromatrizz[65][380] = 9'b111111111;
assign micromatrizz[65][381] = 9'b111111111;
assign micromatrizz[65][382] = 9'b111111111;
assign micromatrizz[65][383] = 9'b111111111;
assign micromatrizz[65][384] = 9'b111110010;
assign micromatrizz[65][385] = 9'b111110010;
assign micromatrizz[65][386] = 9'b111110011;
assign micromatrizz[65][387] = 9'b111110011;
assign micromatrizz[65][388] = 9'b111110011;
assign micromatrizz[65][389] = 9'b111110011;
assign micromatrizz[65][390] = 9'b111110011;
assign micromatrizz[65][391] = 9'b111111111;
assign micromatrizz[65][392] = 9'b111111111;
assign micromatrizz[65][393] = 9'b111111111;
assign micromatrizz[65][394] = 9'b111111111;
assign micromatrizz[65][395] = 9'b111110010;
assign micromatrizz[65][396] = 9'b111110010;
assign micromatrizz[65][397] = 9'b111110010;
assign micromatrizz[65][398] = 9'b111110010;
assign micromatrizz[65][399] = 9'b111110011;
assign micromatrizz[65][400] = 9'b111110011;
assign micromatrizz[65][401] = 9'b111110011;
assign micromatrizz[65][402] = 9'b111110111;
assign micromatrizz[65][403] = 9'b111111111;
assign micromatrizz[65][404] = 9'b111111111;
assign micromatrizz[65][405] = 9'b111111111;
assign micromatrizz[65][406] = 9'b111111111;
assign micromatrizz[65][407] = 9'b111111111;
assign micromatrizz[65][408] = 9'b111111111;
assign micromatrizz[65][409] = 9'b111111111;
assign micromatrizz[65][410] = 9'b111111111;
assign micromatrizz[65][411] = 9'b111111111;
assign micromatrizz[65][412] = 9'b111110010;
assign micromatrizz[65][413] = 9'b111110010;
assign micromatrizz[65][414] = 9'b111110010;
assign micromatrizz[65][415] = 9'b111110011;
assign micromatrizz[65][416] = 9'b111110011;
assign micromatrizz[65][417] = 9'b111110111;
assign micromatrizz[65][418] = 9'b111111111;
assign micromatrizz[65][419] = 9'b111111111;
assign micromatrizz[65][420] = 9'b111111111;
assign micromatrizz[65][421] = 9'b111111111;
assign micromatrizz[65][422] = 9'b111111111;
assign micromatrizz[65][423] = 9'b111111111;
assign micromatrizz[65][424] = 9'b111111111;
assign micromatrizz[65][425] = 9'b111111111;
assign micromatrizz[65][426] = 9'b111110010;
assign micromatrizz[65][427] = 9'b111111111;
assign micromatrizz[65][428] = 9'b111111111;
assign micromatrizz[65][429] = 9'b111111111;
assign micromatrizz[65][430] = 9'b111110111;
assign micromatrizz[65][431] = 9'b111110010;
assign micromatrizz[65][432] = 9'b111110010;
assign micromatrizz[65][433] = 9'b111110010;
assign micromatrizz[65][434] = 9'b111110010;
assign micromatrizz[65][435] = 9'b111110011;
assign micromatrizz[65][436] = 9'b111110011;
assign micromatrizz[65][437] = 9'b111110011;
assign micromatrizz[65][438] = 9'b111111111;
assign micromatrizz[65][439] = 9'b111111111;
assign micromatrizz[65][440] = 9'b111111111;
assign micromatrizz[65][441] = 9'b111111111;
assign micromatrizz[65][442] = 9'b111111111;
assign micromatrizz[65][443] = 9'b111111111;
assign micromatrizz[65][444] = 9'b111111111;
assign micromatrizz[65][445] = 9'b111111111;
assign micromatrizz[65][446] = 9'b111111111;
assign micromatrizz[65][447] = 9'b111110111;
assign micromatrizz[65][448] = 9'b111110010;
assign micromatrizz[65][449] = 9'b111110010;
assign micromatrizz[65][450] = 9'b111110010;
assign micromatrizz[65][451] = 9'b111110011;
assign micromatrizz[65][452] = 9'b111110011;
assign micromatrizz[65][453] = 9'b111110011;
assign micromatrizz[65][454] = 9'b111111111;
assign micromatrizz[65][455] = 9'b111111111;
assign micromatrizz[65][456] = 9'b111111111;
assign micromatrizz[65][457] = 9'b111111111;
assign micromatrizz[65][458] = 9'b111111111;
assign micromatrizz[65][459] = 9'b111111111;
assign micromatrizz[65][460] = 9'b111111111;
assign micromatrizz[65][461] = 9'b111110111;
assign micromatrizz[65][462] = 9'b111111111;
assign micromatrizz[65][463] = 9'b111111111;
assign micromatrizz[65][464] = 9'b111111111;
assign micromatrizz[65][465] = 9'b111111111;
assign micromatrizz[65][466] = 9'b111111111;
assign micromatrizz[65][467] = 9'b111111111;
assign micromatrizz[65][468] = 9'b111111111;
assign micromatrizz[65][469] = 9'b111111111;
assign micromatrizz[65][470] = 9'b111110010;
assign micromatrizz[65][471] = 9'b111110010;
assign micromatrizz[65][472] = 9'b111110011;
assign micromatrizz[65][473] = 9'b111110010;
assign micromatrizz[65][474] = 9'b111110011;
assign micromatrizz[65][475] = 9'b111110011;
assign micromatrizz[65][476] = 9'b111110011;
assign micromatrizz[65][477] = 9'b111110011;
assign micromatrizz[65][478] = 9'b111111111;
assign micromatrizz[65][479] = 9'b111111111;
assign micromatrizz[65][480] = 9'b111111111;
assign micromatrizz[65][481] = 9'b111110010;
assign micromatrizz[65][482] = 9'b111110010;
assign micromatrizz[65][483] = 9'b111110010;
assign micromatrizz[65][484] = 9'b111110010;
assign micromatrizz[65][485] = 9'b111110011;
assign micromatrizz[65][486] = 9'b111110011;
assign micromatrizz[65][487] = 9'b111110011;
assign micromatrizz[65][488] = 9'b111110111;
assign micromatrizz[65][489] = 9'b111111111;
assign micromatrizz[65][490] = 9'b111111111;
assign micromatrizz[65][491] = 9'b111111111;
assign micromatrizz[65][492] = 9'b111111111;
assign micromatrizz[65][493] = 9'b111111111;
assign micromatrizz[65][494] = 9'b111111111;
assign micromatrizz[65][495] = 9'b111111111;
assign micromatrizz[65][496] = 9'b111111111;
assign micromatrizz[65][497] = 9'b111111111;
assign micromatrizz[65][498] = 9'b111110010;
assign micromatrizz[65][499] = 9'b111110010;
assign micromatrizz[65][500] = 9'b111110010;
assign micromatrizz[65][501] = 9'b111110010;
assign micromatrizz[65][502] = 9'b111110010;
assign micromatrizz[65][503] = 9'b111110111;
assign micromatrizz[65][504] = 9'b111111111;
assign micromatrizz[65][505] = 9'b111111111;
assign micromatrizz[65][506] = 9'b111111111;
assign micromatrizz[65][507] = 9'b111111111;
assign micromatrizz[65][508] = 9'b111111111;
assign micromatrizz[65][509] = 9'b111111111;
assign micromatrizz[65][510] = 9'b111111111;
assign micromatrizz[65][511] = 9'b111110111;
assign micromatrizz[65][512] = 9'b111110010;
assign micromatrizz[65][513] = 9'b111111111;
assign micromatrizz[65][514] = 9'b111111111;
assign micromatrizz[65][515] = 9'b111111111;
assign micromatrizz[65][516] = 9'b111110111;
assign micromatrizz[65][517] = 9'b111110010;
assign micromatrizz[65][518] = 9'b111110011;
assign micromatrizz[65][519] = 9'b111110011;
assign micromatrizz[65][520] = 9'b111110010;
assign micromatrizz[65][521] = 9'b111110010;
assign micromatrizz[65][522] = 9'b111110011;
assign micromatrizz[65][523] = 9'b111110111;
assign micromatrizz[65][524] = 9'b111111111;
assign micromatrizz[65][525] = 9'b111111111;
assign micromatrizz[65][526] = 9'b111111111;
assign micromatrizz[65][527] = 9'b111111111;
assign micromatrizz[65][528] = 9'b111110111;
assign micromatrizz[65][529] = 9'b111110010;
assign micromatrizz[65][530] = 9'b111110010;
assign micromatrizz[65][531] = 9'b111110010;
assign micromatrizz[65][532] = 9'b111110011;
assign micromatrizz[65][533] = 9'b111110011;
assign micromatrizz[65][534] = 9'b111110011;
assign micromatrizz[65][535] = 9'b111110111;
assign micromatrizz[65][536] = 9'b111111111;
assign micromatrizz[65][537] = 9'b111111111;
assign micromatrizz[65][538] = 9'b111111111;
assign micromatrizz[65][539] = 9'b111110111;
assign micromatrizz[65][540] = 9'b111110010;
assign micromatrizz[65][541] = 9'b111110011;
assign micromatrizz[65][542] = 9'b111110011;
assign micromatrizz[65][543] = 9'b111110011;
assign micromatrizz[65][544] = 9'b111110011;
assign micromatrizz[65][545] = 9'b111111111;
assign micromatrizz[65][546] = 9'b111111111;
assign micromatrizz[65][547] = 9'b111111111;
assign micromatrizz[65][548] = 9'b111111111;
assign micromatrizz[65][549] = 9'b111111111;
assign micromatrizz[65][550] = 9'b111111111;
assign micromatrizz[65][551] = 9'b111111111;
assign micromatrizz[65][552] = 9'b111111111;
assign micromatrizz[65][553] = 9'b111110111;
assign micromatrizz[65][554] = 9'b111110111;
assign micromatrizz[65][555] = 9'b111111111;
assign micromatrizz[65][556] = 9'b111111111;
assign micromatrizz[65][557] = 9'b111111111;
assign micromatrizz[65][558] = 9'b111110010;
assign micromatrizz[65][559] = 9'b111110010;
assign micromatrizz[65][560] = 9'b111110010;
assign micromatrizz[65][561] = 9'b111110010;
assign micromatrizz[65][562] = 9'b111110011;
assign micromatrizz[65][563] = 9'b111110011;
assign micromatrizz[65][564] = 9'b111110010;
assign micromatrizz[65][565] = 9'b111111111;
assign micromatrizz[65][566] = 9'b111111111;
assign micromatrizz[65][567] = 9'b111111111;
assign micromatrizz[65][568] = 9'b111111111;
assign micromatrizz[65][569] = 9'b111110111;
assign micromatrizz[65][570] = 9'b111110010;
assign micromatrizz[65][571] = 9'b111110010;
assign micromatrizz[65][572] = 9'b111110010;
assign micromatrizz[65][573] = 9'b111110011;
assign micromatrizz[65][574] = 9'b111110011;
assign micromatrizz[65][575] = 9'b111110011;
assign micromatrizz[65][576] = 9'b111111111;
assign micromatrizz[65][577] = 9'b111111111;
assign micromatrizz[65][578] = 9'b111111111;
assign micromatrizz[65][579] = 9'b111111111;
assign micromatrizz[65][580] = 9'b111111111;
assign micromatrizz[65][581] = 9'b111110010;
assign micromatrizz[65][582] = 9'b111110011;
assign micromatrizz[65][583] = 9'b111110011;
assign micromatrizz[65][584] = 9'b111110011;
assign micromatrizz[65][585] = 9'b111110011;
assign micromatrizz[65][586] = 9'b111110011;
assign micromatrizz[65][587] = 9'b111110011;
assign micromatrizz[65][588] = 9'b111111111;
assign micromatrizz[65][589] = 9'b111111111;
assign micromatrizz[65][590] = 9'b111111111;
assign micromatrizz[65][591] = 9'b111111111;
assign micromatrizz[65][592] = 9'b111110111;
assign micromatrizz[65][593] = 9'b111110010;
assign micromatrizz[65][594] = 9'b111110010;
assign micromatrizz[65][595] = 9'b111110011;
assign micromatrizz[65][596] = 9'b111110011;
assign micromatrizz[65][597] = 9'b111110010;
assign micromatrizz[65][598] = 9'b111111111;
assign micromatrizz[65][599] = 9'b111111111;
assign micromatrizz[65][600] = 9'b111111111;
assign micromatrizz[65][601] = 9'b111111111;
assign micromatrizz[65][602] = 9'b111111111;
assign micromatrizz[65][603] = 9'b111111111;
assign micromatrizz[65][604] = 9'b111111111;
assign micromatrizz[65][605] = 9'b111111111;
assign micromatrizz[65][606] = 9'b111110111;
assign micromatrizz[65][607] = 9'b111110111;
assign micromatrizz[65][608] = 9'b111111111;
assign micromatrizz[65][609] = 9'b111111111;
assign micromatrizz[65][610] = 9'b111111111;
assign micromatrizz[65][611] = 9'b111111111;
assign micromatrizz[65][612] = 9'b111111111;
assign micromatrizz[65][613] = 9'b111111111;
assign micromatrizz[65][614] = 9'b111111111;
assign micromatrizz[65][615] = 9'b111110111;
assign micromatrizz[65][616] = 9'b111110010;
assign micromatrizz[65][617] = 9'b111110010;
assign micromatrizz[65][618] = 9'b111110010;
assign micromatrizz[65][619] = 9'b111110011;
assign micromatrizz[65][620] = 9'b111110011;
assign micromatrizz[65][621] = 9'b111110011;
assign micromatrizz[65][622] = 9'b111110011;
assign micromatrizz[65][623] = 9'b111111111;
assign micromatrizz[65][624] = 9'b111111111;
assign micromatrizz[65][625] = 9'b111111111;
assign micromatrizz[65][626] = 9'b111111111;
assign micromatrizz[65][627] = 9'b111111111;
assign micromatrizz[65][628] = 9'b111111111;
assign micromatrizz[65][629] = 9'b111111111;
assign micromatrizz[65][630] = 9'b111111111;
assign micromatrizz[65][631] = 9'b111111111;
assign micromatrizz[65][632] = 9'b111111111;
assign micromatrizz[65][633] = 9'b111111111;
assign micromatrizz[65][634] = 9'b111111111;
assign micromatrizz[65][635] = 9'b111111111;
assign micromatrizz[65][636] = 9'b111111111;
assign micromatrizz[65][637] = 9'b111111111;
assign micromatrizz[65][638] = 9'b111111111;
assign micromatrizz[65][639] = 9'b111111111;
assign micromatrizz[66][0] = 9'b111111111;
assign micromatrizz[66][1] = 9'b111111111;
assign micromatrizz[66][2] = 9'b111111111;
assign micromatrizz[66][3] = 9'b111111111;
assign micromatrizz[66][4] = 9'b111111111;
assign micromatrizz[66][5] = 9'b111111111;
assign micromatrizz[66][6] = 9'b111111111;
assign micromatrizz[66][7] = 9'b111111111;
assign micromatrizz[66][8] = 9'b111111111;
assign micromatrizz[66][9] = 9'b111111111;
assign micromatrizz[66][10] = 9'b111111111;
assign micromatrizz[66][11] = 9'b111111111;
assign micromatrizz[66][12] = 9'b111111111;
assign micromatrizz[66][13] = 9'b111111111;
assign micromatrizz[66][14] = 9'b111110010;
assign micromatrizz[66][15] = 9'b111110010;
assign micromatrizz[66][16] = 9'b111110011;
assign micromatrizz[66][17] = 9'b111110011;
assign micromatrizz[66][18] = 9'b111110011;
assign micromatrizz[66][19] = 9'b111110010;
assign micromatrizz[66][20] = 9'b111110111;
assign micromatrizz[66][21] = 9'b111111111;
assign micromatrizz[66][22] = 9'b111111111;
assign micromatrizz[66][23] = 9'b111111111;
assign micromatrizz[66][24] = 9'b111110010;
assign micromatrizz[66][25] = 9'b111110010;
assign micromatrizz[66][26] = 9'b111110010;
assign micromatrizz[66][27] = 9'b111110011;
assign micromatrizz[66][28] = 9'b111110011;
assign micromatrizz[66][29] = 9'b111110011;
assign micromatrizz[66][30] = 9'b111110011;
assign micromatrizz[66][31] = 9'b111111111;
assign micromatrizz[66][32] = 9'b111111111;
assign micromatrizz[66][33] = 9'b111111111;
assign micromatrizz[66][34] = 9'b111111111;
assign micromatrizz[66][35] = 9'b111110111;
assign micromatrizz[66][36] = 9'b111110010;
assign micromatrizz[66][37] = 9'b111110011;
assign micromatrizz[66][38] = 9'b111110011;
assign micromatrizz[66][39] = 9'b111110011;
assign micromatrizz[66][40] = 9'b111110011;
assign micromatrizz[66][41] = 9'b111110011;
assign micromatrizz[66][42] = 9'b111110011;
assign micromatrizz[66][43] = 9'b111111111;
assign micromatrizz[66][44] = 9'b111111111;
assign micromatrizz[66][45] = 9'b111111111;
assign micromatrizz[66][46] = 9'b111111111;
assign micromatrizz[66][47] = 9'b111110010;
assign micromatrizz[66][48] = 9'b111110010;
assign micromatrizz[66][49] = 9'b111110011;
assign micromatrizz[66][50] = 9'b111110011;
assign micromatrizz[66][51] = 9'b111110011;
assign micromatrizz[66][52] = 9'b111110010;
assign micromatrizz[66][53] = 9'b111110011;
assign micromatrizz[66][54] = 9'b111110111;
assign micromatrizz[66][55] = 9'b111110111;
assign micromatrizz[66][56] = 9'b111110111;
assign micromatrizz[66][57] = 9'b111111111;
assign micromatrizz[66][58] = 9'b111110111;
assign micromatrizz[66][59] = 9'b111110010;
assign micromatrizz[66][60] = 9'b111110010;
assign micromatrizz[66][61] = 9'b111110010;
assign micromatrizz[66][62] = 9'b111110010;
assign micromatrizz[66][63] = 9'b111110011;
assign micromatrizz[66][64] = 9'b111111111;
assign micromatrizz[66][65] = 9'b111111111;
assign micromatrizz[66][66] = 9'b111111111;
assign micromatrizz[66][67] = 9'b111111111;
assign micromatrizz[66][68] = 9'b111111111;
assign micromatrizz[66][69] = 9'b111111111;
assign micromatrizz[66][70] = 9'b111110010;
assign micromatrizz[66][71] = 9'b111110010;
assign micromatrizz[66][72] = 9'b111110011;
assign micromatrizz[66][73] = 9'b111110011;
assign micromatrizz[66][74] = 9'b111110011;
assign micromatrizz[66][75] = 9'b111111111;
assign micromatrizz[66][76] = 9'b111111111;
assign micromatrizz[66][77] = 9'b111111111;
assign micromatrizz[66][78] = 9'b111111111;
assign micromatrizz[66][79] = 9'b111111111;
assign micromatrizz[66][80] = 9'b111111111;
assign micromatrizz[66][81] = 9'b111111111;
assign micromatrizz[66][82] = 9'b111110111;
assign micromatrizz[66][83] = 9'b111110010;
assign micromatrizz[66][84] = 9'b111111111;
assign micromatrizz[66][85] = 9'b111111111;
assign micromatrizz[66][86] = 9'b111111111;
assign micromatrizz[66][87] = 9'b111111111;
assign micromatrizz[66][88] = 9'b111110110;
assign micromatrizz[66][89] = 9'b111110010;
assign micromatrizz[66][90] = 9'b111110010;
assign micromatrizz[66][91] = 9'b111110011;
assign micromatrizz[66][92] = 9'b111110010;
assign micromatrizz[66][93] = 9'b111110011;
assign micromatrizz[66][94] = 9'b111110011;
assign micromatrizz[66][95] = 9'b111110111;
assign micromatrizz[66][96] = 9'b111111111;
assign micromatrizz[66][97] = 9'b111111111;
assign micromatrizz[66][98] = 9'b111111111;
assign micromatrizz[66][99] = 9'b111111111;
assign micromatrizz[66][100] = 9'b111111111;
assign micromatrizz[66][101] = 9'b111111111;
assign micromatrizz[66][102] = 9'b111111111;
assign micromatrizz[66][103] = 9'b111111111;
assign micromatrizz[66][104] = 9'b111111111;
assign micromatrizz[66][105] = 9'b111111111;
assign micromatrizz[66][106] = 9'b111111111;
assign micromatrizz[66][107] = 9'b111111111;
assign micromatrizz[66][108] = 9'b111111111;
assign micromatrizz[66][109] = 9'b111111111;
assign micromatrizz[66][110] = 9'b111110010;
assign micromatrizz[66][111] = 9'b111110010;
assign micromatrizz[66][112] = 9'b111110011;
assign micromatrizz[66][113] = 9'b111110011;
assign micromatrizz[66][114] = 9'b111110011;
assign micromatrizz[66][115] = 9'b111110011;
assign micromatrizz[66][116] = 9'b111110011;
assign micromatrizz[66][117] = 9'b111111111;
assign micromatrizz[66][118] = 9'b111111111;
assign micromatrizz[66][119] = 9'b111111111;
assign micromatrizz[66][120] = 9'b111110111;
assign micromatrizz[66][121] = 9'b111110010;
assign micromatrizz[66][122] = 9'b111110010;
assign micromatrizz[66][123] = 9'b111110010;
assign micromatrizz[66][124] = 9'b111110011;
assign micromatrizz[66][125] = 9'b111110011;
assign micromatrizz[66][126] = 9'b111110011;
assign micromatrizz[66][127] = 9'b111111111;
assign micromatrizz[66][128] = 9'b111111111;
assign micromatrizz[66][129] = 9'b111111111;
assign micromatrizz[66][130] = 9'b111111111;
assign micromatrizz[66][131] = 9'b111111111;
assign micromatrizz[66][132] = 9'b111111111;
assign micromatrizz[66][133] = 9'b111110110;
assign micromatrizz[66][134] = 9'b111111111;
assign micromatrizz[66][135] = 9'b111111111;
assign micromatrizz[66][136] = 9'b111111111;
assign micromatrizz[66][137] = 9'b111111111;
assign micromatrizz[66][138] = 9'b111110111;
assign micromatrizz[66][139] = 9'b111110010;
assign micromatrizz[66][140] = 9'b111110010;
assign micromatrizz[66][141] = 9'b111110010;
assign micromatrizz[66][142] = 9'b111110010;
assign micromatrizz[66][143] = 9'b111110011;
assign micromatrizz[66][144] = 9'b111110011;
assign micromatrizz[66][145] = 9'b111110011;
assign micromatrizz[66][146] = 9'b111111111;
assign micromatrizz[66][147] = 9'b111111111;
assign micromatrizz[66][148] = 9'b111111111;
assign micromatrizz[66][149] = 9'b111111111;
assign micromatrizz[66][150] = 9'b111110111;
assign micromatrizz[66][151] = 9'b111110010;
assign micromatrizz[66][152] = 9'b111110010;
assign micromatrizz[66][153] = 9'b111110011;
assign micromatrizz[66][154] = 9'b111110011;
assign micromatrizz[66][155] = 9'b111110011;
assign micromatrizz[66][156] = 9'b111110011;
assign micromatrizz[66][157] = 9'b111110111;
assign micromatrizz[66][158] = 9'b111111111;
assign micromatrizz[66][159] = 9'b111111111;
assign micromatrizz[66][160] = 9'b111111111;
assign micromatrizz[66][161] = 9'b111110010;
assign micromatrizz[66][162] = 9'b111110010;
assign micromatrizz[66][163] = 9'b111110010;
assign micromatrizz[66][164] = 9'b111110011;
assign micromatrizz[66][165] = 9'b111110011;
assign micromatrizz[66][166] = 9'b111110011;
assign micromatrizz[66][167] = 9'b111110011;
assign micromatrizz[66][168] = 9'b111111111;
assign micromatrizz[66][169] = 9'b111111111;
assign micromatrizz[66][170] = 9'b111111111;
assign micromatrizz[66][171] = 9'b111111111;
assign micromatrizz[66][172] = 9'b111110010;
assign micromatrizz[66][173] = 9'b111110010;
assign micromatrizz[66][174] = 9'b111110011;
assign micromatrizz[66][175] = 9'b111110011;
assign micromatrizz[66][176] = 9'b111110011;
assign micromatrizz[66][177] = 9'b111110011;
assign micromatrizz[66][178] = 9'b111110010;
assign micromatrizz[66][179] = 9'b111110111;
assign micromatrizz[66][180] = 9'b111111111;
assign micromatrizz[66][181] = 9'b111111111;
assign micromatrizz[66][182] = 9'b111111111;
assign micromatrizz[66][183] = 9'b111111111;
assign micromatrizz[66][184] = 9'b111110010;
assign micromatrizz[66][185] = 9'b111110010;
assign micromatrizz[66][186] = 9'b111110010;
assign micromatrizz[66][187] = 9'b111110010;
assign micromatrizz[66][188] = 9'b111110011;
assign micromatrizz[66][189] = 9'b111110011;
assign micromatrizz[66][190] = 9'b111110111;
assign micromatrizz[66][191] = 9'b111111111;
assign micromatrizz[66][192] = 9'b111111111;
assign micromatrizz[66][193] = 9'b111111111;
assign micromatrizz[66][194] = 9'b111110111;
assign micromatrizz[66][195] = 9'b111110010;
assign micromatrizz[66][196] = 9'b111110010;
assign micromatrizz[66][197] = 9'b111110011;
assign micromatrizz[66][198] = 9'b111110011;
assign micromatrizz[66][199] = 9'b111110010;
assign micromatrizz[66][200] = 9'b111110010;
assign micromatrizz[66][201] = 9'b111110011;
assign micromatrizz[66][202] = 9'b111110111;
assign micromatrizz[66][203] = 9'b111111111;
assign micromatrizz[66][204] = 9'b111111111;
assign micromatrizz[66][205] = 9'b111111111;
assign micromatrizz[66][206] = 9'b111111111;
assign micromatrizz[66][207] = 9'b111110111;
assign micromatrizz[66][208] = 9'b111110010;
assign micromatrizz[66][209] = 9'b111110010;
assign micromatrizz[66][210] = 9'b111110011;
assign micromatrizz[66][211] = 9'b111110011;
assign micromatrizz[66][212] = 9'b111110011;
assign micromatrizz[66][213] = 9'b111110111;
assign micromatrizz[66][214] = 9'b111111111;
assign micromatrizz[66][215] = 9'b111111111;
assign micromatrizz[66][216] = 9'b111111111;
assign micromatrizz[66][217] = 9'b111111111;
assign micromatrizz[66][218] = 9'b111111111;
assign micromatrizz[66][219] = 9'b111111111;
assign micromatrizz[66][220] = 9'b111110111;
assign micromatrizz[66][221] = 9'b111111111;
assign micromatrizz[66][222] = 9'b111111111;
assign micromatrizz[66][223] = 9'b111111111;
assign micromatrizz[66][224] = 9'b111111111;
assign micromatrizz[66][225] = 9'b111110011;
assign micromatrizz[66][226] = 9'b111110010;
assign micromatrizz[66][227] = 9'b111110010;
assign micromatrizz[66][228] = 9'b111110010;
assign micromatrizz[66][229] = 9'b111110011;
assign micromatrizz[66][230] = 9'b111110011;
assign micromatrizz[66][231] = 9'b111110011;
assign micromatrizz[66][232] = 9'b111110111;
assign micromatrizz[66][233] = 9'b111111111;
assign micromatrizz[66][234] = 9'b111111111;
assign micromatrizz[66][235] = 9'b111111111;
assign micromatrizz[66][236] = 9'b111111111;
assign micromatrizz[66][237] = 9'b111111111;
assign micromatrizz[66][238] = 9'b111111111;
assign micromatrizz[66][239] = 9'b111111111;
assign micromatrizz[66][240] = 9'b111111111;
assign micromatrizz[66][241] = 9'b111111111;
assign micromatrizz[66][242] = 9'b111110111;
assign micromatrizz[66][243] = 9'b111110010;
assign micromatrizz[66][244] = 9'b111110010;
assign micromatrizz[66][245] = 9'b111110010;
assign micromatrizz[66][246] = 9'b111110010;
assign micromatrizz[66][247] = 9'b111110111;
assign micromatrizz[66][248] = 9'b111111111;
assign micromatrizz[66][249] = 9'b111111111;
assign micromatrizz[66][250] = 9'b111111111;
assign micromatrizz[66][251] = 9'b111111111;
assign micromatrizz[66][252] = 9'b111111111;
assign micromatrizz[66][253] = 9'b111111111;
assign micromatrizz[66][254] = 9'b111111111;
assign micromatrizz[66][255] = 9'b111110010;
assign micromatrizz[66][256] = 9'b111110111;
assign micromatrizz[66][257] = 9'b111111111;
assign micromatrizz[66][258] = 9'b111111111;
assign micromatrizz[66][259] = 9'b111111111;
assign micromatrizz[66][260] = 9'b111111111;
assign micromatrizz[66][261] = 9'b111111111;
assign micromatrizz[66][262] = 9'b111111111;
assign micromatrizz[66][263] = 9'b111111111;
assign micromatrizz[66][264] = 9'b111111111;
assign micromatrizz[66][265] = 9'b111110111;
assign micromatrizz[66][266] = 9'b111110010;
assign micromatrizz[66][267] = 9'b111110011;
assign micromatrizz[66][268] = 9'b111110011;
assign micromatrizz[66][269] = 9'b111110011;
assign micromatrizz[66][270] = 9'b111110011;
assign micromatrizz[66][271] = 9'b111110010;
assign micromatrizz[66][272] = 9'b111111111;
assign micromatrizz[66][273] = 9'b111111111;
assign micromatrizz[66][274] = 9'b111111111;
assign micromatrizz[66][275] = 9'b111110010;
assign micromatrizz[66][276] = 9'b111110010;
assign micromatrizz[66][277] = 9'b111110011;
assign micromatrizz[66][278] = 9'b111110011;
assign micromatrizz[66][279] = 9'b111110011;
assign micromatrizz[66][280] = 9'b111110011;
assign micromatrizz[66][281] = 9'b111110011;
assign micromatrizz[66][282] = 9'b111111111;
assign micromatrizz[66][283] = 9'b111111111;
assign micromatrizz[66][284] = 9'b111111111;
assign micromatrizz[66][285] = 9'b111111111;
assign micromatrizz[66][286] = 9'b111110010;
assign micromatrizz[66][287] = 9'b111110010;
assign micromatrizz[66][288] = 9'b111110011;
assign micromatrizz[66][289] = 9'b111110011;
assign micromatrizz[66][290] = 9'b111110011;
assign micromatrizz[66][291] = 9'b111110011;
assign micromatrizz[66][292] = 9'b111110011;
assign micromatrizz[66][293] = 9'b111110111;
assign micromatrizz[66][294] = 9'b111111111;
assign micromatrizz[66][295] = 9'b111111111;
assign micromatrizz[66][296] = 9'b111111111;
assign micromatrizz[66][297] = 9'b111111111;
assign micromatrizz[66][298] = 9'b111111111;
assign micromatrizz[66][299] = 9'b111111111;
assign micromatrizz[66][300] = 9'b111111111;
assign micromatrizz[66][301] = 9'b111111111;
assign micromatrizz[66][302] = 9'b111111111;
assign micromatrizz[66][303] = 9'b111110111;
assign micromatrizz[66][304] = 9'b111110010;
assign micromatrizz[66][305] = 9'b111110011;
assign micromatrizz[66][306] = 9'b111110011;
assign micromatrizz[66][307] = 9'b111110111;
assign micromatrizz[66][308] = 9'b111111111;
assign micromatrizz[66][309] = 9'b111111111;
assign micromatrizz[66][310] = 9'b111111111;
assign micromatrizz[66][311] = 9'b111111111;
assign micromatrizz[66][312] = 9'b111111111;
assign micromatrizz[66][313] = 9'b111111111;
assign micromatrizz[66][314] = 9'b111111111;
assign micromatrizz[66][315] = 9'b111111111;
assign micromatrizz[66][316] = 9'b111111111;
assign micromatrizz[66][317] = 9'b111110010;
assign micromatrizz[66][318] = 9'b111110010;
assign micromatrizz[66][319] = 9'b111110011;
assign micromatrizz[66][320] = 9'b111110011;
assign micromatrizz[66][321] = 9'b111110011;
assign micromatrizz[66][322] = 9'b111111111;
assign micromatrizz[66][323] = 9'b111111111;
assign micromatrizz[66][324] = 9'b111111111;
assign micromatrizz[66][325] = 9'b111111111;
assign micromatrizz[66][326] = 9'b111111111;
assign micromatrizz[66][327] = 9'b111111111;
assign micromatrizz[66][328] = 9'b111111111;
assign micromatrizz[66][329] = 9'b111110111;
assign micromatrizz[66][330] = 9'b111110010;
assign micromatrizz[66][331] = 9'b111111111;
assign micromatrizz[66][332] = 9'b111111111;
assign micromatrizz[66][333] = 9'b111111111;
assign micromatrizz[66][334] = 9'b111111111;
assign micromatrizz[66][335] = 9'b111110010;
assign micromatrizz[66][336] = 9'b111110011;
assign micromatrizz[66][337] = 9'b111110011;
assign micromatrizz[66][338] = 9'b111110011;
assign micromatrizz[66][339] = 9'b111110010;
assign micromatrizz[66][340] = 9'b111110010;
assign micromatrizz[66][341] = 9'b111110010;
assign micromatrizz[66][342] = 9'b111111111;
assign micromatrizz[66][343] = 9'b111111111;
assign micromatrizz[66][344] = 9'b111111111;
assign micromatrizz[66][345] = 9'b111111111;
assign micromatrizz[66][346] = 9'b111111111;
assign micromatrizz[66][347] = 9'b111110010;
assign micromatrizz[66][348] = 9'b111110010;
assign micromatrizz[66][349] = 9'b111110010;
assign micromatrizz[66][350] = 9'b111110010;
assign micromatrizz[66][351] = 9'b111110010;
assign micromatrizz[66][352] = 9'b111110011;
assign micromatrizz[66][353] = 9'b111110011;
assign micromatrizz[66][354] = 9'b111111111;
assign micromatrizz[66][355] = 9'b111111111;
assign micromatrizz[66][356] = 9'b111111111;
assign micromatrizz[66][357] = 9'b111111111;
assign micromatrizz[66][358] = 9'b111111111;
assign micromatrizz[66][359] = 9'b111110010;
assign micromatrizz[66][360] = 9'b111110011;
assign micromatrizz[66][361] = 9'b111110010;
assign micromatrizz[66][362] = 9'b111110010;
assign micromatrizz[66][363] = 9'b111110010;
assign micromatrizz[66][364] = 9'b111110010;
assign micromatrizz[66][365] = 9'b111110011;
assign micromatrizz[66][366] = 9'b111111111;
assign micromatrizz[66][367] = 9'b111111111;
assign micromatrizz[66][368] = 9'b111111111;
assign micromatrizz[66][369] = 9'b111110010;
assign micromatrizz[66][370] = 9'b111111111;
assign micromatrizz[66][371] = 9'b111111111;
assign micromatrizz[66][372] = 9'b111110010;
assign micromatrizz[66][373] = 9'b111110011;
assign micromatrizz[66][374] = 9'b111110011;
assign micromatrizz[66][375] = 9'b111110011;
assign micromatrizz[66][376] = 9'b111110011;
assign micromatrizz[66][377] = 9'b111110010;
assign micromatrizz[66][378] = 9'b111110010;
assign micromatrizz[66][379] = 9'b111111111;
assign micromatrizz[66][380] = 9'b111111111;
assign micromatrizz[66][381] = 9'b111111111;
assign micromatrizz[66][382] = 9'b111111111;
assign micromatrizz[66][383] = 9'b111110111;
assign micromatrizz[66][384] = 9'b111110010;
assign micromatrizz[66][385] = 9'b111110010;
assign micromatrizz[66][386] = 9'b111110011;
assign micromatrizz[66][387] = 9'b111110011;
assign micromatrizz[66][388] = 9'b111110011;
assign micromatrizz[66][389] = 9'b111110011;
assign micromatrizz[66][390] = 9'b111110011;
assign micromatrizz[66][391] = 9'b111111111;
assign micromatrizz[66][392] = 9'b111111111;
assign micromatrizz[66][393] = 9'b111111111;
assign micromatrizz[66][394] = 9'b111111111;
assign micromatrizz[66][395] = 9'b111110010;
assign micromatrizz[66][396] = 9'b111110010;
assign micromatrizz[66][397] = 9'b111110010;
assign micromatrizz[66][398] = 9'b111110010;
assign micromatrizz[66][399] = 9'b111110011;
assign micromatrizz[66][400] = 9'b111110011;
assign micromatrizz[66][401] = 9'b111110011;
assign micromatrizz[66][402] = 9'b111110111;
assign micromatrizz[66][403] = 9'b111111111;
assign micromatrizz[66][404] = 9'b111111111;
assign micromatrizz[66][405] = 9'b111111111;
assign micromatrizz[66][406] = 9'b111111111;
assign micromatrizz[66][407] = 9'b111111111;
assign micromatrizz[66][408] = 9'b111111111;
assign micromatrizz[66][409] = 9'b111111111;
assign micromatrizz[66][410] = 9'b111111111;
assign micromatrizz[66][411] = 9'b111111111;
assign micromatrizz[66][412] = 9'b111110111;
assign micromatrizz[66][413] = 9'b111110010;
assign micromatrizz[66][414] = 9'b111110010;
assign micromatrizz[66][415] = 9'b111110011;
assign micromatrizz[66][416] = 9'b111110011;
assign micromatrizz[66][417] = 9'b111110111;
assign micromatrizz[66][418] = 9'b111111111;
assign micromatrizz[66][419] = 9'b111111111;
assign micromatrizz[66][420] = 9'b111111111;
assign micromatrizz[66][421] = 9'b111111111;
assign micromatrizz[66][422] = 9'b111111111;
assign micromatrizz[66][423] = 9'b111111111;
assign micromatrizz[66][424] = 9'b111111111;
assign micromatrizz[66][425] = 9'b111110010;
assign micromatrizz[66][426] = 9'b111110111;
assign micromatrizz[66][427] = 9'b111111111;
assign micromatrizz[66][428] = 9'b111111111;
assign micromatrizz[66][429] = 9'b111111111;
assign micromatrizz[66][430] = 9'b111110111;
assign micromatrizz[66][431] = 9'b111110010;
assign micromatrizz[66][432] = 9'b111110010;
assign micromatrizz[66][433] = 9'b111110010;
assign micromatrizz[66][434] = 9'b111110010;
assign micromatrizz[66][435] = 9'b111110011;
assign micromatrizz[66][436] = 9'b111110011;
assign micromatrizz[66][437] = 9'b111110011;
assign micromatrizz[66][438] = 9'b111111111;
assign micromatrizz[66][439] = 9'b111111111;
assign micromatrizz[66][440] = 9'b111111111;
assign micromatrizz[66][441] = 9'b111111111;
assign micromatrizz[66][442] = 9'b111111111;
assign micromatrizz[66][443] = 9'b111111111;
assign micromatrizz[66][444] = 9'b111111111;
assign micromatrizz[66][445] = 9'b111111111;
assign micromatrizz[66][446] = 9'b111111111;
assign micromatrizz[66][447] = 9'b111111111;
assign micromatrizz[66][448] = 9'b111110010;
assign micromatrizz[66][449] = 9'b111110010;
assign micromatrizz[66][450] = 9'b111110010;
assign micromatrizz[66][451] = 9'b111110011;
assign micromatrizz[66][452] = 9'b111110011;
assign micromatrizz[66][453] = 9'b111110011;
assign micromatrizz[66][454] = 9'b111111111;
assign micromatrizz[66][455] = 9'b111111111;
assign micromatrizz[66][456] = 9'b111111111;
assign micromatrizz[66][457] = 9'b111111111;
assign micromatrizz[66][458] = 9'b111111111;
assign micromatrizz[66][459] = 9'b111111111;
assign micromatrizz[66][460] = 9'b111110110;
assign micromatrizz[66][461] = 9'b111111111;
assign micromatrizz[66][462] = 9'b111111111;
assign micromatrizz[66][463] = 9'b111111111;
assign micromatrizz[66][464] = 9'b111111111;
assign micromatrizz[66][465] = 9'b111111111;
assign micromatrizz[66][466] = 9'b111111111;
assign micromatrizz[66][467] = 9'b111111111;
assign micromatrizz[66][468] = 9'b111111111;
assign micromatrizz[66][469] = 9'b111111111;
assign micromatrizz[66][470] = 9'b111111111;
assign micromatrizz[66][471] = 9'b111110010;
assign micromatrizz[66][472] = 9'b111110010;
assign micromatrizz[66][473] = 9'b111110011;
assign micromatrizz[66][474] = 9'b111110010;
assign micromatrizz[66][475] = 9'b111110011;
assign micromatrizz[66][476] = 9'b111110011;
assign micromatrizz[66][477] = 9'b111110111;
assign micromatrizz[66][478] = 9'b111111111;
assign micromatrizz[66][479] = 9'b111111111;
assign micromatrizz[66][480] = 9'b111111111;
assign micromatrizz[66][481] = 9'b111110010;
assign micromatrizz[66][482] = 9'b111110010;
assign micromatrizz[66][483] = 9'b111110010;
assign micromatrizz[66][484] = 9'b111110010;
assign micromatrizz[66][485] = 9'b111110011;
assign micromatrizz[66][486] = 9'b111110011;
assign micromatrizz[66][487] = 9'b111110011;
assign micromatrizz[66][488] = 9'b111110111;
assign micromatrizz[66][489] = 9'b111111111;
assign micromatrizz[66][490] = 9'b111111111;
assign micromatrizz[66][491] = 9'b111111111;
assign micromatrizz[66][492] = 9'b111111111;
assign micromatrizz[66][493] = 9'b111111111;
assign micromatrizz[66][494] = 9'b111111111;
assign micromatrizz[66][495] = 9'b111111111;
assign micromatrizz[66][496] = 9'b111111111;
assign micromatrizz[66][497] = 9'b111111111;
assign micromatrizz[66][498] = 9'b111110111;
assign micromatrizz[66][499] = 9'b111110010;
assign micromatrizz[66][500] = 9'b111110010;
assign micromatrizz[66][501] = 9'b111110010;
assign micromatrizz[66][502] = 9'b111110010;
assign micromatrizz[66][503] = 9'b111111111;
assign micromatrizz[66][504] = 9'b111111111;
assign micromatrizz[66][505] = 9'b111111111;
assign micromatrizz[66][506] = 9'b111111111;
assign micromatrizz[66][507] = 9'b111111111;
assign micromatrizz[66][508] = 9'b111111111;
assign micromatrizz[66][509] = 9'b111111111;
assign micromatrizz[66][510] = 9'b111111111;
assign micromatrizz[66][511] = 9'b111110010;
assign micromatrizz[66][512] = 9'b111110111;
assign micromatrizz[66][513] = 9'b111111111;
assign micromatrizz[66][514] = 9'b111111111;
assign micromatrizz[66][515] = 9'b111111111;
assign micromatrizz[66][516] = 9'b111110111;
assign micromatrizz[66][517] = 9'b111110010;
assign micromatrizz[66][518] = 9'b111110011;
assign micromatrizz[66][519] = 9'b111110011;
assign micromatrizz[66][520] = 9'b111110010;
assign micromatrizz[66][521] = 9'b111110010;
assign micromatrizz[66][522] = 9'b111110011;
assign micromatrizz[66][523] = 9'b111110011;
assign micromatrizz[66][524] = 9'b111111111;
assign micromatrizz[66][525] = 9'b111111111;
assign micromatrizz[66][526] = 9'b111111111;
assign micromatrizz[66][527] = 9'b111111111;
assign micromatrizz[66][528] = 9'b111111111;
assign micromatrizz[66][529] = 9'b111110010;
assign micromatrizz[66][530] = 9'b111110010;
assign micromatrizz[66][531] = 9'b111110010;
assign micromatrizz[66][532] = 9'b111110011;
assign micromatrizz[66][533] = 9'b111110011;
assign micromatrizz[66][534] = 9'b111110011;
assign micromatrizz[66][535] = 9'b111111111;
assign micromatrizz[66][536] = 9'b111111111;
assign micromatrizz[66][537] = 9'b111111111;
assign micromatrizz[66][538] = 9'b111111111;
assign micromatrizz[66][539] = 9'b111111111;
assign micromatrizz[66][540] = 9'b111110010;
assign micromatrizz[66][541] = 9'b111110010;
assign micromatrizz[66][542] = 9'b111110011;
assign micromatrizz[66][543] = 9'b111110010;
assign micromatrizz[66][544] = 9'b111110011;
assign micromatrizz[66][545] = 9'b111111111;
assign micromatrizz[66][546] = 9'b111111111;
assign micromatrizz[66][547] = 9'b111111111;
assign micromatrizz[66][548] = 9'b111111111;
assign micromatrizz[66][549] = 9'b111111111;
assign micromatrizz[66][550] = 9'b111111111;
assign micromatrizz[66][551] = 9'b111111111;
assign micromatrizz[66][552] = 9'b111110111;
assign micromatrizz[66][553] = 9'b111110010;
assign micromatrizz[66][554] = 9'b111111111;
assign micromatrizz[66][555] = 9'b111111111;
assign micromatrizz[66][556] = 9'b111111111;
assign micromatrizz[66][557] = 9'b111111111;
assign micromatrizz[66][558] = 9'b111110010;
assign micromatrizz[66][559] = 9'b111110010;
assign micromatrizz[66][560] = 9'b111110010;
assign micromatrizz[66][561] = 9'b111110010;
assign micromatrizz[66][562] = 9'b111110011;
assign micromatrizz[66][563] = 9'b111110011;
assign micromatrizz[66][564] = 9'b111110010;
assign micromatrizz[66][565] = 9'b111111111;
assign micromatrizz[66][566] = 9'b111111111;
assign micromatrizz[66][567] = 9'b111111111;
assign micromatrizz[66][568] = 9'b111111111;
assign micromatrizz[66][569] = 9'b111111111;
assign micromatrizz[66][570] = 9'b111110010;
assign micromatrizz[66][571] = 9'b111110010;
assign micromatrizz[66][572] = 9'b111110010;
assign micromatrizz[66][573] = 9'b111110010;
assign micromatrizz[66][574] = 9'b111110011;
assign micromatrizz[66][575] = 9'b111110011;
assign micromatrizz[66][576] = 9'b111111111;
assign micromatrizz[66][577] = 9'b111111111;
assign micromatrizz[66][578] = 9'b111111111;
assign micromatrizz[66][579] = 9'b111111111;
assign micromatrizz[66][580] = 9'b111110111;
assign micromatrizz[66][581] = 9'b111110010;
assign micromatrizz[66][582] = 9'b111110010;
assign micromatrizz[66][583] = 9'b111110011;
assign micromatrizz[66][584] = 9'b111110011;
assign micromatrizz[66][585] = 9'b111110011;
assign micromatrizz[66][586] = 9'b111110011;
assign micromatrizz[66][587] = 9'b111110011;
assign micromatrizz[66][588] = 9'b111111111;
assign micromatrizz[66][589] = 9'b111111111;
assign micromatrizz[66][590] = 9'b111111111;
assign micromatrizz[66][591] = 9'b111111111;
assign micromatrizz[66][592] = 9'b111111111;
assign micromatrizz[66][593] = 9'b111110010;
assign micromatrizz[66][594] = 9'b111110010;
assign micromatrizz[66][595] = 9'b111110011;
assign micromatrizz[66][596] = 9'b111110011;
assign micromatrizz[66][597] = 9'b111110011;
assign micromatrizz[66][598] = 9'b111111111;
assign micromatrizz[66][599] = 9'b111111111;
assign micromatrizz[66][600] = 9'b111111111;
assign micromatrizz[66][601] = 9'b111111111;
assign micromatrizz[66][602] = 9'b111111111;
assign micromatrizz[66][603] = 9'b111111111;
assign micromatrizz[66][604] = 9'b111111111;
assign micromatrizz[66][605] = 9'b111110111;
assign micromatrizz[66][606] = 9'b111110010;
assign micromatrizz[66][607] = 9'b111111111;
assign micromatrizz[66][608] = 9'b111111111;
assign micromatrizz[66][609] = 9'b111111111;
assign micromatrizz[66][610] = 9'b111111111;
assign micromatrizz[66][611] = 9'b111111111;
assign micromatrizz[66][612] = 9'b111111111;
assign micromatrizz[66][613] = 9'b111111111;
assign micromatrizz[66][614] = 9'b111111111;
assign micromatrizz[66][615] = 9'b111111111;
assign micromatrizz[66][616] = 9'b111110111;
assign micromatrizz[66][617] = 9'b111110010;
assign micromatrizz[66][618] = 9'b111110010;
assign micromatrizz[66][619] = 9'b111110010;
assign micromatrizz[66][620] = 9'b111110011;
assign micromatrizz[66][621] = 9'b111110011;
assign micromatrizz[66][622] = 9'b111110111;
assign micromatrizz[66][623] = 9'b111111111;
assign micromatrizz[66][624] = 9'b111111111;
assign micromatrizz[66][625] = 9'b111111111;
assign micromatrizz[66][626] = 9'b111111111;
assign micromatrizz[66][627] = 9'b111111111;
assign micromatrizz[66][628] = 9'b111111111;
assign micromatrizz[66][629] = 9'b111111111;
assign micromatrizz[66][630] = 9'b111111111;
assign micromatrizz[66][631] = 9'b111111111;
assign micromatrizz[66][632] = 9'b111111111;
assign micromatrizz[66][633] = 9'b111111111;
assign micromatrizz[66][634] = 9'b111111111;
assign micromatrizz[66][635] = 9'b111111111;
assign micromatrizz[66][636] = 9'b111111111;
assign micromatrizz[66][637] = 9'b111111111;
assign micromatrizz[66][638] = 9'b111111111;
assign micromatrizz[66][639] = 9'b111111111;
assign micromatrizz[67][0] = 9'b111111111;
assign micromatrizz[67][1] = 9'b111111111;
assign micromatrizz[67][2] = 9'b111111111;
assign micromatrizz[67][3] = 9'b111111111;
assign micromatrizz[67][4] = 9'b111111111;
assign micromatrizz[67][5] = 9'b111111111;
assign micromatrizz[67][6] = 9'b111111111;
assign micromatrizz[67][7] = 9'b111111111;
assign micromatrizz[67][8] = 9'b111110010;
assign micromatrizz[67][9] = 9'b111111111;
assign micromatrizz[67][10] = 9'b111111111;
assign micromatrizz[67][11] = 9'b111111111;
assign micromatrizz[67][12] = 9'b111111111;
assign micromatrizz[67][13] = 9'b111111111;
assign micromatrizz[67][14] = 9'b111110111;
assign micromatrizz[67][15] = 9'b111110010;
assign micromatrizz[67][16] = 9'b111110011;
assign micromatrizz[67][17] = 9'b111110011;
assign micromatrizz[67][18] = 9'b111110011;
assign micromatrizz[67][19] = 9'b111110010;
assign micromatrizz[67][20] = 9'b111111111;
assign micromatrizz[67][21] = 9'b111111111;
assign micromatrizz[67][22] = 9'b111111111;
assign micromatrizz[67][23] = 9'b111111111;
assign micromatrizz[67][24] = 9'b111110010;
assign micromatrizz[67][25] = 9'b111110010;
assign micromatrizz[67][26] = 9'b111110010;
assign micromatrizz[67][27] = 9'b111110011;
assign micromatrizz[67][28] = 9'b111110011;
assign micromatrizz[67][29] = 9'b111110011;
assign micromatrizz[67][30] = 9'b111110011;
assign micromatrizz[67][31] = 9'b111111111;
assign micromatrizz[67][32] = 9'b111111111;
assign micromatrizz[67][33] = 9'b111111111;
assign micromatrizz[67][34] = 9'b111110111;
assign micromatrizz[67][35] = 9'b111110010;
assign micromatrizz[67][36] = 9'b111110010;
assign micromatrizz[67][37] = 9'b111110011;
assign micromatrizz[67][38] = 9'b111110011;
assign micromatrizz[67][39] = 9'b111110010;
assign micromatrizz[67][40] = 9'b111110011;
assign micromatrizz[67][41] = 9'b111110011;
assign micromatrizz[67][42] = 9'b111110010;
assign micromatrizz[67][43] = 9'b111111111;
assign micromatrizz[67][44] = 9'b111111111;
assign micromatrizz[67][45] = 9'b111111111;
assign micromatrizz[67][46] = 9'b111111111;
assign micromatrizz[67][47] = 9'b111110010;
assign micromatrizz[67][48] = 9'b111110010;
assign micromatrizz[67][49] = 9'b111110011;
assign micromatrizz[67][50] = 9'b111110011;
assign micromatrizz[67][51] = 9'b111110011;
assign micromatrizz[67][52] = 9'b111110010;
assign micromatrizz[67][53] = 9'b111110010;
assign micromatrizz[67][54] = 9'b111111111;
assign micromatrizz[67][55] = 9'b111111111;
assign micromatrizz[67][56] = 9'b111111111;
assign micromatrizz[67][57] = 9'b111110111;
assign micromatrizz[67][58] = 9'b111110010;
assign micromatrizz[67][59] = 9'b111110010;
assign micromatrizz[67][60] = 9'b111110010;
assign micromatrizz[67][61] = 9'b111110010;
assign micromatrizz[67][62] = 9'b111110111;
assign micromatrizz[67][63] = 9'b111111111;
assign micromatrizz[67][64] = 9'b111111111;
assign micromatrizz[67][65] = 9'b111111111;
assign micromatrizz[67][66] = 9'b111111111;
assign micromatrizz[67][67] = 9'b111111111;
assign micromatrizz[67][68] = 9'b111111111;
assign micromatrizz[67][69] = 9'b111111111;
assign micromatrizz[67][70] = 9'b111111111;
assign micromatrizz[67][71] = 9'b111110010;
assign micromatrizz[67][72] = 9'b111110010;
assign micromatrizz[67][73] = 9'b111110010;
assign micromatrizz[67][74] = 9'b111110011;
assign micromatrizz[67][75] = 9'b111111111;
assign micromatrizz[67][76] = 9'b111111111;
assign micromatrizz[67][77] = 9'b111111111;
assign micromatrizz[67][78] = 9'b111111111;
assign micromatrizz[67][79] = 9'b111111111;
assign micromatrizz[67][80] = 9'b111111111;
assign micromatrizz[67][81] = 9'b111110111;
assign micromatrizz[67][82] = 9'b111110010;
assign micromatrizz[67][83] = 9'b111110111;
assign micromatrizz[67][84] = 9'b111111111;
assign micromatrizz[67][85] = 9'b111111111;
assign micromatrizz[67][86] = 9'b111111111;
assign micromatrizz[67][87] = 9'b111111111;
assign micromatrizz[67][88] = 9'b111110010;
assign micromatrizz[67][89] = 9'b111110010;
assign micromatrizz[67][90] = 9'b111110011;
assign micromatrizz[67][91] = 9'b111110011;
assign micromatrizz[67][92] = 9'b111110011;
assign micromatrizz[67][93] = 9'b111110011;
assign micromatrizz[67][94] = 9'b111110010;
assign micromatrizz[67][95] = 9'b111110111;
assign micromatrizz[67][96] = 9'b111111111;
assign micromatrizz[67][97] = 9'b111111111;
assign micromatrizz[67][98] = 9'b111111111;
assign micromatrizz[67][99] = 9'b111111111;
assign micromatrizz[67][100] = 9'b111111111;
assign micromatrizz[67][101] = 9'b111111111;
assign micromatrizz[67][102] = 9'b111111111;
assign micromatrizz[67][103] = 9'b111111111;
assign micromatrizz[67][104] = 9'b111110010;
assign micromatrizz[67][105] = 9'b111110111;
assign micromatrizz[67][106] = 9'b111111111;
assign micromatrizz[67][107] = 9'b111111111;
assign micromatrizz[67][108] = 9'b111111111;
assign micromatrizz[67][109] = 9'b111111111;
assign micromatrizz[67][110] = 9'b111111111;
assign micromatrizz[67][111] = 9'b111110010;
assign micromatrizz[67][112] = 9'b111110011;
assign micromatrizz[67][113] = 9'b111110011;
assign micromatrizz[67][114] = 9'b111110011;
assign micromatrizz[67][115] = 9'b111110010;
assign micromatrizz[67][116] = 9'b111111111;
assign micromatrizz[67][117] = 9'b111111111;
assign micromatrizz[67][118] = 9'b111111111;
assign micromatrizz[67][119] = 9'b111111111;
assign micromatrizz[67][120] = 9'b111111111;
assign micromatrizz[67][121] = 9'b111110111;
assign micromatrizz[67][122] = 9'b111110010;
assign micromatrizz[67][123] = 9'b111110011;
assign micromatrizz[67][124] = 9'b111110010;
assign micromatrizz[67][125] = 9'b111110011;
assign micromatrizz[67][126] = 9'b111110111;
assign micromatrizz[67][127] = 9'b111111111;
assign micromatrizz[67][128] = 9'b111111111;
assign micromatrizz[67][129] = 9'b111111111;
assign micromatrizz[67][130] = 9'b111111111;
assign micromatrizz[67][131] = 9'b111111111;
assign micromatrizz[67][132] = 9'b111110111;
assign micromatrizz[67][133] = 9'b111111111;
assign micromatrizz[67][134] = 9'b111111111;
assign micromatrizz[67][135] = 9'b111111111;
assign micromatrizz[67][136] = 9'b111111111;
assign micromatrizz[67][137] = 9'b111111111;
assign micromatrizz[67][138] = 9'b111110111;
assign micromatrizz[67][139] = 9'b111110010;
assign micromatrizz[67][140] = 9'b111110010;
assign micromatrizz[67][141] = 9'b111110010;
assign micromatrizz[67][142] = 9'b111110010;
assign micromatrizz[67][143] = 9'b111110010;
assign micromatrizz[67][144] = 9'b111110011;
assign micromatrizz[67][145] = 9'b111110111;
assign micromatrizz[67][146] = 9'b111111111;
assign micromatrizz[67][147] = 9'b111111111;
assign micromatrizz[67][148] = 9'b111111111;
assign micromatrizz[67][149] = 9'b111111111;
assign micromatrizz[67][150] = 9'b111110111;
assign micromatrizz[67][151] = 9'b111110010;
assign micromatrizz[67][152] = 9'b111110010;
assign micromatrizz[67][153] = 9'b111110010;
assign micromatrizz[67][154] = 9'b111110011;
assign micromatrizz[67][155] = 9'b111110011;
assign micromatrizz[67][156] = 9'b111110011;
assign micromatrizz[67][157] = 9'b111110111;
assign micromatrizz[67][158] = 9'b111111111;
assign micromatrizz[67][159] = 9'b111111111;
assign micromatrizz[67][160] = 9'b111111111;
assign micromatrizz[67][161] = 9'b111111111;
assign micromatrizz[67][162] = 9'b111110010;
assign micromatrizz[67][163] = 9'b111110010;
assign micromatrizz[67][164] = 9'b111110011;
assign micromatrizz[67][165] = 9'b111110011;
assign micromatrizz[67][166] = 9'b111110011;
assign micromatrizz[67][167] = 9'b111110010;
assign micromatrizz[67][168] = 9'b111111111;
assign micromatrizz[67][169] = 9'b111111111;
assign micromatrizz[67][170] = 9'b111111111;
assign micromatrizz[67][171] = 9'b111110111;
assign micromatrizz[67][172] = 9'b111110010;
assign micromatrizz[67][173] = 9'b111110011;
assign micromatrizz[67][174] = 9'b111110011;
assign micromatrizz[67][175] = 9'b111110011;
assign micromatrizz[67][176] = 9'b111110011;
assign micromatrizz[67][177] = 9'b111110011;
assign micromatrizz[67][178] = 9'b111110010;
assign micromatrizz[67][179] = 9'b111110111;
assign micromatrizz[67][180] = 9'b111111111;
assign micromatrizz[67][181] = 9'b111111111;
assign micromatrizz[67][182] = 9'b111111111;
assign micromatrizz[67][183] = 9'b111111111;
assign micromatrizz[67][184] = 9'b111111111;
assign micromatrizz[67][185] = 9'b111110010;
assign micromatrizz[67][186] = 9'b111110010;
assign micromatrizz[67][187] = 9'b111110011;
assign micromatrizz[67][188] = 9'b111110011;
assign micromatrizz[67][189] = 9'b111110011;
assign micromatrizz[67][190] = 9'b111110111;
assign micromatrizz[67][191] = 9'b111111111;
assign micromatrizz[67][192] = 9'b111111111;
assign micromatrizz[67][193] = 9'b111110111;
assign micromatrizz[67][194] = 9'b111110010;
assign micromatrizz[67][195] = 9'b111110010;
assign micromatrizz[67][196] = 9'b111110011;
assign micromatrizz[67][197] = 9'b111110011;
assign micromatrizz[67][198] = 9'b111110011;
assign micromatrizz[67][199] = 9'b111110010;
assign micromatrizz[67][200] = 9'b111110010;
assign micromatrizz[67][201] = 9'b111110011;
assign micromatrizz[67][202] = 9'b111110111;
assign micromatrizz[67][203] = 9'b111111111;
assign micromatrizz[67][204] = 9'b111111111;
assign micromatrizz[67][205] = 9'b111111111;
assign micromatrizz[67][206] = 9'b111111111;
assign micromatrizz[67][207] = 9'b111111111;
assign micromatrizz[67][208] = 9'b111110010;
assign micromatrizz[67][209] = 9'b111110010;
assign micromatrizz[67][210] = 9'b111110010;
assign micromatrizz[67][211] = 9'b111110011;
assign micromatrizz[67][212] = 9'b111110011;
assign micromatrizz[67][213] = 9'b111110111;
assign micromatrizz[67][214] = 9'b111111111;
assign micromatrizz[67][215] = 9'b111111111;
assign micromatrizz[67][216] = 9'b111111111;
assign micromatrizz[67][217] = 9'b111111111;
assign micromatrizz[67][218] = 9'b111111111;
assign micromatrizz[67][219] = 9'b111110110;
assign micromatrizz[67][220] = 9'b111111111;
assign micromatrizz[67][221] = 9'b111111111;
assign micromatrizz[67][222] = 9'b111111111;
assign micromatrizz[67][223] = 9'b111111111;
assign micromatrizz[67][224] = 9'b111111111;
assign micromatrizz[67][225] = 9'b111110010;
assign micromatrizz[67][226] = 9'b111110010;
assign micromatrizz[67][227] = 9'b111110010;
assign micromatrizz[67][228] = 9'b111110010;
assign micromatrizz[67][229] = 9'b111110011;
assign micromatrizz[67][230] = 9'b111110011;
assign micromatrizz[67][231] = 9'b111110011;
assign micromatrizz[67][232] = 9'b111110111;
assign micromatrizz[67][233] = 9'b111111111;
assign micromatrizz[67][234] = 9'b111111111;
assign micromatrizz[67][235] = 9'b111111111;
assign micromatrizz[67][236] = 9'b111111111;
assign micromatrizz[67][237] = 9'b111111111;
assign micromatrizz[67][238] = 9'b111111111;
assign micromatrizz[67][239] = 9'b111111111;
assign micromatrizz[67][240] = 9'b111111111;
assign micromatrizz[67][241] = 9'b111111111;
assign micromatrizz[67][242] = 9'b111111111;
assign micromatrizz[67][243] = 9'b111110111;
assign micromatrizz[67][244] = 9'b111110010;
assign micromatrizz[67][245] = 9'b111110010;
assign micromatrizz[67][246] = 9'b111110010;
assign micromatrizz[67][247] = 9'b111110111;
assign micromatrizz[67][248] = 9'b111111111;
assign micromatrizz[67][249] = 9'b111111111;
assign micromatrizz[67][250] = 9'b111111111;
assign micromatrizz[67][251] = 9'b111111111;
assign micromatrizz[67][252] = 9'b111111111;
assign micromatrizz[67][253] = 9'b111111111;
assign micromatrizz[67][254] = 9'b111110010;
assign micromatrizz[67][255] = 9'b111110111;
assign micromatrizz[67][256] = 9'b111111111;
assign micromatrizz[67][257] = 9'b111111111;
assign micromatrizz[67][258] = 9'b111111111;
assign micromatrizz[67][259] = 9'b111110111;
assign micromatrizz[67][260] = 9'b111110010;
assign micromatrizz[67][261] = 9'b111111111;
assign micromatrizz[67][262] = 9'b111111111;
assign micromatrizz[67][263] = 9'b111111111;
assign micromatrizz[67][264] = 9'b111111111;
assign micromatrizz[67][265] = 9'b111111111;
assign micromatrizz[67][266] = 9'b111110111;
assign micromatrizz[67][267] = 9'b111110010;
assign micromatrizz[67][268] = 9'b111110011;
assign micromatrizz[67][269] = 9'b111110010;
assign micromatrizz[67][270] = 9'b111110010;
assign micromatrizz[67][271] = 9'b111110010;
assign micromatrizz[67][272] = 9'b111111111;
assign micromatrizz[67][273] = 9'b111111111;
assign micromatrizz[67][274] = 9'b111111111;
assign micromatrizz[67][275] = 9'b111110111;
assign micromatrizz[67][276] = 9'b111110010;
assign micromatrizz[67][277] = 9'b111110010;
assign micromatrizz[67][278] = 9'b111110011;
assign micromatrizz[67][279] = 9'b111110011;
assign micromatrizz[67][280] = 9'b111110011;
assign micromatrizz[67][281] = 9'b111110011;
assign micromatrizz[67][282] = 9'b111111111;
assign micromatrizz[67][283] = 9'b111111111;
assign micromatrizz[67][284] = 9'b111111111;
assign micromatrizz[67][285] = 9'b111110111;
assign micromatrizz[67][286] = 9'b111110011;
assign micromatrizz[67][287] = 9'b111110010;
assign micromatrizz[67][288] = 9'b111110010;
assign micromatrizz[67][289] = 9'b111110011;
assign micromatrizz[67][290] = 9'b111110011;
assign micromatrizz[67][291] = 9'b111110011;
assign micromatrizz[67][292] = 9'b111110011;
assign micromatrizz[67][293] = 9'b111111111;
assign micromatrizz[67][294] = 9'b111111111;
assign micromatrizz[67][295] = 9'b111111111;
assign micromatrizz[67][296] = 9'b111111111;
assign micromatrizz[67][297] = 9'b111111111;
assign micromatrizz[67][298] = 9'b111111111;
assign micromatrizz[67][299] = 9'b111111111;
assign micromatrizz[67][300] = 9'b111111111;
assign micromatrizz[67][301] = 9'b111111111;
assign micromatrizz[67][302] = 9'b111111111;
assign micromatrizz[67][303] = 9'b111111111;
assign micromatrizz[67][304] = 9'b111110010;
assign micromatrizz[67][305] = 9'b111110011;
assign micromatrizz[67][306] = 9'b111110010;
assign micromatrizz[67][307] = 9'b111111111;
assign micromatrizz[67][308] = 9'b111111111;
assign micromatrizz[67][309] = 9'b111111111;
assign micromatrizz[67][310] = 9'b111111111;
assign micromatrizz[67][311] = 9'b111111111;
assign micromatrizz[67][312] = 9'b111111111;
assign micromatrizz[67][313] = 9'b111111111;
assign micromatrizz[67][314] = 9'b111111111;
assign micromatrizz[67][315] = 9'b111111111;
assign micromatrizz[67][316] = 9'b111111111;
assign micromatrizz[67][317] = 9'b111111111;
assign micromatrizz[67][318] = 9'b111110010;
assign micromatrizz[67][319] = 9'b111110010;
assign micromatrizz[67][320] = 9'b111110010;
assign micromatrizz[67][321] = 9'b111110011;
assign micromatrizz[67][322] = 9'b111111111;
assign micromatrizz[67][323] = 9'b111111111;
assign micromatrizz[67][324] = 9'b111111111;
assign micromatrizz[67][325] = 9'b111111111;
assign micromatrizz[67][326] = 9'b111111111;
assign micromatrizz[67][327] = 9'b111111111;
assign micromatrizz[67][328] = 9'b111110111;
assign micromatrizz[67][329] = 9'b111110010;
assign micromatrizz[67][330] = 9'b111111111;
assign micromatrizz[67][331] = 9'b111111111;
assign micromatrizz[67][332] = 9'b111111111;
assign micromatrizz[67][333] = 9'b111111111;
assign micromatrizz[67][334] = 9'b111111111;
assign micromatrizz[67][335] = 9'b111110010;
assign micromatrizz[67][336] = 9'b111110011;
assign micromatrizz[67][337] = 9'b111110011;
assign micromatrizz[67][338] = 9'b111110011;
assign micromatrizz[67][339] = 9'b111110010;
assign micromatrizz[67][340] = 9'b111110010;
assign micromatrizz[67][341] = 9'b111110010;
assign micromatrizz[67][342] = 9'b111111111;
assign micromatrizz[67][343] = 9'b111111111;
assign micromatrizz[67][344] = 9'b111111111;
assign micromatrizz[67][345] = 9'b111111111;
assign micromatrizz[67][346] = 9'b111111111;
assign micromatrizz[67][347] = 9'b111110010;
assign micromatrizz[67][348] = 9'b111110010;
assign micromatrizz[67][349] = 9'b111110010;
assign micromatrizz[67][350] = 9'b111110010;
assign micromatrizz[67][351] = 9'b111110010;
assign micromatrizz[67][352] = 9'b111110011;
assign micromatrizz[67][353] = 9'b111110011;
assign micromatrizz[67][354] = 9'b111111111;
assign micromatrizz[67][355] = 9'b111111111;
assign micromatrizz[67][356] = 9'b111111111;
assign micromatrizz[67][357] = 9'b111111111;
assign micromatrizz[67][358] = 9'b111111111;
assign micromatrizz[67][359] = 9'b111110111;
assign micromatrizz[67][360] = 9'b111110010;
assign micromatrizz[67][361] = 9'b111110010;
assign micromatrizz[67][362] = 9'b111110010;
assign micromatrizz[67][363] = 9'b111110010;
assign micromatrizz[67][364] = 9'b111110011;
assign micromatrizz[67][365] = 9'b111110010;
assign micromatrizz[67][366] = 9'b111110111;
assign micromatrizz[67][367] = 9'b111111111;
assign micromatrizz[67][368] = 9'b111110011;
assign micromatrizz[67][369] = 9'b111111111;
assign micromatrizz[67][370] = 9'b111111111;
assign micromatrizz[67][371] = 9'b111111111;
assign micromatrizz[67][372] = 9'b111110010;
assign micromatrizz[67][373] = 9'b111110010;
assign micromatrizz[67][374] = 9'b111110011;
assign micromatrizz[67][375] = 9'b111110011;
assign micromatrizz[67][376] = 9'b111110011;
assign micromatrizz[67][377] = 9'b111110010;
assign micromatrizz[67][378] = 9'b111110010;
assign micromatrizz[67][379] = 9'b111111111;
assign micromatrizz[67][380] = 9'b111111111;
assign micromatrizz[67][381] = 9'b111111111;
assign micromatrizz[67][382] = 9'b111110111;
assign micromatrizz[67][383] = 9'b111110010;
assign micromatrizz[67][384] = 9'b111110010;
assign micromatrizz[67][385] = 9'b111110010;
assign micromatrizz[67][386] = 9'b111110011;
assign micromatrizz[67][387] = 9'b111110011;
assign micromatrizz[67][388] = 9'b111110011;
assign micromatrizz[67][389] = 9'b111110011;
assign micromatrizz[67][390] = 9'b111110011;
assign micromatrizz[67][391] = 9'b111111111;
assign micromatrizz[67][392] = 9'b111111111;
assign micromatrizz[67][393] = 9'b111111111;
assign micromatrizz[67][394] = 9'b111111111;
assign micromatrizz[67][395] = 9'b111110110;
assign micromatrizz[67][396] = 9'b111110010;
assign micromatrizz[67][397] = 9'b111110010;
assign micromatrizz[67][398] = 9'b111110010;
assign micromatrizz[67][399] = 9'b111110011;
assign micromatrizz[67][400] = 9'b111110011;
assign micromatrizz[67][401] = 9'b111110011;
assign micromatrizz[67][402] = 9'b111110111;
assign micromatrizz[67][403] = 9'b111111111;
assign micromatrizz[67][404] = 9'b111111111;
assign micromatrizz[67][405] = 9'b111111111;
assign micromatrizz[67][406] = 9'b111111111;
assign micromatrizz[67][407] = 9'b111111111;
assign micromatrizz[67][408] = 9'b111111111;
assign micromatrizz[67][409] = 9'b111111111;
assign micromatrizz[67][410] = 9'b111111111;
assign micromatrizz[67][411] = 9'b111111111;
assign micromatrizz[67][412] = 9'b111111111;
assign micromatrizz[67][413] = 9'b111110111;
assign micromatrizz[67][414] = 9'b111110010;
assign micromatrizz[67][415] = 9'b111110010;
assign micromatrizz[67][416] = 9'b111110010;
assign micromatrizz[67][417] = 9'b111110111;
assign micromatrizz[67][418] = 9'b111111111;
assign micromatrizz[67][419] = 9'b111111111;
assign micromatrizz[67][420] = 9'b111111111;
assign micromatrizz[67][421] = 9'b111111111;
assign micromatrizz[67][422] = 9'b111111111;
assign micromatrizz[67][423] = 9'b111111111;
assign micromatrizz[67][424] = 9'b111110110;
assign micromatrizz[67][425] = 9'b111110111;
assign micromatrizz[67][426] = 9'b111111111;
assign micromatrizz[67][427] = 9'b111111111;
assign micromatrizz[67][428] = 9'b111111111;
assign micromatrizz[67][429] = 9'b111111111;
assign micromatrizz[67][430] = 9'b111110111;
assign micromatrizz[67][431] = 9'b111110010;
assign micromatrizz[67][432] = 9'b111110010;
assign micromatrizz[67][433] = 9'b111110010;
assign micromatrizz[67][434] = 9'b111110010;
assign micromatrizz[67][435] = 9'b111110011;
assign micromatrizz[67][436] = 9'b111110011;
assign micromatrizz[67][437] = 9'b111110011;
assign micromatrizz[67][438] = 9'b111111111;
assign micromatrizz[67][439] = 9'b111111111;
assign micromatrizz[67][440] = 9'b111111111;
assign micromatrizz[67][441] = 9'b111111111;
assign micromatrizz[67][442] = 9'b111111111;
assign micromatrizz[67][443] = 9'b111111111;
assign micromatrizz[67][444] = 9'b111111111;
assign micromatrizz[67][445] = 9'b111111111;
assign micromatrizz[67][446] = 9'b111111111;
assign micromatrizz[67][447] = 9'b111111111;
assign micromatrizz[67][448] = 9'b111110111;
assign micromatrizz[67][449] = 9'b111110010;
assign micromatrizz[67][450] = 9'b111110011;
assign micromatrizz[67][451] = 9'b111110010;
assign micromatrizz[67][452] = 9'b111110011;
assign micromatrizz[67][453] = 9'b111110011;
assign micromatrizz[67][454] = 9'b111111111;
assign micromatrizz[67][455] = 9'b111111111;
assign micromatrizz[67][456] = 9'b111111111;
assign micromatrizz[67][457] = 9'b111111111;
assign micromatrizz[67][458] = 9'b111111111;
assign micromatrizz[67][459] = 9'b111110111;
assign micromatrizz[67][460] = 9'b111110111;
assign micromatrizz[67][461] = 9'b111111111;
assign micromatrizz[67][462] = 9'b111111111;
assign micromatrizz[67][463] = 9'b111111111;
assign micromatrizz[67][464] = 9'b111111111;
assign micromatrizz[67][465] = 9'b111110010;
assign micromatrizz[67][466] = 9'b111110111;
assign micromatrizz[67][467] = 9'b111111111;
assign micromatrizz[67][468] = 9'b111111111;
assign micromatrizz[67][469] = 9'b111111111;
assign micromatrizz[67][470] = 9'b111111111;
assign micromatrizz[67][471] = 9'b111110111;
assign micromatrizz[67][472] = 9'b111110010;
assign micromatrizz[67][473] = 9'b111110011;
assign micromatrizz[67][474] = 9'b111110011;
assign micromatrizz[67][475] = 9'b111110011;
assign micromatrizz[67][476] = 9'b111110010;
assign micromatrizz[67][477] = 9'b111111111;
assign micromatrizz[67][478] = 9'b111111111;
assign micromatrizz[67][479] = 9'b111111111;
assign micromatrizz[67][480] = 9'b111111111;
assign micromatrizz[67][481] = 9'b111110010;
assign micromatrizz[67][482] = 9'b111110010;
assign micromatrizz[67][483] = 9'b111110011;
assign micromatrizz[67][484] = 9'b111110011;
assign micromatrizz[67][485] = 9'b111110011;
assign micromatrizz[67][486] = 9'b111110011;
assign micromatrizz[67][487] = 9'b111110011;
assign micromatrizz[67][488] = 9'b111110111;
assign micromatrizz[67][489] = 9'b111111111;
assign micromatrizz[67][490] = 9'b111111111;
assign micromatrizz[67][491] = 9'b111111111;
assign micromatrizz[67][492] = 9'b111111111;
assign micromatrizz[67][493] = 9'b111111111;
assign micromatrizz[67][494] = 9'b111111111;
assign micromatrizz[67][495] = 9'b111111111;
assign micromatrizz[67][496] = 9'b111111111;
assign micromatrizz[67][497] = 9'b111111111;
assign micromatrizz[67][498] = 9'b111111111;
assign micromatrizz[67][499] = 9'b111110111;
assign micromatrizz[67][500] = 9'b111110010;
assign micromatrizz[67][501] = 9'b111110010;
assign micromatrizz[67][502] = 9'b111110010;
assign micromatrizz[67][503] = 9'b111110111;
assign micromatrizz[67][504] = 9'b111111111;
assign micromatrizz[67][505] = 9'b111111111;
assign micromatrizz[67][506] = 9'b111111111;
assign micromatrizz[67][507] = 9'b111111111;
assign micromatrizz[67][508] = 9'b111111111;
assign micromatrizz[67][509] = 9'b111111111;
assign micromatrizz[67][510] = 9'b111110010;
assign micromatrizz[67][511] = 9'b111110111;
assign micromatrizz[67][512] = 9'b111111111;
assign micromatrizz[67][513] = 9'b111111111;
assign micromatrizz[67][514] = 9'b111111111;
assign micromatrizz[67][515] = 9'b111111111;
assign micromatrizz[67][516] = 9'b111110110;
assign micromatrizz[67][517] = 9'b111110010;
assign micromatrizz[67][518] = 9'b111110011;
assign micromatrizz[67][519] = 9'b111110010;
assign micromatrizz[67][520] = 9'b111110010;
assign micromatrizz[67][521] = 9'b111110010;
assign micromatrizz[67][522] = 9'b111110011;
assign micromatrizz[67][523] = 9'b111110011;
assign micromatrizz[67][524] = 9'b111110111;
assign micromatrizz[67][525] = 9'b111111111;
assign micromatrizz[67][526] = 9'b111111111;
assign micromatrizz[67][527] = 9'b111111111;
assign micromatrizz[67][528] = 9'b111110111;
assign micromatrizz[67][529] = 9'b111110010;
assign micromatrizz[67][530] = 9'b111110010;
assign micromatrizz[67][531] = 9'b111110010;
assign micromatrizz[67][532] = 9'b111110011;
assign micromatrizz[67][533] = 9'b111110010;
assign micromatrizz[67][534] = 9'b111111111;
assign micromatrizz[67][535] = 9'b111111111;
assign micromatrizz[67][536] = 9'b111111111;
assign micromatrizz[67][537] = 9'b111111111;
assign micromatrizz[67][538] = 9'b111111111;
assign micromatrizz[67][539] = 9'b111111111;
assign micromatrizz[67][540] = 9'b111111111;
assign micromatrizz[67][541] = 9'b111110010;
assign micromatrizz[67][542] = 9'b111110010;
assign micromatrizz[67][543] = 9'b111110011;
assign micromatrizz[67][544] = 9'b111110010;
assign micromatrizz[67][545] = 9'b111111111;
assign micromatrizz[67][546] = 9'b111111111;
assign micromatrizz[67][547] = 9'b111111111;
assign micromatrizz[67][548] = 9'b111111111;
assign micromatrizz[67][549] = 9'b111111111;
assign micromatrizz[67][550] = 9'b111111111;
assign micromatrizz[67][551] = 9'b111110111;
assign micromatrizz[67][552] = 9'b111110010;
assign micromatrizz[67][553] = 9'b111111111;
assign micromatrizz[67][554] = 9'b111111111;
assign micromatrizz[67][555] = 9'b111111111;
assign micromatrizz[67][556] = 9'b111111111;
assign micromatrizz[67][557] = 9'b111111111;
assign micromatrizz[67][558] = 9'b111110010;
assign micromatrizz[67][559] = 9'b111110010;
assign micromatrizz[67][560] = 9'b111110010;
assign micromatrizz[67][561] = 9'b111110010;
assign micromatrizz[67][562] = 9'b111110011;
assign micromatrizz[67][563] = 9'b111110011;
assign micromatrizz[67][564] = 9'b111110010;
assign micromatrizz[67][565] = 9'b111111111;
assign micromatrizz[67][566] = 9'b111111111;
assign micromatrizz[67][567] = 9'b111111111;
assign micromatrizz[67][568] = 9'b111111111;
assign micromatrizz[67][569] = 9'b111111111;
assign micromatrizz[67][570] = 9'b111110111;
assign micromatrizz[67][571] = 9'b111110010;
assign micromatrizz[67][572] = 9'b111110010;
assign micromatrizz[67][573] = 9'b111110011;
assign micromatrizz[67][574] = 9'b111110011;
assign micromatrizz[67][575] = 9'b111110010;
assign micromatrizz[67][576] = 9'b111111111;
assign micromatrizz[67][577] = 9'b111111111;
assign micromatrizz[67][578] = 9'b111111111;
assign micromatrizz[67][579] = 9'b111110110;
assign micromatrizz[67][580] = 9'b111110010;
assign micromatrizz[67][581] = 9'b111110011;
assign micromatrizz[67][582] = 9'b111110010;
assign micromatrizz[67][583] = 9'b111110011;
assign micromatrizz[67][584] = 9'b111110011;
assign micromatrizz[67][585] = 9'b111110011;
assign micromatrizz[67][586] = 9'b111110011;
assign micromatrizz[67][587] = 9'b111110011;
assign micromatrizz[67][588] = 9'b111111111;
assign micromatrizz[67][589] = 9'b111111111;
assign micromatrizz[67][590] = 9'b111111111;
assign micromatrizz[67][591] = 9'b111111111;
assign micromatrizz[67][592] = 9'b111111111;
assign micromatrizz[67][593] = 9'b111111111;
assign micromatrizz[67][594] = 9'b111110010;
assign micromatrizz[67][595] = 9'b111110010;
assign micromatrizz[67][596] = 9'b111110010;
assign micromatrizz[67][597] = 9'b111110010;
assign micromatrizz[67][598] = 9'b111111111;
assign micromatrizz[67][599] = 9'b111111111;
assign micromatrizz[67][600] = 9'b111111111;
assign micromatrizz[67][601] = 9'b111111111;
assign micromatrizz[67][602] = 9'b111111111;
assign micromatrizz[67][603] = 9'b111111111;
assign micromatrizz[67][604] = 9'b111110111;
assign micromatrizz[67][605] = 9'b111110010;
assign micromatrizz[67][606] = 9'b111111111;
assign micromatrizz[67][607] = 9'b111111111;
assign micromatrizz[67][608] = 9'b111111111;
assign micromatrizz[67][609] = 9'b111111111;
assign micromatrizz[67][610] = 9'b111110010;
assign micromatrizz[67][611] = 9'b111110111;
assign micromatrizz[67][612] = 9'b111111111;
assign micromatrizz[67][613] = 9'b111111111;
assign micromatrizz[67][614] = 9'b111111111;
assign micromatrizz[67][615] = 9'b111111111;
assign micromatrizz[67][616] = 9'b111111111;
assign micromatrizz[67][617] = 9'b111110010;
assign micromatrizz[67][618] = 9'b111110010;
assign micromatrizz[67][619] = 9'b111110011;
assign micromatrizz[67][620] = 9'b111110011;
assign micromatrizz[67][621] = 9'b111110010;
assign micromatrizz[67][622] = 9'b111111111;
assign micromatrizz[67][623] = 9'b111111111;
assign micromatrizz[67][624] = 9'b111111111;
assign micromatrizz[67][625] = 9'b111111111;
assign micromatrizz[67][626] = 9'b111111111;
assign micromatrizz[67][627] = 9'b111111111;
assign micromatrizz[67][628] = 9'b111111111;
assign micromatrizz[67][629] = 9'b111111111;
assign micromatrizz[67][630] = 9'b111111111;
assign micromatrizz[67][631] = 9'b111111111;
assign micromatrizz[67][632] = 9'b111111111;
assign micromatrizz[67][633] = 9'b111111111;
assign micromatrizz[67][634] = 9'b111111111;
assign micromatrizz[67][635] = 9'b111111111;
assign micromatrizz[67][636] = 9'b111111111;
assign micromatrizz[67][637] = 9'b111111111;
assign micromatrizz[67][638] = 9'b111111111;
assign micromatrizz[67][639] = 9'b111111111;
assign micromatrizz[68][0] = 9'b111111111;
assign micromatrizz[68][1] = 9'b111111111;
assign micromatrizz[68][2] = 9'b111111111;
assign micromatrizz[68][3] = 9'b111111111;
assign micromatrizz[68][4] = 9'b111111111;
assign micromatrizz[68][5] = 9'b111111111;
assign micromatrizz[68][6] = 9'b111111111;
assign micromatrizz[68][7] = 9'b111111111;
assign micromatrizz[68][8] = 9'b111111111;
assign micromatrizz[68][9] = 9'b111110010;
assign micromatrizz[68][10] = 9'b111110111;
assign micromatrizz[68][11] = 9'b111111111;
assign micromatrizz[68][12] = 9'b111111111;
assign micromatrizz[68][13] = 9'b111111111;
assign micromatrizz[68][14] = 9'b111111111;
assign micromatrizz[68][15] = 9'b111110010;
assign micromatrizz[68][16] = 9'b111110010;
assign micromatrizz[68][17] = 9'b111110010;
assign micromatrizz[68][18] = 9'b111110011;
assign micromatrizz[68][19] = 9'b111111111;
assign micromatrizz[68][20] = 9'b111111111;
assign micromatrizz[68][21] = 9'b111111111;
assign micromatrizz[68][22] = 9'b111111111;
assign micromatrizz[68][23] = 9'b111111111;
assign micromatrizz[68][24] = 9'b111110111;
assign micromatrizz[68][25] = 9'b111110010;
assign micromatrizz[68][26] = 9'b111110010;
assign micromatrizz[68][27] = 9'b111110010;
assign micromatrizz[68][28] = 9'b111110011;
assign micromatrizz[68][29] = 9'b111110011;
assign micromatrizz[68][30] = 9'b111110011;
assign micromatrizz[68][31] = 9'b111110111;
assign micromatrizz[68][32] = 9'b111111111;
assign micromatrizz[68][33] = 9'b111110111;
assign micromatrizz[68][34] = 9'b111110111;
assign micromatrizz[68][35] = 9'b111110111;
assign micromatrizz[68][36] = 9'b111110010;
assign micromatrizz[68][37] = 9'b111110010;
assign micromatrizz[68][38] = 9'b111110011;
assign micromatrizz[68][39] = 9'b111110010;
assign micromatrizz[68][40] = 9'b111110011;
assign micromatrizz[68][41] = 9'b111110011;
assign micromatrizz[68][42] = 9'b111110010;
assign micromatrizz[68][43] = 9'b111111111;
assign micromatrizz[68][44] = 9'b111111111;
assign micromatrizz[68][45] = 9'b111111111;
assign micromatrizz[68][46] = 9'b111111111;
assign micromatrizz[68][47] = 9'b111110010;
assign micromatrizz[68][48] = 9'b111110010;
assign micromatrizz[68][49] = 9'b111110011;
assign micromatrizz[68][50] = 9'b111110011;
assign micromatrizz[68][51] = 9'b111110011;
assign micromatrizz[68][52] = 9'b111110011;
assign micromatrizz[68][53] = 9'b111110010;
assign micromatrizz[68][54] = 9'b111110111;
assign micromatrizz[68][55] = 9'b111111111;
assign micromatrizz[68][56] = 9'b111111111;
assign micromatrizz[68][57] = 9'b111111111;
assign micromatrizz[68][58] = 9'b111111111;
assign micromatrizz[68][59] = 9'b111111111;
assign micromatrizz[68][60] = 9'b111111111;
assign micromatrizz[68][61] = 9'b111111111;
assign micromatrizz[68][62] = 9'b111111111;
assign micromatrizz[68][63] = 9'b111111111;
assign micromatrizz[68][64] = 9'b111111111;
assign micromatrizz[68][65] = 9'b111111111;
assign micromatrizz[68][66] = 9'b111111111;
assign micromatrizz[68][67] = 9'b111111111;
assign micromatrizz[68][68] = 9'b111111111;
assign micromatrizz[68][69] = 9'b111111111;
assign micromatrizz[68][70] = 9'b111111111;
assign micromatrizz[68][71] = 9'b111111111;
assign micromatrizz[68][72] = 9'b111110111;
assign micromatrizz[68][73] = 9'b111110010;
assign micromatrizz[68][74] = 9'b111110010;
assign micromatrizz[68][75] = 9'b111110111;
assign micromatrizz[68][76] = 9'b111111111;
assign micromatrizz[68][77] = 9'b111111111;
assign micromatrizz[68][78] = 9'b111111111;
assign micromatrizz[68][79] = 9'b111111111;
assign micromatrizz[68][80] = 9'b111110111;
assign micromatrizz[68][81] = 9'b111110111;
assign micromatrizz[68][82] = 9'b111111111;
assign micromatrizz[68][83] = 9'b111111111;
assign micromatrizz[68][84] = 9'b111111111;
assign micromatrizz[68][85] = 9'b111111111;
assign micromatrizz[68][86] = 9'b111111111;
assign micromatrizz[68][87] = 9'b111111111;
assign micromatrizz[68][88] = 9'b111110010;
assign micromatrizz[68][89] = 9'b111110010;
assign micromatrizz[68][90] = 9'b111110011;
assign micromatrizz[68][91] = 9'b111110011;
assign micromatrizz[68][92] = 9'b111110011;
assign micromatrizz[68][93] = 9'b111110010;
assign micromatrizz[68][94] = 9'b111110010;
assign micromatrizz[68][95] = 9'b111110111;
assign micromatrizz[68][96] = 9'b111111111;
assign micromatrizz[68][97] = 9'b111111111;
assign micromatrizz[68][98] = 9'b111111111;
assign micromatrizz[68][99] = 9'b111111111;
assign micromatrizz[68][100] = 9'b111111111;
assign micromatrizz[68][101] = 9'b111111111;
assign micromatrizz[68][102] = 9'b111111111;
assign micromatrizz[68][103] = 9'b111111111;
assign micromatrizz[68][104] = 9'b111111111;
assign micromatrizz[68][105] = 9'b111110110;
assign micromatrizz[68][106] = 9'b111110111;
assign micromatrizz[68][107] = 9'b111111111;
assign micromatrizz[68][108] = 9'b111111111;
assign micromatrizz[68][109] = 9'b111111111;
assign micromatrizz[68][110] = 9'b111111111;
assign micromatrizz[68][111] = 9'b111110010;
assign micromatrizz[68][112] = 9'b111110010;
assign micromatrizz[68][113] = 9'b111110010;
assign micromatrizz[68][114] = 9'b111110010;
assign micromatrizz[68][115] = 9'b111111111;
assign micromatrizz[68][116] = 9'b111111111;
assign micromatrizz[68][117] = 9'b111111111;
assign micromatrizz[68][118] = 9'b111111111;
assign micromatrizz[68][119] = 9'b111111111;
assign micromatrizz[68][120] = 9'b111111111;
assign micromatrizz[68][121] = 9'b111111111;
assign micromatrizz[68][122] = 9'b111110111;
assign micromatrizz[68][123] = 9'b111110010;
assign micromatrizz[68][124] = 9'b111110010;
assign micromatrizz[68][125] = 9'b111110011;
assign micromatrizz[68][126] = 9'b111110011;
assign micromatrizz[68][127] = 9'b111111111;
assign micromatrizz[68][128] = 9'b111111111;
assign micromatrizz[68][129] = 9'b111111111;
assign micromatrizz[68][130] = 9'b111111111;
assign micromatrizz[68][131] = 9'b111110110;
assign micromatrizz[68][132] = 9'b111111111;
assign micromatrizz[68][133] = 9'b111111111;
assign micromatrizz[68][134] = 9'b111111111;
assign micromatrizz[68][135] = 9'b111111111;
assign micromatrizz[68][136] = 9'b111111111;
assign micromatrizz[68][137] = 9'b111111111;
assign micromatrizz[68][138] = 9'b111110111;
assign micromatrizz[68][139] = 9'b111110010;
assign micromatrizz[68][140] = 9'b111110010;
assign micromatrizz[68][141] = 9'b111110010;
assign micromatrizz[68][142] = 9'b111110010;
assign micromatrizz[68][143] = 9'b111110010;
assign micromatrizz[68][144] = 9'b111110011;
assign micromatrizz[68][145] = 9'b111110011;
assign micromatrizz[68][146] = 9'b111111111;
assign micromatrizz[68][147] = 9'b111111111;
assign micromatrizz[68][148] = 9'b111111111;
assign micromatrizz[68][149] = 9'b111111111;
assign micromatrizz[68][150] = 9'b111110111;
assign micromatrizz[68][151] = 9'b111110010;
assign micromatrizz[68][152] = 9'b111110011;
assign micromatrizz[68][153] = 9'b111110011;
assign micromatrizz[68][154] = 9'b111110010;
assign micromatrizz[68][155] = 9'b111110011;
assign micromatrizz[68][156] = 9'b111110011;
assign micromatrizz[68][157] = 9'b111110011;
assign micromatrizz[68][158] = 9'b111111111;
assign micromatrizz[68][159] = 9'b111111111;
assign micromatrizz[68][160] = 9'b111111111;
assign micromatrizz[68][161] = 9'b111111111;
assign micromatrizz[68][162] = 9'b111110111;
assign micromatrizz[68][163] = 9'b111110010;
assign micromatrizz[68][164] = 9'b111110010;
assign micromatrizz[68][165] = 9'b111110011;
assign micromatrizz[68][166] = 9'b111110011;
assign micromatrizz[68][167] = 9'b111110011;
assign micromatrizz[68][168] = 9'b111110111;
assign micromatrizz[68][169] = 9'b111111111;
assign micromatrizz[68][170] = 9'b111110111;
assign micromatrizz[68][171] = 9'b111110111;
assign micromatrizz[68][172] = 9'b111110010;
assign micromatrizz[68][173] = 9'b111110010;
assign micromatrizz[68][174] = 9'b111110011;
assign micromatrizz[68][175] = 9'b111110011;
assign micromatrizz[68][176] = 9'b111110011;
assign micromatrizz[68][177] = 9'b111110011;
assign micromatrizz[68][178] = 9'b111110010;
assign micromatrizz[68][179] = 9'b111110111;
assign micromatrizz[68][180] = 9'b111111111;
assign micromatrizz[68][181] = 9'b111111111;
assign micromatrizz[68][182] = 9'b111111111;
assign micromatrizz[68][183] = 9'b111111111;
assign micromatrizz[68][184] = 9'b111111111;
assign micromatrizz[68][185] = 9'b111111111;
assign micromatrizz[68][186] = 9'b111110010;
assign micromatrizz[68][187] = 9'b111110010;
assign micromatrizz[68][188] = 9'b111110011;
assign micromatrizz[68][189] = 9'b111110011;
assign micromatrizz[68][190] = 9'b111110011;
assign micromatrizz[68][191] = 9'b111111111;
assign micromatrizz[68][192] = 9'b111110111;
assign micromatrizz[68][193] = 9'b111110111;
assign micromatrizz[68][194] = 9'b111110111;
assign micromatrizz[68][195] = 9'b111110010;
assign micromatrizz[68][196] = 9'b111110011;
assign micromatrizz[68][197] = 9'b111110011;
assign micromatrizz[68][198] = 9'b111110011;
assign micromatrizz[68][199] = 9'b111110010;
assign micromatrizz[68][200] = 9'b111110010;
assign micromatrizz[68][201] = 9'b111110010;
assign micromatrizz[68][202] = 9'b111110111;
assign micromatrizz[68][203] = 9'b111111111;
assign micromatrizz[68][204] = 9'b111111111;
assign micromatrizz[68][205] = 9'b111111111;
assign micromatrizz[68][206] = 9'b111111111;
assign micromatrizz[68][207] = 9'b111111111;
assign micromatrizz[68][208] = 9'b111111111;
assign micromatrizz[68][209] = 9'b111110111;
assign micromatrizz[68][210] = 9'b111110010;
assign micromatrizz[68][211] = 9'b111110010;
assign micromatrizz[68][212] = 9'b111110010;
assign micromatrizz[68][213] = 9'b111110111;
assign micromatrizz[68][214] = 9'b111111111;
assign micromatrizz[68][215] = 9'b111111111;
assign micromatrizz[68][216] = 9'b111111111;
assign micromatrizz[68][217] = 9'b111110111;
assign micromatrizz[68][218] = 9'b111110111;
assign micromatrizz[68][219] = 9'b111111111;
assign micromatrizz[68][220] = 9'b111111111;
assign micromatrizz[68][221] = 9'b111111111;
assign micromatrizz[68][222] = 9'b111111111;
assign micromatrizz[68][223] = 9'b111111111;
assign micromatrizz[68][224] = 9'b111111111;
assign micromatrizz[68][225] = 9'b111110011;
assign micromatrizz[68][226] = 9'b111110010;
assign micromatrizz[68][227] = 9'b111110010;
assign micromatrizz[68][228] = 9'b111110010;
assign micromatrizz[68][229] = 9'b111110011;
assign micromatrizz[68][230] = 9'b111110011;
assign micromatrizz[68][231] = 9'b111110011;
assign micromatrizz[68][232] = 9'b111110111;
assign micromatrizz[68][233] = 9'b111111111;
assign micromatrizz[68][234] = 9'b111111111;
assign micromatrizz[68][235] = 9'b111111111;
assign micromatrizz[68][236] = 9'b111111111;
assign micromatrizz[68][237] = 9'b111111111;
assign micromatrizz[68][238] = 9'b111111111;
assign micromatrizz[68][239] = 9'b111111111;
assign micromatrizz[68][240] = 9'b111111111;
assign micromatrizz[68][241] = 9'b111111111;
assign micromatrizz[68][242] = 9'b111111111;
assign micromatrizz[68][243] = 9'b111111111;
assign micromatrizz[68][244] = 9'b111110111;
assign micromatrizz[68][245] = 9'b111110010;
assign micromatrizz[68][246] = 9'b111110010;
assign micromatrizz[68][247] = 9'b111110011;
assign micromatrizz[68][248] = 9'b111111111;
assign micromatrizz[68][249] = 9'b111111111;
assign micromatrizz[68][250] = 9'b111111111;
assign micromatrizz[68][251] = 9'b111111111;
assign micromatrizz[68][252] = 9'b111111111;
assign micromatrizz[68][253] = 9'b111110110;
assign micromatrizz[68][254] = 9'b111111111;
assign micromatrizz[68][255] = 9'b111111111;
assign micromatrizz[68][256] = 9'b111111111;
assign micromatrizz[68][257] = 9'b111111111;
assign micromatrizz[68][258] = 9'b111111111;
assign micromatrizz[68][259] = 9'b111111111;
assign micromatrizz[68][260] = 9'b111110111;
assign micromatrizz[68][261] = 9'b111110110;
assign micromatrizz[68][262] = 9'b111111111;
assign micromatrizz[68][263] = 9'b111111111;
assign micromatrizz[68][264] = 9'b111111111;
assign micromatrizz[68][265] = 9'b111111111;
assign micromatrizz[68][266] = 9'b111110111;
assign micromatrizz[68][267] = 9'b111110010;
assign micromatrizz[68][268] = 9'b111110010;
assign micromatrizz[68][269] = 9'b111110010;
assign micromatrizz[68][270] = 9'b111110111;
assign micromatrizz[68][271] = 9'b111111111;
assign micromatrizz[68][272] = 9'b111111111;
assign micromatrizz[68][273] = 9'b111111111;
assign micromatrizz[68][274] = 9'b111111111;
assign micromatrizz[68][275] = 9'b111111111;
assign micromatrizz[68][276] = 9'b111110111;
assign micromatrizz[68][277] = 9'b111110010;
assign micromatrizz[68][278] = 9'b111110010;
assign micromatrizz[68][279] = 9'b111110011;
assign micromatrizz[68][280] = 9'b111110011;
assign micromatrizz[68][281] = 9'b111110011;
assign micromatrizz[68][282] = 9'b111110111;
assign micromatrizz[68][283] = 9'b111111111;
assign micromatrizz[68][284] = 9'b111110111;
assign micromatrizz[68][285] = 9'b111110111;
assign micromatrizz[68][286] = 9'b111110011;
assign micromatrizz[68][287] = 9'b111110010;
assign micromatrizz[68][288] = 9'b111110010;
assign micromatrizz[68][289] = 9'b111110011;
assign micromatrizz[68][290] = 9'b111110011;
assign micromatrizz[68][291] = 9'b111110011;
assign micromatrizz[68][292] = 9'b111110011;
assign micromatrizz[68][293] = 9'b111110111;
assign micromatrizz[68][294] = 9'b111111111;
assign micromatrizz[68][295] = 9'b111111111;
assign micromatrizz[68][296] = 9'b111111111;
assign micromatrizz[68][297] = 9'b111111111;
assign micromatrizz[68][298] = 9'b111111111;
assign micromatrizz[68][299] = 9'b111111111;
assign micromatrizz[68][300] = 9'b111111111;
assign micromatrizz[68][301] = 9'b111111111;
assign micromatrizz[68][302] = 9'b111111111;
assign micromatrizz[68][303] = 9'b111111111;
assign micromatrizz[68][304] = 9'b111110111;
assign micromatrizz[68][305] = 9'b111110010;
assign micromatrizz[68][306] = 9'b111110111;
assign micromatrizz[68][307] = 9'b111111111;
assign micromatrizz[68][308] = 9'b111111111;
assign micromatrizz[68][309] = 9'b111111111;
assign micromatrizz[68][310] = 9'b111111111;
assign micromatrizz[68][311] = 9'b111111111;
assign micromatrizz[68][312] = 9'b111111111;
assign micromatrizz[68][313] = 9'b111111111;
assign micromatrizz[68][314] = 9'b111111111;
assign micromatrizz[68][315] = 9'b111111111;
assign micromatrizz[68][316] = 9'b111111111;
assign micromatrizz[68][317] = 9'b111111111;
assign micromatrizz[68][318] = 9'b111111111;
assign micromatrizz[68][319] = 9'b111110111;
assign micromatrizz[68][320] = 9'b111110010;
assign micromatrizz[68][321] = 9'b111110010;
assign micromatrizz[68][322] = 9'b111110111;
assign micromatrizz[68][323] = 9'b111111111;
assign micromatrizz[68][324] = 9'b111111111;
assign micromatrizz[68][325] = 9'b111111111;
assign micromatrizz[68][326] = 9'b111111111;
assign micromatrizz[68][327] = 9'b111110111;
assign micromatrizz[68][328] = 9'b111110111;
assign micromatrizz[68][329] = 9'b111111111;
assign micromatrizz[68][330] = 9'b111111111;
assign micromatrizz[68][331] = 9'b111111111;
assign micromatrizz[68][332] = 9'b111111111;
assign micromatrizz[68][333] = 9'b111111111;
assign micromatrizz[68][334] = 9'b111111111;
assign micromatrizz[68][335] = 9'b111110010;
assign micromatrizz[68][336] = 9'b111110011;
assign micromatrizz[68][337] = 9'b111110011;
assign micromatrizz[68][338] = 9'b111110010;
assign micromatrizz[68][339] = 9'b111110010;
assign micromatrizz[68][340] = 9'b111110011;
assign micromatrizz[68][341] = 9'b111110010;
assign micromatrizz[68][342] = 9'b111110111;
assign micromatrizz[68][343] = 9'b111111111;
assign micromatrizz[68][344] = 9'b111111111;
assign micromatrizz[68][345] = 9'b111111111;
assign micromatrizz[68][346] = 9'b111111111;
assign micromatrizz[68][347] = 9'b111110010;
assign micromatrizz[68][348] = 9'b111110010;
assign micromatrizz[68][349] = 9'b111110010;
assign micromatrizz[68][350] = 9'b111110010;
assign micromatrizz[68][351] = 9'b111110010;
assign micromatrizz[68][352] = 9'b111110011;
assign micromatrizz[68][353] = 9'b111110011;
assign micromatrizz[68][354] = 9'b111111111;
assign micromatrizz[68][355] = 9'b111111111;
assign micromatrizz[68][356] = 9'b111111111;
assign micromatrizz[68][357] = 9'b111111111;
assign micromatrizz[68][358] = 9'b111111111;
assign micromatrizz[68][359] = 9'b111111111;
assign micromatrizz[68][360] = 9'b111110011;
assign micromatrizz[68][361] = 9'b111110010;
assign micromatrizz[68][362] = 9'b111110010;
assign micromatrizz[68][363] = 9'b111110010;
assign micromatrizz[68][364] = 9'b111110010;
assign micromatrizz[68][365] = 9'b111110011;
assign micromatrizz[68][366] = 9'b111110011;
assign micromatrizz[68][367] = 9'b111110010;
assign micromatrizz[68][368] = 9'b111110111;
assign micromatrizz[68][369] = 9'b111111111;
assign micromatrizz[68][370] = 9'b111111111;
assign micromatrizz[68][371] = 9'b111111111;
assign micromatrizz[68][372] = 9'b111111111;
assign micromatrizz[68][373] = 9'b111110010;
assign micromatrizz[68][374] = 9'b111110011;
assign micromatrizz[68][375] = 9'b111110011;
assign micromatrizz[68][376] = 9'b111110010;
assign micromatrizz[68][377] = 9'b111110010;
assign micromatrizz[68][378] = 9'b111110011;
assign micromatrizz[68][379] = 9'b111110111;
assign micromatrizz[68][380] = 9'b111111111;
assign micromatrizz[68][381] = 9'b111110111;
assign micromatrizz[68][382] = 9'b111110110;
assign micromatrizz[68][383] = 9'b111110111;
assign micromatrizz[68][384] = 9'b111110010;
assign micromatrizz[68][385] = 9'b111110010;
assign micromatrizz[68][386] = 9'b111110011;
assign micromatrizz[68][387] = 9'b111110011;
assign micromatrizz[68][388] = 9'b111110010;
assign micromatrizz[68][389] = 9'b111110011;
assign micromatrizz[68][390] = 9'b111110011;
assign micromatrizz[68][391] = 9'b111111111;
assign micromatrizz[68][392] = 9'b111111111;
assign micromatrizz[68][393] = 9'b111111111;
assign micromatrizz[68][394] = 9'b111111111;
assign micromatrizz[68][395] = 9'b111110111;
assign micromatrizz[68][396] = 9'b111110010;
assign micromatrizz[68][397] = 9'b111110010;
assign micromatrizz[68][398] = 9'b111110011;
assign micromatrizz[68][399] = 9'b111110011;
assign micromatrizz[68][400] = 9'b111110011;
assign micromatrizz[68][401] = 9'b111110011;
assign micromatrizz[68][402] = 9'b111110111;
assign micromatrizz[68][403] = 9'b111111111;
assign micromatrizz[68][404] = 9'b111111111;
assign micromatrizz[68][405] = 9'b111111111;
assign micromatrizz[68][406] = 9'b111111111;
assign micromatrizz[68][407] = 9'b111111111;
assign micromatrizz[68][408] = 9'b111111111;
assign micromatrizz[68][409] = 9'b111111111;
assign micromatrizz[68][410] = 9'b111111111;
assign micromatrizz[68][411] = 9'b111111111;
assign micromatrizz[68][412] = 9'b111111111;
assign micromatrizz[68][413] = 9'b111111111;
assign micromatrizz[68][414] = 9'b111110111;
assign micromatrizz[68][415] = 9'b111110010;
assign micromatrizz[68][416] = 9'b111110010;
assign micromatrizz[68][417] = 9'b111110011;
assign micromatrizz[68][418] = 9'b111111111;
assign micromatrizz[68][419] = 9'b111111111;
assign micromatrizz[68][420] = 9'b111111111;
assign micromatrizz[68][421] = 9'b111111111;
assign micromatrizz[68][422] = 9'b111111111;
assign micromatrizz[68][423] = 9'b111110110;
assign micromatrizz[68][424] = 9'b111111111;
assign micromatrizz[68][425] = 9'b111111111;
assign micromatrizz[68][426] = 9'b111111111;
assign micromatrizz[68][427] = 9'b111111111;
assign micromatrizz[68][428] = 9'b111111111;
assign micromatrizz[68][429] = 9'b111111111;
assign micromatrizz[68][430] = 9'b111110111;
assign micromatrizz[68][431] = 9'b111110010;
assign micromatrizz[68][432] = 9'b111110010;
assign micromatrizz[68][433] = 9'b111110010;
assign micromatrizz[68][434] = 9'b111110010;
assign micromatrizz[68][435] = 9'b111110011;
assign micromatrizz[68][436] = 9'b111110011;
assign micromatrizz[68][437] = 9'b111110011;
assign micromatrizz[68][438] = 9'b111111111;
assign micromatrizz[68][439] = 9'b111111111;
assign micromatrizz[68][440] = 9'b111111111;
assign micromatrizz[68][441] = 9'b111111111;
assign micromatrizz[68][442] = 9'b111111111;
assign micromatrizz[68][443] = 9'b111111111;
assign micromatrizz[68][444] = 9'b111111111;
assign micromatrizz[68][445] = 9'b111111111;
assign micromatrizz[68][446] = 9'b111111111;
assign micromatrizz[68][447] = 9'b111111111;
assign micromatrizz[68][448] = 9'b111111111;
assign micromatrizz[68][449] = 9'b111111111;
assign micromatrizz[68][450] = 9'b111110110;
assign micromatrizz[68][451] = 9'b111110010;
assign micromatrizz[68][452] = 9'b111110011;
assign micromatrizz[68][453] = 9'b111110011;
assign micromatrizz[68][454] = 9'b111111111;
assign micromatrizz[68][455] = 9'b111111111;
assign micromatrizz[68][456] = 9'b111111111;
assign micromatrizz[68][457] = 9'b111111111;
assign micromatrizz[68][458] = 9'b111110111;
assign micromatrizz[68][459] = 9'b111110111;
assign micromatrizz[68][460] = 9'b111111111;
assign micromatrizz[68][461] = 9'b111111111;
assign micromatrizz[68][462] = 9'b111111111;
assign micromatrizz[68][463] = 9'b111111111;
assign micromatrizz[68][464] = 9'b111111111;
assign micromatrizz[68][465] = 9'b111111111;
assign micromatrizz[68][466] = 9'b111110010;
assign micromatrizz[68][467] = 9'b111110111;
assign micromatrizz[68][468] = 9'b111111111;
assign micromatrizz[68][469] = 9'b111111111;
assign micromatrizz[68][470] = 9'b111111111;
assign micromatrizz[68][471] = 9'b111111111;
assign micromatrizz[68][472] = 9'b111110010;
assign micromatrizz[68][473] = 9'b111110010;
assign micromatrizz[68][474] = 9'b111110010;
assign micromatrizz[68][475] = 9'b111110010;
assign micromatrizz[68][476] = 9'b111111111;
assign micromatrizz[68][477] = 9'b111111111;
assign micromatrizz[68][478] = 9'b111111111;
assign micromatrizz[68][479] = 9'b111111111;
assign micromatrizz[68][480] = 9'b111111111;
assign micromatrizz[68][481] = 9'b111110011;
assign micromatrizz[68][482] = 9'b111110010;
assign micromatrizz[68][483] = 9'b111110011;
assign micromatrizz[68][484] = 9'b111110011;
assign micromatrizz[68][485] = 9'b111110011;
assign micromatrizz[68][486] = 9'b111110011;
assign micromatrizz[68][487] = 9'b111110010;
assign micromatrizz[68][488] = 9'b111110111;
assign micromatrizz[68][489] = 9'b111111111;
assign micromatrizz[68][490] = 9'b111111111;
assign micromatrizz[68][491] = 9'b111111111;
assign micromatrizz[68][492] = 9'b111111111;
assign micromatrizz[68][493] = 9'b111111111;
assign micromatrizz[68][494] = 9'b111111111;
assign micromatrizz[68][495] = 9'b111111111;
assign micromatrizz[68][496] = 9'b111111111;
assign micromatrizz[68][497] = 9'b111111111;
assign micromatrizz[68][498] = 9'b111111111;
assign micromatrizz[68][499] = 9'b111111111;
assign micromatrizz[68][500] = 9'b111110111;
assign micromatrizz[68][501] = 9'b111110010;
assign micromatrizz[68][502] = 9'b111110010;
assign micromatrizz[68][503] = 9'b111110111;
assign micromatrizz[68][504] = 9'b111111111;
assign micromatrizz[68][505] = 9'b111111111;
assign micromatrizz[68][506] = 9'b111111111;
assign micromatrizz[68][507] = 9'b111111111;
assign micromatrizz[68][508] = 9'b111111111;
assign micromatrizz[68][509] = 9'b111110110;
assign micromatrizz[68][510] = 9'b111111111;
assign micromatrizz[68][511] = 9'b111111111;
assign micromatrizz[68][512] = 9'b111111111;
assign micromatrizz[68][513] = 9'b111111111;
assign micromatrizz[68][514] = 9'b111111111;
assign micromatrizz[68][515] = 9'b111111111;
assign micromatrizz[68][516] = 9'b111110110;
assign micromatrizz[68][517] = 9'b111110010;
assign micromatrizz[68][518] = 9'b111110011;
assign micromatrizz[68][519] = 9'b111110011;
assign micromatrizz[68][520] = 9'b111110010;
assign micromatrizz[68][521] = 9'b111110011;
assign micromatrizz[68][522] = 9'b111110011;
assign micromatrizz[68][523] = 9'b111110011;
assign micromatrizz[68][524] = 9'b111110111;
assign micromatrizz[68][525] = 9'b111110111;
assign micromatrizz[68][526] = 9'b111111111;
assign micromatrizz[68][527] = 9'b111111111;
assign micromatrizz[68][528] = 9'b111110111;
assign micromatrizz[68][529] = 9'b111110010;
assign micromatrizz[68][530] = 9'b111110010;
assign micromatrizz[68][531] = 9'b111110010;
assign micromatrizz[68][532] = 9'b111110111;
assign micromatrizz[68][533] = 9'b111111111;
assign micromatrizz[68][534] = 9'b111111111;
assign micromatrizz[68][535] = 9'b111111111;
assign micromatrizz[68][536] = 9'b111111111;
assign micromatrizz[68][537] = 9'b111111111;
assign micromatrizz[68][538] = 9'b111111111;
assign micromatrizz[68][539] = 9'b111111111;
assign micromatrizz[68][540] = 9'b111111111;
assign micromatrizz[68][541] = 9'b111111111;
assign micromatrizz[68][542] = 9'b111110010;
assign micromatrizz[68][543] = 9'b111110010;
assign micromatrizz[68][544] = 9'b111110010;
assign micromatrizz[68][545] = 9'b111110111;
assign micromatrizz[68][546] = 9'b111111111;
assign micromatrizz[68][547] = 9'b111111111;
assign micromatrizz[68][548] = 9'b111111111;
assign micromatrizz[68][549] = 9'b111111111;
assign micromatrizz[68][550] = 9'b111110111;
assign micromatrizz[68][551] = 9'b111110110;
assign micromatrizz[68][552] = 9'b111111111;
assign micromatrizz[68][553] = 9'b111111111;
assign micromatrizz[68][554] = 9'b111111111;
assign micromatrizz[68][555] = 9'b111111111;
assign micromatrizz[68][556] = 9'b111111111;
assign micromatrizz[68][557] = 9'b111111111;
assign micromatrizz[68][558] = 9'b111110010;
assign micromatrizz[68][559] = 9'b111110010;
assign micromatrizz[68][560] = 9'b111110010;
assign micromatrizz[68][561] = 9'b111110011;
assign micromatrizz[68][562] = 9'b111110011;
assign micromatrizz[68][563] = 9'b111110011;
assign micromatrizz[68][564] = 9'b111110010;
assign micromatrizz[68][565] = 9'b111111111;
assign micromatrizz[68][566] = 9'b111111111;
assign micromatrizz[68][567] = 9'b111111111;
assign micromatrizz[68][568] = 9'b111111111;
assign micromatrizz[68][569] = 9'b111111111;
assign micromatrizz[68][570] = 9'b111111111;
assign micromatrizz[68][571] = 9'b111110111;
assign micromatrizz[68][572] = 9'b111110010;
assign micromatrizz[68][573] = 9'b111110010;
assign micromatrizz[68][574] = 9'b111110011;
assign micromatrizz[68][575] = 9'b111110011;
assign micromatrizz[68][576] = 9'b111110111;
assign micromatrizz[68][577] = 9'b111111111;
assign micromatrizz[68][578] = 9'b111110110;
assign micromatrizz[68][579] = 9'b111110111;
assign micromatrizz[68][580] = 9'b111110111;
assign micromatrizz[68][581] = 9'b111110010;
assign micromatrizz[68][582] = 9'b111110010;
assign micromatrizz[68][583] = 9'b111110010;
assign micromatrizz[68][584] = 9'b111110011;
assign micromatrizz[68][585] = 9'b111110011;
assign micromatrizz[68][586] = 9'b111110011;
assign micromatrizz[68][587] = 9'b111110010;
assign micromatrizz[68][588] = 9'b111111111;
assign micromatrizz[68][589] = 9'b111111111;
assign micromatrizz[68][590] = 9'b111111111;
assign micromatrizz[68][591] = 9'b111111111;
assign micromatrizz[68][592] = 9'b111111111;
assign micromatrizz[68][593] = 9'b111111111;
assign micromatrizz[68][594] = 9'b111111111;
assign micromatrizz[68][595] = 9'b111110011;
assign micromatrizz[68][596] = 9'b111110010;
assign micromatrizz[68][597] = 9'b111110010;
assign micromatrizz[68][598] = 9'b111111111;
assign micromatrizz[68][599] = 9'b111111111;
assign micromatrizz[68][600] = 9'b111111111;
assign micromatrizz[68][601] = 9'b111111111;
assign micromatrizz[68][602] = 9'b111111111;
assign micromatrizz[68][603] = 9'b111110111;
assign micromatrizz[68][604] = 9'b111110111;
assign micromatrizz[68][605] = 9'b111111111;
assign micromatrizz[68][606] = 9'b111111111;
assign micromatrizz[68][607] = 9'b111111111;
assign micromatrizz[68][608] = 9'b111111111;
assign micromatrizz[68][609] = 9'b111111111;
assign micromatrizz[68][610] = 9'b111111111;
assign micromatrizz[68][611] = 9'b111110110;
assign micromatrizz[68][612] = 9'b111110111;
assign micromatrizz[68][613] = 9'b111111111;
assign micromatrizz[68][614] = 9'b111111111;
assign micromatrizz[68][615] = 9'b111111111;
assign micromatrizz[68][616] = 9'b111111111;
assign micromatrizz[68][617] = 9'b111110011;
assign micromatrizz[68][618] = 9'b111110010;
assign micromatrizz[68][619] = 9'b111110010;
assign micromatrizz[68][620] = 9'b111110010;
assign micromatrizz[68][621] = 9'b111110111;
assign micromatrizz[68][622] = 9'b111111111;
assign micromatrizz[68][623] = 9'b111111111;
assign micromatrizz[68][624] = 9'b111111111;
assign micromatrizz[68][625] = 9'b111111111;
assign micromatrizz[68][626] = 9'b111111111;
assign micromatrizz[68][627] = 9'b111111111;
assign micromatrizz[68][628] = 9'b111111111;
assign micromatrizz[68][629] = 9'b111111111;
assign micromatrizz[68][630] = 9'b111111111;
assign micromatrizz[68][631] = 9'b111111111;
assign micromatrizz[68][632] = 9'b111111111;
assign micromatrizz[68][633] = 9'b111111111;
assign micromatrizz[68][634] = 9'b111111111;
assign micromatrizz[68][635] = 9'b111111111;
assign micromatrizz[68][636] = 9'b111111111;
assign micromatrizz[68][637] = 9'b111111111;
assign micromatrizz[68][638] = 9'b111111111;
assign micromatrizz[68][639] = 9'b111111111;
assign micromatrizz[69][0] = 9'b111111111;
assign micromatrizz[69][1] = 9'b111111111;
assign micromatrizz[69][2] = 9'b111111111;
assign micromatrizz[69][3] = 9'b111111111;
assign micromatrizz[69][4] = 9'b111111111;
assign micromatrizz[69][5] = 9'b111111111;
assign micromatrizz[69][6] = 9'b111111111;
assign micromatrizz[69][7] = 9'b111111111;
assign micromatrizz[69][8] = 9'b111111111;
assign micromatrizz[69][9] = 9'b111111111;
assign micromatrizz[69][10] = 9'b111111111;
assign micromatrizz[69][11] = 9'b111110111;
assign micromatrizz[69][12] = 9'b111110111;
assign micromatrizz[69][13] = 9'b111111111;
assign micromatrizz[69][14] = 9'b111110111;
assign micromatrizz[69][15] = 9'b111110010;
assign micromatrizz[69][16] = 9'b111110111;
assign micromatrizz[69][17] = 9'b111111111;
assign micromatrizz[69][18] = 9'b111111111;
assign micromatrizz[69][19] = 9'b111111111;
assign micromatrizz[69][20] = 9'b111111111;
assign micromatrizz[69][21] = 9'b111111111;
assign micromatrizz[69][22] = 9'b111111111;
assign micromatrizz[69][23] = 9'b111111111;
assign micromatrizz[69][24] = 9'b111111111;
assign micromatrizz[69][25] = 9'b111111111;
assign micromatrizz[69][26] = 9'b111110111;
assign micromatrizz[69][27] = 9'b111110010;
assign micromatrizz[69][28] = 9'b111110010;
assign micromatrizz[69][29] = 9'b111110011;
assign micromatrizz[69][30] = 9'b111110010;
assign micromatrizz[69][31] = 9'b111110011;
assign micromatrizz[69][32] = 9'b111110111;
assign micromatrizz[69][33] = 9'b111111111;
assign micromatrizz[69][34] = 9'b111111111;
assign micromatrizz[69][35] = 9'b111110111;
assign micromatrizz[69][36] = 9'b111110010;
assign micromatrizz[69][37] = 9'b111110010;
assign micromatrizz[69][38] = 9'b111110010;
assign micromatrizz[69][39] = 9'b111110010;
assign micromatrizz[69][40] = 9'b111110010;
assign micromatrizz[69][41] = 9'b111110010;
assign micromatrizz[69][42] = 9'b111110010;
assign micromatrizz[69][43] = 9'b111111111;
assign micromatrizz[69][44] = 9'b111111111;
assign micromatrizz[69][45] = 9'b111111111;
assign micromatrizz[69][46] = 9'b111111111;
assign micromatrizz[69][47] = 9'b111110010;
assign micromatrizz[69][48] = 9'b111110011;
assign micromatrizz[69][49] = 9'b111110011;
assign micromatrizz[69][50] = 9'b111110011;
assign micromatrizz[69][51] = 9'b111110011;
assign micromatrizz[69][52] = 9'b111110010;
assign micromatrizz[69][53] = 9'b111110010;
assign micromatrizz[69][54] = 9'b111110111;
assign micromatrizz[69][55] = 9'b111111111;
assign micromatrizz[69][56] = 9'b111111111;
assign micromatrizz[69][57] = 9'b111111111;
assign micromatrizz[69][58] = 9'b111111111;
assign micromatrizz[69][59] = 9'b111111111;
assign micromatrizz[69][60] = 9'b111111111;
assign micromatrizz[69][61] = 9'b111111111;
assign micromatrizz[69][62] = 9'b111111111;
assign micromatrizz[69][63] = 9'b111111111;
assign micromatrizz[69][64] = 9'b111111111;
assign micromatrizz[69][65] = 9'b111111111;
assign micromatrizz[69][66] = 9'b111111111;
assign micromatrizz[69][67] = 9'b111111111;
assign micromatrizz[69][68] = 9'b111111111;
assign micromatrizz[69][69] = 9'b111111111;
assign micromatrizz[69][70] = 9'b111111111;
assign micromatrizz[69][71] = 9'b111111111;
assign micromatrizz[69][72] = 9'b111111111;
assign micromatrizz[69][73] = 9'b111111111;
assign micromatrizz[69][74] = 9'b111110011;
assign micromatrizz[69][75] = 9'b111110010;
assign micromatrizz[69][76] = 9'b111111111;
assign micromatrizz[69][77] = 9'b111111111;
assign micromatrizz[69][78] = 9'b111110111;
assign micromatrizz[69][79] = 9'b111110111;
assign micromatrizz[69][80] = 9'b111111111;
assign micromatrizz[69][81] = 9'b111111111;
assign micromatrizz[69][82] = 9'b111111111;
assign micromatrizz[69][83] = 9'b111111111;
assign micromatrizz[69][84] = 9'b111111111;
assign micromatrizz[69][85] = 9'b111111111;
assign micromatrizz[69][86] = 9'b111111111;
assign micromatrizz[69][87] = 9'b111111111;
assign micromatrizz[69][88] = 9'b111110010;
assign micromatrizz[69][89] = 9'b111110010;
assign micromatrizz[69][90] = 9'b111110010;
assign micromatrizz[69][91] = 9'b111110010;
assign micromatrizz[69][92] = 9'b111110010;
assign micromatrizz[69][93] = 9'b111110010;
assign micromatrizz[69][94] = 9'b111110010;
assign micromatrizz[69][95] = 9'b111110111;
assign micromatrizz[69][96] = 9'b111111111;
assign micromatrizz[69][97] = 9'b111111111;
assign micromatrizz[69][98] = 9'b111111111;
assign micromatrizz[69][99] = 9'b111111111;
assign micromatrizz[69][100] = 9'b111111111;
assign micromatrizz[69][101] = 9'b111111111;
assign micromatrizz[69][102] = 9'b111111111;
assign micromatrizz[69][103] = 9'b111111111;
assign micromatrizz[69][104] = 9'b111111111;
assign micromatrizz[69][105] = 9'b111111111;
assign micromatrizz[69][106] = 9'b111111111;
assign micromatrizz[69][107] = 9'b111110111;
assign micromatrizz[69][108] = 9'b111110111;
assign micromatrizz[69][109] = 9'b111111111;
assign micromatrizz[69][110] = 9'b111110111;
assign micromatrizz[69][111] = 9'b111110010;
assign micromatrizz[69][112] = 9'b111110010;
assign micromatrizz[69][113] = 9'b111110111;
assign micromatrizz[69][114] = 9'b111111111;
assign micromatrizz[69][115] = 9'b111111111;
assign micromatrizz[69][116] = 9'b111111111;
assign micromatrizz[69][117] = 9'b111111111;
assign micromatrizz[69][118] = 9'b111111111;
assign micromatrizz[69][119] = 9'b111111111;
assign micromatrizz[69][120] = 9'b111111111;
assign micromatrizz[69][121] = 9'b111111111;
assign micromatrizz[69][122] = 9'b111111111;
assign micromatrizz[69][123] = 9'b111111111;
assign micromatrizz[69][124] = 9'b111110111;
assign micromatrizz[69][125] = 9'b111110010;
assign micromatrizz[69][126] = 9'b111110010;
assign micromatrizz[69][127] = 9'b111110111;
assign micromatrizz[69][128] = 9'b111111111;
assign micromatrizz[69][129] = 9'b111110111;
assign micromatrizz[69][130] = 9'b111110111;
assign micromatrizz[69][131] = 9'b111111111;
assign micromatrizz[69][132] = 9'b111111111;
assign micromatrizz[69][133] = 9'b111111111;
assign micromatrizz[69][134] = 9'b111111111;
assign micromatrizz[69][135] = 9'b111111111;
assign micromatrizz[69][136] = 9'b111111111;
assign micromatrizz[69][137] = 9'b111111111;
assign micromatrizz[69][138] = 9'b111110111;
assign micromatrizz[69][139] = 9'b111110010;
assign micromatrizz[69][140] = 9'b111110010;
assign micromatrizz[69][141] = 9'b111110010;
assign micromatrizz[69][142] = 9'b111110010;
assign micromatrizz[69][143] = 9'b111110010;
assign micromatrizz[69][144] = 9'b111110010;
assign micromatrizz[69][145] = 9'b111110011;
assign micromatrizz[69][146] = 9'b111111111;
assign micromatrizz[69][147] = 9'b111111111;
assign micromatrizz[69][148] = 9'b111111111;
assign micromatrizz[69][149] = 9'b111111111;
assign micromatrizz[69][150] = 9'b111110110;
assign micromatrizz[69][151] = 9'b111110010;
assign micromatrizz[69][152] = 9'b111110010;
assign micromatrizz[69][153] = 9'b111110010;
assign micromatrizz[69][154] = 9'b111110010;
assign micromatrizz[69][155] = 9'b111110010;
assign micromatrizz[69][156] = 9'b111110010;
assign micromatrizz[69][157] = 9'b111110011;
assign micromatrizz[69][158] = 9'b111111111;
assign micromatrizz[69][159] = 9'b111111111;
assign micromatrizz[69][160] = 9'b111111111;
assign micromatrizz[69][161] = 9'b111111111;
assign micromatrizz[69][162] = 9'b111111111;
assign micromatrizz[69][163] = 9'b111111111;
assign micromatrizz[69][164] = 9'b111110011;
assign micromatrizz[69][165] = 9'b111110010;
assign micromatrizz[69][166] = 9'b111110010;
assign micromatrizz[69][167] = 9'b111110011;
assign micromatrizz[69][168] = 9'b111110011;
assign micromatrizz[69][169] = 9'b111110111;
assign micromatrizz[69][170] = 9'b111111111;
assign micromatrizz[69][171] = 9'b111111111;
assign micromatrizz[69][172] = 9'b111110010;
assign micromatrizz[69][173] = 9'b111110010;
assign micromatrizz[69][174] = 9'b111110010;
assign micromatrizz[69][175] = 9'b111110010;
assign micromatrizz[69][176] = 9'b111110010;
assign micromatrizz[69][177] = 9'b111110010;
assign micromatrizz[69][178] = 9'b111110010;
assign micromatrizz[69][179] = 9'b111110010;
assign micromatrizz[69][180] = 9'b111111111;
assign micromatrizz[69][181] = 9'b111111111;
assign micromatrizz[69][182] = 9'b111111111;
assign micromatrizz[69][183] = 9'b111111111;
assign micromatrizz[69][184] = 9'b111111111;
assign micromatrizz[69][185] = 9'b111111111;
assign micromatrizz[69][186] = 9'b111111111;
assign micromatrizz[69][187] = 9'b111110111;
assign micromatrizz[69][188] = 9'b111110011;
assign micromatrizz[69][189] = 9'b111110011;
assign micromatrizz[69][190] = 9'b111110010;
assign micromatrizz[69][191] = 9'b111110010;
assign micromatrizz[69][192] = 9'b111110111;
assign micromatrizz[69][193] = 9'b111111111;
assign micromatrizz[69][194] = 9'b111111111;
assign micromatrizz[69][195] = 9'b111110010;
assign micromatrizz[69][196] = 9'b111110010;
assign micromatrizz[69][197] = 9'b111110010;
assign micromatrizz[69][198] = 9'b111110010;
assign micromatrizz[69][199] = 9'b111110010;
assign micromatrizz[69][200] = 9'b111110010;
assign micromatrizz[69][201] = 9'b111110010;
assign micromatrizz[69][202] = 9'b111110111;
assign micromatrizz[69][203] = 9'b111111111;
assign micromatrizz[69][204] = 9'b111111111;
assign micromatrizz[69][205] = 9'b111111111;
assign micromatrizz[69][206] = 9'b111111111;
assign micromatrizz[69][207] = 9'b111111111;
assign micromatrizz[69][208] = 9'b111111111;
assign micromatrizz[69][209] = 9'b111111111;
assign micromatrizz[69][210] = 9'b111111111;
assign micromatrizz[69][211] = 9'b111110111;
assign micromatrizz[69][212] = 9'b111110010;
assign micromatrizz[69][213] = 9'b111110011;
assign micromatrizz[69][214] = 9'b111111111;
assign micromatrizz[69][215] = 9'b111110111;
assign micromatrizz[69][216] = 9'b111110111;
assign micromatrizz[69][217] = 9'b111111111;
assign micromatrizz[69][218] = 9'b111111111;
assign micromatrizz[69][219] = 9'b111111111;
assign micromatrizz[69][220] = 9'b111111111;
assign micromatrizz[69][221] = 9'b111111111;
assign micromatrizz[69][222] = 9'b111111111;
assign micromatrizz[69][223] = 9'b111111111;
assign micromatrizz[69][224] = 9'b111111111;
assign micromatrizz[69][225] = 9'b111110010;
assign micromatrizz[69][226] = 9'b111110010;
assign micromatrizz[69][227] = 9'b111110010;
assign micromatrizz[69][228] = 9'b111110010;
assign micromatrizz[69][229] = 9'b111110010;
assign micromatrizz[69][230] = 9'b111110011;
assign micromatrizz[69][231] = 9'b111110010;
assign micromatrizz[69][232] = 9'b111110111;
assign micromatrizz[69][233] = 9'b111111111;
assign micromatrizz[69][234] = 9'b111111111;
assign micromatrizz[69][235] = 9'b111111111;
assign micromatrizz[69][236] = 9'b111111111;
assign micromatrizz[69][237] = 9'b111111111;
assign micromatrizz[69][238] = 9'b111111111;
assign micromatrizz[69][239] = 9'b111111111;
assign micromatrizz[69][240] = 9'b111111111;
assign micromatrizz[69][241] = 9'b111111111;
assign micromatrizz[69][242] = 9'b111111111;
assign micromatrizz[69][243] = 9'b111111111;
assign micromatrizz[69][244] = 9'b111111111;
assign micromatrizz[69][245] = 9'b111111111;
assign micromatrizz[69][246] = 9'b111110111;
assign micromatrizz[69][247] = 9'b111110010;
assign micromatrizz[69][248] = 9'b111110111;
assign micromatrizz[69][249] = 9'b111111111;
assign micromatrizz[69][250] = 9'b111111111;
assign micromatrizz[69][251] = 9'b111110111;
assign micromatrizz[69][252] = 9'b111110111;
assign micromatrizz[69][253] = 9'b111111111;
assign micromatrizz[69][254] = 9'b111111111;
assign micromatrizz[69][255] = 9'b111111111;
assign micromatrizz[69][256] = 9'b111111111;
assign micromatrizz[69][257] = 9'b111111111;
assign micromatrizz[69][258] = 9'b111111111;
assign micromatrizz[69][259] = 9'b111111111;
assign micromatrizz[69][260] = 9'b111111111;
assign micromatrizz[69][261] = 9'b111111111;
assign micromatrizz[69][262] = 9'b111110111;
assign micromatrizz[69][263] = 9'b111110111;
assign micromatrizz[69][264] = 9'b111110111;
assign micromatrizz[69][265] = 9'b111111111;
assign micromatrizz[69][266] = 9'b111110111;
assign micromatrizz[69][267] = 9'b111110010;
assign micromatrizz[69][268] = 9'b111110111;
assign micromatrizz[69][269] = 9'b111111111;
assign micromatrizz[69][270] = 9'b111111111;
assign micromatrizz[69][271] = 9'b111111111;
assign micromatrizz[69][272] = 9'b111111111;
assign micromatrizz[69][273] = 9'b111111111;
assign micromatrizz[69][274] = 9'b111111111;
assign micromatrizz[69][275] = 9'b111111111;
assign micromatrizz[69][276] = 9'b111111111;
assign micromatrizz[69][277] = 9'b111111111;
assign micromatrizz[69][278] = 9'b111110111;
assign micromatrizz[69][279] = 9'b111110010;
assign micromatrizz[69][280] = 9'b111110010;
assign micromatrizz[69][281] = 9'b111110010;
assign micromatrizz[69][282] = 9'b111110011;
assign micromatrizz[69][283] = 9'b111110111;
assign micromatrizz[69][284] = 9'b111111111;
assign micromatrizz[69][285] = 9'b111111111;
assign micromatrizz[69][286] = 9'b111110010;
assign micromatrizz[69][287] = 9'b111110010;
assign micromatrizz[69][288] = 9'b111110010;
assign micromatrizz[69][289] = 9'b111110010;
assign micromatrizz[69][290] = 9'b111110010;
assign micromatrizz[69][291] = 9'b111110010;
assign micromatrizz[69][292] = 9'b111110010;
assign micromatrizz[69][293] = 9'b111110010;
assign micromatrizz[69][294] = 9'b111111111;
assign micromatrizz[69][295] = 9'b111111111;
assign micromatrizz[69][296] = 9'b111111111;
assign micromatrizz[69][297] = 9'b111111111;
assign micromatrizz[69][298] = 9'b111111111;
assign micromatrizz[69][299] = 9'b111111111;
assign micromatrizz[69][300] = 9'b111111111;
assign micromatrizz[69][301] = 9'b111111111;
assign micromatrizz[69][302] = 9'b111111111;
assign micromatrizz[69][303] = 9'b111111111;
assign micromatrizz[69][304] = 9'b111111111;
assign micromatrizz[69][305] = 9'b111110111;
assign micromatrizz[69][306] = 9'b111111111;
assign micromatrizz[69][307] = 9'b111111111;
assign micromatrizz[69][308] = 9'b111111111;
assign micromatrizz[69][309] = 9'b111111111;
assign micromatrizz[69][310] = 9'b111111111;
assign micromatrizz[69][311] = 9'b111111111;
assign micromatrizz[69][312] = 9'b111111111;
assign micromatrizz[69][313] = 9'b111111111;
assign micromatrizz[69][314] = 9'b111111111;
assign micromatrizz[69][315] = 9'b111111111;
assign micromatrizz[69][316] = 9'b111111111;
assign micromatrizz[69][317] = 9'b111111111;
assign micromatrizz[69][318] = 9'b111111111;
assign micromatrizz[69][319] = 9'b111111111;
assign micromatrizz[69][320] = 9'b111110111;
assign micromatrizz[69][321] = 9'b111110011;
assign micromatrizz[69][322] = 9'b111110010;
assign micromatrizz[69][323] = 9'b111111111;
assign micromatrizz[69][324] = 9'b111111111;
assign micromatrizz[69][325] = 9'b111111111;
assign micromatrizz[69][326] = 9'b111110111;
assign micromatrizz[69][327] = 9'b111111111;
assign micromatrizz[69][328] = 9'b111111111;
assign micromatrizz[69][329] = 9'b111111111;
assign micromatrizz[69][330] = 9'b111111111;
assign micromatrizz[69][331] = 9'b111111111;
assign micromatrizz[69][332] = 9'b111111111;
assign micromatrizz[69][333] = 9'b111111111;
assign micromatrizz[69][334] = 9'b111111111;
assign micromatrizz[69][335] = 9'b111110010;
assign micromatrizz[69][336] = 9'b111110010;
assign micromatrizz[69][337] = 9'b111110011;
assign micromatrizz[69][338] = 9'b111110010;
assign micromatrizz[69][339] = 9'b111110010;
assign micromatrizz[69][340] = 9'b111110010;
assign micromatrizz[69][341] = 9'b111110010;
assign micromatrizz[69][342] = 9'b111110111;
assign micromatrizz[69][343] = 9'b111111111;
assign micromatrizz[69][344] = 9'b111111111;
assign micromatrizz[69][345] = 9'b111111111;
assign micromatrizz[69][346] = 9'b111111111;
assign micromatrizz[69][347] = 9'b111110010;
assign micromatrizz[69][348] = 9'b111110010;
assign micromatrizz[69][349] = 9'b111110010;
assign micromatrizz[69][350] = 9'b111110010;
assign micromatrizz[69][351] = 9'b111110010;
assign micromatrizz[69][352] = 9'b111110010;
assign micromatrizz[69][353] = 9'b111110010;
assign micromatrizz[69][354] = 9'b111111111;
assign micromatrizz[69][355] = 9'b111111111;
assign micromatrizz[69][356] = 9'b111111111;
assign micromatrizz[69][357] = 9'b111111111;
assign micromatrizz[69][358] = 9'b111111111;
assign micromatrizz[69][359] = 9'b111111111;
assign micromatrizz[69][360] = 9'b111111111;
assign micromatrizz[69][361] = 9'b111110111;
assign micromatrizz[69][362] = 9'b111110010;
assign micromatrizz[69][363] = 9'b111110010;
assign micromatrizz[69][364] = 9'b111110010;
assign micromatrizz[69][365] = 9'b111110010;
assign micromatrizz[69][366] = 9'b111110111;
assign micromatrizz[69][367] = 9'b111111111;
assign micromatrizz[69][368] = 9'b111111111;
assign micromatrizz[69][369] = 9'b111111111;
assign micromatrizz[69][370] = 9'b111111111;
assign micromatrizz[69][371] = 9'b111111111;
assign micromatrizz[69][372] = 9'b111111111;
assign micromatrizz[69][373] = 9'b111111111;
assign micromatrizz[69][374] = 9'b111110111;
assign micromatrizz[69][375] = 9'b111110011;
assign micromatrizz[69][376] = 9'b111110010;
assign micromatrizz[69][377] = 9'b111110010;
assign micromatrizz[69][378] = 9'b111110010;
assign micromatrizz[69][379] = 9'b111110011;
assign micromatrizz[69][380] = 9'b111110111;
assign micromatrizz[69][381] = 9'b111111111;
assign micromatrizz[69][382] = 9'b111111111;
assign micromatrizz[69][383] = 9'b111110111;
assign micromatrizz[69][384] = 9'b111110010;
assign micromatrizz[69][385] = 9'b111110010;
assign micromatrizz[69][386] = 9'b111110010;
assign micromatrizz[69][387] = 9'b111110010;
assign micromatrizz[69][388] = 9'b111110010;
assign micromatrizz[69][389] = 9'b111110010;
assign micromatrizz[69][390] = 9'b111110010;
assign micromatrizz[69][391] = 9'b111111111;
assign micromatrizz[69][392] = 9'b111111111;
assign micromatrizz[69][393] = 9'b111111111;
assign micromatrizz[69][394] = 9'b111111111;
assign micromatrizz[69][395] = 9'b111110110;
assign micromatrizz[69][396] = 9'b111110010;
assign micromatrizz[69][397] = 9'b111110010;
assign micromatrizz[69][398] = 9'b111110010;
assign micromatrizz[69][399] = 9'b111110010;
assign micromatrizz[69][400] = 9'b111110010;
assign micromatrizz[69][401] = 9'b111110010;
assign micromatrizz[69][402] = 9'b111110111;
assign micromatrizz[69][403] = 9'b111111111;
assign micromatrizz[69][404] = 9'b111111111;
assign micromatrizz[69][405] = 9'b111111111;
assign micromatrizz[69][406] = 9'b111111111;
assign micromatrizz[69][407] = 9'b111111111;
assign micromatrizz[69][408] = 9'b111111111;
assign micromatrizz[69][409] = 9'b111111111;
assign micromatrizz[69][410] = 9'b111111111;
assign micromatrizz[69][411] = 9'b111111111;
assign micromatrizz[69][412] = 9'b111111111;
assign micromatrizz[69][413] = 9'b111111111;
assign micromatrizz[69][414] = 9'b111111111;
assign micromatrizz[69][415] = 9'b111111111;
assign micromatrizz[69][416] = 9'b111110111;
assign micromatrizz[69][417] = 9'b111110010;
assign micromatrizz[69][418] = 9'b111110111;
assign micromatrizz[69][419] = 9'b111111111;
assign micromatrizz[69][420] = 9'b111111111;
assign micromatrizz[69][421] = 9'b111110111;
assign micromatrizz[69][422] = 9'b111110111;
assign micromatrizz[69][423] = 9'b111111111;
assign micromatrizz[69][424] = 9'b111111111;
assign micromatrizz[69][425] = 9'b111111111;
assign micromatrizz[69][426] = 9'b111111111;
assign micromatrizz[69][427] = 9'b111111111;
assign micromatrizz[69][428] = 9'b111111111;
assign micromatrizz[69][429] = 9'b111111111;
assign micromatrizz[69][430] = 9'b111110111;
assign micromatrizz[69][431] = 9'b111110010;
assign micromatrizz[69][432] = 9'b111110010;
assign micromatrizz[69][433] = 9'b111110010;
assign micromatrizz[69][434] = 9'b111110010;
assign micromatrizz[69][435] = 9'b111110010;
assign micromatrizz[69][436] = 9'b111110010;
assign micromatrizz[69][437] = 9'b111110111;
assign micromatrizz[69][438] = 9'b111111111;
assign micromatrizz[69][439] = 9'b111111111;
assign micromatrizz[69][440] = 9'b111111111;
assign micromatrizz[69][441] = 9'b111111111;
assign micromatrizz[69][442] = 9'b111111111;
assign micromatrizz[69][443] = 9'b111111111;
assign micromatrizz[69][444] = 9'b111111111;
assign micromatrizz[69][445] = 9'b111111111;
assign micromatrizz[69][446] = 9'b111111111;
assign micromatrizz[69][447] = 9'b111111111;
assign micromatrizz[69][448] = 9'b111111111;
assign micromatrizz[69][449] = 9'b111111111;
assign micromatrizz[69][450] = 9'b111111111;
assign micromatrizz[69][451] = 9'b111110111;
assign micromatrizz[69][452] = 9'b111110011;
assign micromatrizz[69][453] = 9'b111110010;
assign micromatrizz[69][454] = 9'b111110111;
assign micromatrizz[69][455] = 9'b111111111;
assign micromatrizz[69][456] = 9'b111110111;
assign micromatrizz[69][457] = 9'b111110111;
assign micromatrizz[69][458] = 9'b111111111;
assign micromatrizz[69][459] = 9'b111111111;
assign micromatrizz[69][460] = 9'b111111111;
assign micromatrizz[69][461] = 9'b111111111;
assign micromatrizz[69][462] = 9'b111111111;
assign micromatrizz[69][463] = 9'b111111111;
assign micromatrizz[69][464] = 9'b111111111;
assign micromatrizz[69][465] = 9'b111111111;
assign micromatrizz[69][466] = 9'b111111111;
assign micromatrizz[69][467] = 9'b111110111;
assign micromatrizz[69][468] = 9'b111110111;
assign micromatrizz[69][469] = 9'b111111111;
assign micromatrizz[69][470] = 9'b111111111;
assign micromatrizz[69][471] = 9'b111110111;
assign micromatrizz[69][472] = 9'b111110010;
assign micromatrizz[69][473] = 9'b111110010;
assign micromatrizz[69][474] = 9'b111110111;
assign micromatrizz[69][475] = 9'b111111111;
assign micromatrizz[69][476] = 9'b111111111;
assign micromatrizz[69][477] = 9'b111111111;
assign micromatrizz[69][478] = 9'b111111111;
assign micromatrizz[69][479] = 9'b111111111;
assign micromatrizz[69][480] = 9'b111111111;
assign micromatrizz[69][481] = 9'b111110010;
assign micromatrizz[69][482] = 9'b111110010;
assign micromatrizz[69][483] = 9'b111110010;
assign micromatrizz[69][484] = 9'b111110010;
assign micromatrizz[69][485] = 9'b111110010;
assign micromatrizz[69][486] = 9'b111110010;
assign micromatrizz[69][487] = 9'b111110010;
assign micromatrizz[69][488] = 9'b111110111;
assign micromatrizz[69][489] = 9'b111111111;
assign micromatrizz[69][490] = 9'b111111111;
assign micromatrizz[69][491] = 9'b111111111;
assign micromatrizz[69][492] = 9'b111111111;
assign micromatrizz[69][493] = 9'b111111111;
assign micromatrizz[69][494] = 9'b111111111;
assign micromatrizz[69][495] = 9'b111111111;
assign micromatrizz[69][496] = 9'b111111111;
assign micromatrizz[69][497] = 9'b111111111;
assign micromatrizz[69][498] = 9'b111111111;
assign micromatrizz[69][499] = 9'b111111111;
assign micromatrizz[69][500] = 9'b111111111;
assign micromatrizz[69][501] = 9'b111111111;
assign micromatrizz[69][502] = 9'b111110111;
assign micromatrizz[69][503] = 9'b111110010;
assign micromatrizz[69][504] = 9'b111110111;
assign micromatrizz[69][505] = 9'b111111111;
assign micromatrizz[69][506] = 9'b111110111;
assign micromatrizz[69][507] = 9'b111110111;
assign micromatrizz[69][508] = 9'b111111111;
assign micromatrizz[69][509] = 9'b111111111;
assign micromatrizz[69][510] = 9'b111111111;
assign micromatrizz[69][511] = 9'b111111111;
assign micromatrizz[69][512] = 9'b111111111;
assign micromatrizz[69][513] = 9'b111111111;
assign micromatrizz[69][514] = 9'b111111111;
assign micromatrizz[69][515] = 9'b111111111;
assign micromatrizz[69][516] = 9'b111110110;
assign micromatrizz[69][517] = 9'b111110010;
assign micromatrizz[69][518] = 9'b111110011;
assign micromatrizz[69][519] = 9'b111110010;
assign micromatrizz[69][520] = 9'b111110010;
assign micromatrizz[69][521] = 9'b111110010;
assign micromatrizz[69][522] = 9'b111110010;
assign micromatrizz[69][523] = 9'b111110111;
assign micromatrizz[69][524] = 9'b111111111;
assign micromatrizz[69][525] = 9'b111111111;
assign micromatrizz[69][526] = 9'b111110111;
assign micromatrizz[69][527] = 9'b111110010;
assign micromatrizz[69][528] = 9'b111110010;
assign micromatrizz[69][529] = 9'b111110010;
assign micromatrizz[69][530] = 9'b111110010;
assign micromatrizz[69][531] = 9'b111110111;
assign micromatrizz[69][532] = 9'b111111111;
assign micromatrizz[69][533] = 9'b111111111;
assign micromatrizz[69][534] = 9'b111111111;
assign micromatrizz[69][535] = 9'b111111111;
assign micromatrizz[69][536] = 9'b111111111;
assign micromatrizz[69][537] = 9'b111111111;
assign micromatrizz[69][538] = 9'b111111111;
assign micromatrizz[69][539] = 9'b111111111;
assign micromatrizz[69][540] = 9'b111111111;
assign micromatrizz[69][541] = 9'b111111111;
assign micromatrizz[69][542] = 9'b111111111;
assign micromatrizz[69][543] = 9'b111110111;
assign micromatrizz[69][544] = 9'b111110011;
assign micromatrizz[69][545] = 9'b111110011;
assign micromatrizz[69][546] = 9'b111110111;
assign micromatrizz[69][547] = 9'b111111111;
assign micromatrizz[69][548] = 9'b111110111;
assign micromatrizz[69][549] = 9'b111110111;
assign micromatrizz[69][550] = 9'b111111111;
assign micromatrizz[69][551] = 9'b111111111;
assign micromatrizz[69][552] = 9'b111111111;
assign micromatrizz[69][553] = 9'b111111111;
assign micromatrizz[69][554] = 9'b111111111;
assign micromatrizz[69][555] = 9'b111111111;
assign micromatrizz[69][556] = 9'b111111111;
assign micromatrizz[69][557] = 9'b111111111;
assign micromatrizz[69][558] = 9'b111110010;
assign micromatrizz[69][559] = 9'b111110010;
assign micromatrizz[69][560] = 9'b111110010;
assign micromatrizz[69][561] = 9'b111110010;
assign micromatrizz[69][562] = 9'b111110010;
assign micromatrizz[69][563] = 9'b111110010;
assign micromatrizz[69][564] = 9'b111110010;
assign micromatrizz[69][565] = 9'b111111111;
assign micromatrizz[69][566] = 9'b111111111;
assign micromatrizz[69][567] = 9'b111111111;
assign micromatrizz[69][568] = 9'b111111111;
assign micromatrizz[69][569] = 9'b111111111;
assign micromatrizz[69][570] = 9'b111111111;
assign micromatrizz[69][571] = 9'b111111111;
assign micromatrizz[69][572] = 9'b111111111;
assign micromatrizz[69][573] = 9'b111110111;
assign micromatrizz[69][574] = 9'b111110010;
assign micromatrizz[69][575] = 9'b111110010;
assign micromatrizz[69][576] = 9'b111110010;
assign micromatrizz[69][577] = 9'b111110010;
assign micromatrizz[69][578] = 9'b111111111;
assign micromatrizz[69][579] = 9'b111111111;
assign micromatrizz[69][580] = 9'b111111111;
assign micromatrizz[69][581] = 9'b111110010;
assign micromatrizz[69][582] = 9'b111110010;
assign micromatrizz[69][583] = 9'b111110010;
assign micromatrizz[69][584] = 9'b111110010;
assign micromatrizz[69][585] = 9'b111110010;
assign micromatrizz[69][586] = 9'b111110010;
assign micromatrizz[69][587] = 9'b111110010;
assign micromatrizz[69][588] = 9'b111111111;
assign micromatrizz[69][589] = 9'b111111111;
assign micromatrizz[69][590] = 9'b111111111;
assign micromatrizz[69][591] = 9'b111111111;
assign micromatrizz[69][592] = 9'b111111111;
assign micromatrizz[69][593] = 9'b111111111;
assign micromatrizz[69][594] = 9'b111111111;
assign micromatrizz[69][595] = 9'b111111111;
assign micromatrizz[69][596] = 9'b111110111;
assign micromatrizz[69][597] = 9'b111110010;
assign micromatrizz[69][598] = 9'b111110111;
assign micromatrizz[69][599] = 9'b111111111;
assign micromatrizz[69][600] = 9'b111111111;
assign micromatrizz[69][601] = 9'b111110111;
assign micromatrizz[69][602] = 9'b111110111;
assign micromatrizz[69][603] = 9'b111111111;
assign micromatrizz[69][604] = 9'b111111111;
assign micromatrizz[69][605] = 9'b111111111;
assign micromatrizz[69][606] = 9'b111111111;
assign micromatrizz[69][607] = 9'b111111111;
assign micromatrizz[69][608] = 9'b111111111;
assign micromatrizz[69][609] = 9'b111111111;
assign micromatrizz[69][610] = 9'b111111111;
assign micromatrizz[69][611] = 9'b111111111;
assign micromatrizz[69][612] = 9'b111111111;
assign micromatrizz[69][613] = 9'b111110111;
assign micromatrizz[69][614] = 9'b111110111;
assign micromatrizz[69][615] = 9'b111111111;
assign micromatrizz[69][616] = 9'b111111111;
assign micromatrizz[69][617] = 9'b111110010;
assign micromatrizz[69][618] = 9'b111110111;
assign micromatrizz[69][619] = 9'b111110111;
assign micromatrizz[69][620] = 9'b111111111;
assign micromatrizz[69][621] = 9'b111111111;
assign micromatrizz[69][622] = 9'b111111111;
assign micromatrizz[69][623] = 9'b111111111;
assign micromatrizz[69][624] = 9'b111111111;
assign micromatrizz[69][625] = 9'b111111111;
assign micromatrizz[69][626] = 9'b111111111;
assign micromatrizz[69][627] = 9'b111111111;
assign micromatrizz[69][628] = 9'b111111111;
assign micromatrizz[69][629] = 9'b111111111;
assign micromatrizz[69][630] = 9'b111111111;
assign micromatrizz[69][631] = 9'b111111111;
assign micromatrizz[69][632] = 9'b111111111;
assign micromatrizz[69][633] = 9'b111111111;
assign micromatrizz[69][634] = 9'b111111111;
assign micromatrizz[69][635] = 9'b111111111;
assign micromatrizz[69][636] = 9'b111111111;
assign micromatrizz[69][637] = 9'b111111111;
assign micromatrizz[69][638] = 9'b111111111;
assign micromatrizz[69][639] = 9'b111111111;
assign micromatrizz[70][0] = 9'b111111111;
assign micromatrizz[70][1] = 9'b111111111;
assign micromatrizz[70][2] = 9'b111111111;
assign micromatrizz[70][3] = 9'b111111111;
assign micromatrizz[70][4] = 9'b111111111;
assign micromatrizz[70][5] = 9'b111111111;
assign micromatrizz[70][6] = 9'b111111111;
assign micromatrizz[70][7] = 9'b111111111;
assign micromatrizz[70][8] = 9'b111111111;
assign micromatrizz[70][9] = 9'b111111111;
assign micromatrizz[70][10] = 9'b111111111;
assign micromatrizz[70][11] = 9'b111111111;
assign micromatrizz[70][12] = 9'b111111111;
assign micromatrizz[70][13] = 9'b111111111;
assign micromatrizz[70][14] = 9'b111111111;
assign micromatrizz[70][15] = 9'b111111111;
assign micromatrizz[70][16] = 9'b111111111;
assign micromatrizz[70][17] = 9'b111111111;
assign micromatrizz[70][18] = 9'b111111111;
assign micromatrizz[70][19] = 9'b111111111;
assign micromatrizz[70][20] = 9'b111111111;
assign micromatrizz[70][21] = 9'b111111111;
assign micromatrizz[70][22] = 9'b111111111;
assign micromatrizz[70][23] = 9'b111111111;
assign micromatrizz[70][24] = 9'b111111111;
assign micromatrizz[70][25] = 9'b111111111;
assign micromatrizz[70][26] = 9'b111111111;
assign micromatrizz[70][27] = 9'b111111111;
assign micromatrizz[70][28] = 9'b111111111;
assign micromatrizz[70][29] = 9'b111111111;
assign micromatrizz[70][30] = 9'b111111111;
assign micromatrizz[70][31] = 9'b111111111;
assign micromatrizz[70][32] = 9'b111111111;
assign micromatrizz[70][33] = 9'b111111111;
assign micromatrizz[70][34] = 9'b111111111;
assign micromatrizz[70][35] = 9'b111111111;
assign micromatrizz[70][36] = 9'b111111111;
assign micromatrizz[70][37] = 9'b111111111;
assign micromatrizz[70][38] = 9'b111111111;
assign micromatrizz[70][39] = 9'b111111111;
assign micromatrizz[70][40] = 9'b111111111;
assign micromatrizz[70][41] = 9'b111111111;
assign micromatrizz[70][42] = 9'b111111111;
assign micromatrizz[70][43] = 9'b111111111;
assign micromatrizz[70][44] = 9'b111111111;
assign micromatrizz[70][45] = 9'b111111111;
assign micromatrizz[70][46] = 9'b111111111;
assign micromatrizz[70][47] = 9'b111110010;
assign micromatrizz[70][48] = 9'b111110010;
assign micromatrizz[70][49] = 9'b111110010;
assign micromatrizz[70][50] = 9'b111110010;
assign micromatrizz[70][51] = 9'b111110010;
assign micromatrizz[70][52] = 9'b111110010;
assign micromatrizz[70][53] = 9'b111110010;
assign micromatrizz[70][54] = 9'b111110111;
assign micromatrizz[70][55] = 9'b111111111;
assign micromatrizz[70][56] = 9'b111111111;
assign micromatrizz[70][57] = 9'b111111111;
assign micromatrizz[70][58] = 9'b111111111;
assign micromatrizz[70][59] = 9'b111111111;
assign micromatrizz[70][60] = 9'b111111111;
assign micromatrizz[70][61] = 9'b111111111;
assign micromatrizz[70][62] = 9'b111111111;
assign micromatrizz[70][63] = 9'b111111111;
assign micromatrizz[70][64] = 9'b111111111;
assign micromatrizz[70][65] = 9'b111111111;
assign micromatrizz[70][66] = 9'b111111111;
assign micromatrizz[70][67] = 9'b111111111;
assign micromatrizz[70][68] = 9'b111111111;
assign micromatrizz[70][69] = 9'b111111111;
assign micromatrizz[70][70] = 9'b111111111;
assign micromatrizz[70][71] = 9'b111111111;
assign micromatrizz[70][72] = 9'b111111111;
assign micromatrizz[70][73] = 9'b111111111;
assign micromatrizz[70][74] = 9'b111111111;
assign micromatrizz[70][75] = 9'b111111111;
assign micromatrizz[70][76] = 9'b111111111;
assign micromatrizz[70][77] = 9'b111111111;
assign micromatrizz[70][78] = 9'b111111111;
assign micromatrizz[70][79] = 9'b111111111;
assign micromatrizz[70][80] = 9'b111111111;
assign micromatrizz[70][81] = 9'b111111111;
assign micromatrizz[70][82] = 9'b111111111;
assign micromatrizz[70][83] = 9'b111111111;
assign micromatrizz[70][84] = 9'b111111111;
assign micromatrizz[70][85] = 9'b111111111;
assign micromatrizz[70][86] = 9'b111111111;
assign micromatrizz[70][87] = 9'b111111111;
assign micromatrizz[70][88] = 9'b111111111;
assign micromatrizz[70][89] = 9'b111111111;
assign micromatrizz[70][90] = 9'b111111111;
assign micromatrizz[70][91] = 9'b111111111;
assign micromatrizz[70][92] = 9'b111111111;
assign micromatrizz[70][93] = 9'b111111111;
assign micromatrizz[70][94] = 9'b111111111;
assign micromatrizz[70][95] = 9'b111111111;
assign micromatrizz[70][96] = 9'b111111111;
assign micromatrizz[70][97] = 9'b111111111;
assign micromatrizz[70][98] = 9'b111111111;
assign micromatrizz[70][99] = 9'b111111111;
assign micromatrizz[70][100] = 9'b111111111;
assign micromatrizz[70][101] = 9'b111111111;
assign micromatrizz[70][102] = 9'b111111111;
assign micromatrizz[70][103] = 9'b111111111;
assign micromatrizz[70][104] = 9'b111111111;
assign micromatrizz[70][105] = 9'b111111111;
assign micromatrizz[70][106] = 9'b111111111;
assign micromatrizz[70][107] = 9'b111111111;
assign micromatrizz[70][108] = 9'b111111111;
assign micromatrizz[70][109] = 9'b111111111;
assign micromatrizz[70][110] = 9'b111111111;
assign micromatrizz[70][111] = 9'b111111111;
assign micromatrizz[70][112] = 9'b111111111;
assign micromatrizz[70][113] = 9'b111111111;
assign micromatrizz[70][114] = 9'b111111111;
assign micromatrizz[70][115] = 9'b111111111;
assign micromatrizz[70][116] = 9'b111111111;
assign micromatrizz[70][117] = 9'b111111111;
assign micromatrizz[70][118] = 9'b111111111;
assign micromatrizz[70][119] = 9'b111111111;
assign micromatrizz[70][120] = 9'b111111111;
assign micromatrizz[70][121] = 9'b111111111;
assign micromatrizz[70][122] = 9'b111111111;
assign micromatrizz[70][123] = 9'b111111111;
assign micromatrizz[70][124] = 9'b111111111;
assign micromatrizz[70][125] = 9'b111111111;
assign micromatrizz[70][126] = 9'b111111111;
assign micromatrizz[70][127] = 9'b111111111;
assign micromatrizz[70][128] = 9'b111111111;
assign micromatrizz[70][129] = 9'b111111111;
assign micromatrizz[70][130] = 9'b111111111;
assign micromatrizz[70][131] = 9'b111111111;
assign micromatrizz[70][132] = 9'b111111111;
assign micromatrizz[70][133] = 9'b111111111;
assign micromatrizz[70][134] = 9'b111111111;
assign micromatrizz[70][135] = 9'b111111111;
assign micromatrizz[70][136] = 9'b111111111;
assign micromatrizz[70][137] = 9'b111111111;
assign micromatrizz[70][138] = 9'b111111111;
assign micromatrizz[70][139] = 9'b111111111;
assign micromatrizz[70][140] = 9'b111111111;
assign micromatrizz[70][141] = 9'b111111111;
assign micromatrizz[70][142] = 9'b111111111;
assign micromatrizz[70][143] = 9'b111111111;
assign micromatrizz[70][144] = 9'b111111111;
assign micromatrizz[70][145] = 9'b111111111;
assign micromatrizz[70][146] = 9'b111111111;
assign micromatrizz[70][147] = 9'b111111111;
assign micromatrizz[70][148] = 9'b111111111;
assign micromatrizz[70][149] = 9'b111111111;
assign micromatrizz[70][150] = 9'b111111111;
assign micromatrizz[70][151] = 9'b111111111;
assign micromatrizz[70][152] = 9'b111111111;
assign micromatrizz[70][153] = 9'b111111111;
assign micromatrizz[70][154] = 9'b111111111;
assign micromatrizz[70][155] = 9'b111111111;
assign micromatrizz[70][156] = 9'b111111111;
assign micromatrizz[70][157] = 9'b111111111;
assign micromatrizz[70][158] = 9'b111111111;
assign micromatrizz[70][159] = 9'b111111111;
assign micromatrizz[70][160] = 9'b111111111;
assign micromatrizz[70][161] = 9'b111111111;
assign micromatrizz[70][162] = 9'b111111111;
assign micromatrizz[70][163] = 9'b111111111;
assign micromatrizz[70][164] = 9'b111111111;
assign micromatrizz[70][165] = 9'b111111111;
assign micromatrizz[70][166] = 9'b111111111;
assign micromatrizz[70][167] = 9'b111111111;
assign micromatrizz[70][168] = 9'b111111111;
assign micromatrizz[70][169] = 9'b111111111;
assign micromatrizz[70][170] = 9'b111111111;
assign micromatrizz[70][171] = 9'b111111111;
assign micromatrizz[70][172] = 9'b111111111;
assign micromatrizz[70][173] = 9'b111111111;
assign micromatrizz[70][174] = 9'b111111111;
assign micromatrizz[70][175] = 9'b111111111;
assign micromatrizz[70][176] = 9'b111111111;
assign micromatrizz[70][177] = 9'b111111111;
assign micromatrizz[70][178] = 9'b111111111;
assign micromatrizz[70][179] = 9'b111111111;
assign micromatrizz[70][180] = 9'b111111111;
assign micromatrizz[70][181] = 9'b111111111;
assign micromatrizz[70][182] = 9'b111111111;
assign micromatrizz[70][183] = 9'b111111111;
assign micromatrizz[70][184] = 9'b111111111;
assign micromatrizz[70][185] = 9'b111111111;
assign micromatrizz[70][186] = 9'b111111111;
assign micromatrizz[70][187] = 9'b111111111;
assign micromatrizz[70][188] = 9'b111111111;
assign micromatrizz[70][189] = 9'b111111111;
assign micromatrizz[70][190] = 9'b111111111;
assign micromatrizz[70][191] = 9'b111111111;
assign micromatrizz[70][192] = 9'b111111111;
assign micromatrizz[70][193] = 9'b111111111;
assign micromatrizz[70][194] = 9'b111111111;
assign micromatrizz[70][195] = 9'b111111111;
assign micromatrizz[70][196] = 9'b111111111;
assign micromatrizz[70][197] = 9'b111111111;
assign micromatrizz[70][198] = 9'b111111111;
assign micromatrizz[70][199] = 9'b111111111;
assign micromatrizz[70][200] = 9'b111111111;
assign micromatrizz[70][201] = 9'b111111111;
assign micromatrizz[70][202] = 9'b111111111;
assign micromatrizz[70][203] = 9'b111111111;
assign micromatrizz[70][204] = 9'b111111111;
assign micromatrizz[70][205] = 9'b111111111;
assign micromatrizz[70][206] = 9'b111111111;
assign micromatrizz[70][207] = 9'b111111111;
assign micromatrizz[70][208] = 9'b111111111;
assign micromatrizz[70][209] = 9'b111111111;
assign micromatrizz[70][210] = 9'b111111111;
assign micromatrizz[70][211] = 9'b111111111;
assign micromatrizz[70][212] = 9'b111111111;
assign micromatrizz[70][213] = 9'b111111111;
assign micromatrizz[70][214] = 9'b111111111;
assign micromatrizz[70][215] = 9'b111111111;
assign micromatrizz[70][216] = 9'b111111111;
assign micromatrizz[70][217] = 9'b111111111;
assign micromatrizz[70][218] = 9'b111111111;
assign micromatrizz[70][219] = 9'b111111111;
assign micromatrizz[70][220] = 9'b111111111;
assign micromatrizz[70][221] = 9'b111111111;
assign micromatrizz[70][222] = 9'b111111111;
assign micromatrizz[70][223] = 9'b111111111;
assign micromatrizz[70][224] = 9'b111111111;
assign micromatrizz[70][225] = 9'b111111111;
assign micromatrizz[70][226] = 9'b111111111;
assign micromatrizz[70][227] = 9'b111111111;
assign micromatrizz[70][228] = 9'b111111111;
assign micromatrizz[70][229] = 9'b111111111;
assign micromatrizz[70][230] = 9'b111111111;
assign micromatrizz[70][231] = 9'b111111111;
assign micromatrizz[70][232] = 9'b111111111;
assign micromatrizz[70][233] = 9'b111111111;
assign micromatrizz[70][234] = 9'b111111111;
assign micromatrizz[70][235] = 9'b111111111;
assign micromatrizz[70][236] = 9'b111111111;
assign micromatrizz[70][237] = 9'b111111111;
assign micromatrizz[70][238] = 9'b111111111;
assign micromatrizz[70][239] = 9'b111111111;
assign micromatrizz[70][240] = 9'b111111111;
assign micromatrizz[70][241] = 9'b111111111;
assign micromatrizz[70][242] = 9'b111111111;
assign micromatrizz[70][243] = 9'b111111111;
assign micromatrizz[70][244] = 9'b111111111;
assign micromatrizz[70][245] = 9'b111111111;
assign micromatrizz[70][246] = 9'b111111111;
assign micromatrizz[70][247] = 9'b111111111;
assign micromatrizz[70][248] = 9'b111111111;
assign micromatrizz[70][249] = 9'b111111111;
assign micromatrizz[70][250] = 9'b111111111;
assign micromatrizz[70][251] = 9'b111111111;
assign micromatrizz[70][252] = 9'b111111111;
assign micromatrizz[70][253] = 9'b111111111;
assign micromatrizz[70][254] = 9'b111111111;
assign micromatrizz[70][255] = 9'b111111111;
assign micromatrizz[70][256] = 9'b111111111;
assign micromatrizz[70][257] = 9'b111111111;
assign micromatrizz[70][258] = 9'b111111111;
assign micromatrizz[70][259] = 9'b111111111;
assign micromatrizz[70][260] = 9'b111111111;
assign micromatrizz[70][261] = 9'b111111111;
assign micromatrizz[70][262] = 9'b111111111;
assign micromatrizz[70][263] = 9'b111111111;
assign micromatrizz[70][264] = 9'b111111111;
assign micromatrizz[70][265] = 9'b111111111;
assign micromatrizz[70][266] = 9'b111111111;
assign micromatrizz[70][267] = 9'b111111111;
assign micromatrizz[70][268] = 9'b111111111;
assign micromatrizz[70][269] = 9'b111111111;
assign micromatrizz[70][270] = 9'b111111111;
assign micromatrizz[70][271] = 9'b111111111;
assign micromatrizz[70][272] = 9'b111111111;
assign micromatrizz[70][273] = 9'b111111111;
assign micromatrizz[70][274] = 9'b111111111;
assign micromatrizz[70][275] = 9'b111111111;
assign micromatrizz[70][276] = 9'b111111111;
assign micromatrizz[70][277] = 9'b111111111;
assign micromatrizz[70][278] = 9'b111111111;
assign micromatrizz[70][279] = 9'b111111111;
assign micromatrizz[70][280] = 9'b111111111;
assign micromatrizz[70][281] = 9'b111111111;
assign micromatrizz[70][282] = 9'b111111111;
assign micromatrizz[70][283] = 9'b111111111;
assign micromatrizz[70][284] = 9'b111111111;
assign micromatrizz[70][285] = 9'b111111111;
assign micromatrizz[70][286] = 9'b111111111;
assign micromatrizz[70][287] = 9'b111111111;
assign micromatrizz[70][288] = 9'b111111111;
assign micromatrizz[70][289] = 9'b111111111;
assign micromatrizz[70][290] = 9'b111111111;
assign micromatrizz[70][291] = 9'b111111111;
assign micromatrizz[70][292] = 9'b111111111;
assign micromatrizz[70][293] = 9'b111111111;
assign micromatrizz[70][294] = 9'b111111111;
assign micromatrizz[70][295] = 9'b111111111;
assign micromatrizz[70][296] = 9'b111111111;
assign micromatrizz[70][297] = 9'b111111111;
assign micromatrizz[70][298] = 9'b111111111;
assign micromatrizz[70][299] = 9'b111111111;
assign micromatrizz[70][300] = 9'b111111111;
assign micromatrizz[70][301] = 9'b111111111;
assign micromatrizz[70][302] = 9'b111111111;
assign micromatrizz[70][303] = 9'b111111111;
assign micromatrizz[70][304] = 9'b111111111;
assign micromatrizz[70][305] = 9'b111111111;
assign micromatrizz[70][306] = 9'b111111111;
assign micromatrizz[70][307] = 9'b111111111;
assign micromatrizz[70][308] = 9'b111111111;
assign micromatrizz[70][309] = 9'b111111111;
assign micromatrizz[70][310] = 9'b111111111;
assign micromatrizz[70][311] = 9'b111111111;
assign micromatrizz[70][312] = 9'b111111111;
assign micromatrizz[70][313] = 9'b111111111;
assign micromatrizz[70][314] = 9'b111111111;
assign micromatrizz[70][315] = 9'b111111111;
assign micromatrizz[70][316] = 9'b111111111;
assign micromatrizz[70][317] = 9'b111111111;
assign micromatrizz[70][318] = 9'b111111111;
assign micromatrizz[70][319] = 9'b111111111;
assign micromatrizz[70][320] = 9'b111111111;
assign micromatrizz[70][321] = 9'b111111111;
assign micromatrizz[70][322] = 9'b111111111;
assign micromatrizz[70][323] = 9'b111111111;
assign micromatrizz[70][324] = 9'b111111111;
assign micromatrizz[70][325] = 9'b111111111;
assign micromatrizz[70][326] = 9'b111111111;
assign micromatrizz[70][327] = 9'b111111111;
assign micromatrizz[70][328] = 9'b111111111;
assign micromatrizz[70][329] = 9'b111111111;
assign micromatrizz[70][330] = 9'b111111111;
assign micromatrizz[70][331] = 9'b111111111;
assign micromatrizz[70][332] = 9'b111111111;
assign micromatrizz[70][333] = 9'b111111111;
assign micromatrizz[70][334] = 9'b111111111;
assign micromatrizz[70][335] = 9'b111111111;
assign micromatrizz[70][336] = 9'b111111111;
assign micromatrizz[70][337] = 9'b111111111;
assign micromatrizz[70][338] = 9'b111111111;
assign micromatrizz[70][339] = 9'b111111111;
assign micromatrizz[70][340] = 9'b111111111;
assign micromatrizz[70][341] = 9'b111111111;
assign micromatrizz[70][342] = 9'b111111111;
assign micromatrizz[70][343] = 9'b111111111;
assign micromatrizz[70][344] = 9'b111111111;
assign micromatrizz[70][345] = 9'b111111111;
assign micromatrizz[70][346] = 9'b111111111;
assign micromatrizz[70][347] = 9'b111111111;
assign micromatrizz[70][348] = 9'b111111111;
assign micromatrizz[70][349] = 9'b111111111;
assign micromatrizz[70][350] = 9'b111111111;
assign micromatrizz[70][351] = 9'b111111111;
assign micromatrizz[70][352] = 9'b111111111;
assign micromatrizz[70][353] = 9'b111111111;
assign micromatrizz[70][354] = 9'b111111111;
assign micromatrizz[70][355] = 9'b111111111;
assign micromatrizz[70][356] = 9'b111111111;
assign micromatrizz[70][357] = 9'b111111111;
assign micromatrizz[70][358] = 9'b111111111;
assign micromatrizz[70][359] = 9'b111111111;
assign micromatrizz[70][360] = 9'b111111111;
assign micromatrizz[70][361] = 9'b111111111;
assign micromatrizz[70][362] = 9'b111111111;
assign micromatrizz[70][363] = 9'b111111111;
assign micromatrizz[70][364] = 9'b111111111;
assign micromatrizz[70][365] = 9'b111111111;
assign micromatrizz[70][366] = 9'b111111111;
assign micromatrizz[70][367] = 9'b111111111;
assign micromatrizz[70][368] = 9'b111111111;
assign micromatrizz[70][369] = 9'b111111111;
assign micromatrizz[70][370] = 9'b111111111;
assign micromatrizz[70][371] = 9'b111111111;
assign micromatrizz[70][372] = 9'b111111111;
assign micromatrizz[70][373] = 9'b111111111;
assign micromatrizz[70][374] = 9'b111111111;
assign micromatrizz[70][375] = 9'b111111111;
assign micromatrizz[70][376] = 9'b111111111;
assign micromatrizz[70][377] = 9'b111111111;
assign micromatrizz[70][378] = 9'b111111111;
assign micromatrizz[70][379] = 9'b111111111;
assign micromatrizz[70][380] = 9'b111111111;
assign micromatrizz[70][381] = 9'b111111111;
assign micromatrizz[70][382] = 9'b111111111;
assign micromatrizz[70][383] = 9'b111111111;
assign micromatrizz[70][384] = 9'b111111111;
assign micromatrizz[70][385] = 9'b111111111;
assign micromatrizz[70][386] = 9'b111111111;
assign micromatrizz[70][387] = 9'b111111111;
assign micromatrizz[70][388] = 9'b111111111;
assign micromatrizz[70][389] = 9'b111111111;
assign micromatrizz[70][390] = 9'b111111111;
assign micromatrizz[70][391] = 9'b111111111;
assign micromatrizz[70][392] = 9'b111111111;
assign micromatrizz[70][393] = 9'b111111111;
assign micromatrizz[70][394] = 9'b111111111;
assign micromatrizz[70][395] = 9'b111111111;
assign micromatrizz[70][396] = 9'b111111111;
assign micromatrizz[70][397] = 9'b111111111;
assign micromatrizz[70][398] = 9'b111111111;
assign micromatrizz[70][399] = 9'b111111111;
assign micromatrizz[70][400] = 9'b111111111;
assign micromatrizz[70][401] = 9'b111111111;
assign micromatrizz[70][402] = 9'b111111111;
assign micromatrizz[70][403] = 9'b111111111;
assign micromatrizz[70][404] = 9'b111111111;
assign micromatrizz[70][405] = 9'b111111111;
assign micromatrizz[70][406] = 9'b111111111;
assign micromatrizz[70][407] = 9'b111111111;
assign micromatrizz[70][408] = 9'b111111111;
assign micromatrizz[70][409] = 9'b111111111;
assign micromatrizz[70][410] = 9'b111111111;
assign micromatrizz[70][411] = 9'b111111111;
assign micromatrizz[70][412] = 9'b111111111;
assign micromatrizz[70][413] = 9'b111111111;
assign micromatrizz[70][414] = 9'b111111111;
assign micromatrizz[70][415] = 9'b111111111;
assign micromatrizz[70][416] = 9'b111111111;
assign micromatrizz[70][417] = 9'b111111111;
assign micromatrizz[70][418] = 9'b111111111;
assign micromatrizz[70][419] = 9'b111111111;
assign micromatrizz[70][420] = 9'b111111111;
assign micromatrizz[70][421] = 9'b111111111;
assign micromatrizz[70][422] = 9'b111111111;
assign micromatrizz[70][423] = 9'b111111111;
assign micromatrizz[70][424] = 9'b111111111;
assign micromatrizz[70][425] = 9'b111111111;
assign micromatrizz[70][426] = 9'b111111111;
assign micromatrizz[70][427] = 9'b111111111;
assign micromatrizz[70][428] = 9'b111111111;
assign micromatrizz[70][429] = 9'b111111111;
assign micromatrizz[70][430] = 9'b111111111;
assign micromatrizz[70][431] = 9'b111111111;
assign micromatrizz[70][432] = 9'b111111111;
assign micromatrizz[70][433] = 9'b111111111;
assign micromatrizz[70][434] = 9'b111111111;
assign micromatrizz[70][435] = 9'b111111111;
assign micromatrizz[70][436] = 9'b111111111;
assign micromatrizz[70][437] = 9'b111111111;
assign micromatrizz[70][438] = 9'b111111111;
assign micromatrizz[70][439] = 9'b111111111;
assign micromatrizz[70][440] = 9'b111111111;
assign micromatrizz[70][441] = 9'b111111111;
assign micromatrizz[70][442] = 9'b111111111;
assign micromatrizz[70][443] = 9'b111111111;
assign micromatrizz[70][444] = 9'b111111111;
assign micromatrizz[70][445] = 9'b111111111;
assign micromatrizz[70][446] = 9'b111111111;
assign micromatrizz[70][447] = 9'b111111111;
assign micromatrizz[70][448] = 9'b111111111;
assign micromatrizz[70][449] = 9'b111111111;
assign micromatrizz[70][450] = 9'b111111111;
assign micromatrizz[70][451] = 9'b111111111;
assign micromatrizz[70][452] = 9'b111111111;
assign micromatrizz[70][453] = 9'b111111111;
assign micromatrizz[70][454] = 9'b111111111;
assign micromatrizz[70][455] = 9'b111111111;
assign micromatrizz[70][456] = 9'b111111111;
assign micromatrizz[70][457] = 9'b111111111;
assign micromatrizz[70][458] = 9'b111111111;
assign micromatrizz[70][459] = 9'b111111111;
assign micromatrizz[70][460] = 9'b111111111;
assign micromatrizz[70][461] = 9'b111111111;
assign micromatrizz[70][462] = 9'b111111111;
assign micromatrizz[70][463] = 9'b111111111;
assign micromatrizz[70][464] = 9'b111111111;
assign micromatrizz[70][465] = 9'b111111111;
assign micromatrizz[70][466] = 9'b111111111;
assign micromatrizz[70][467] = 9'b111111111;
assign micromatrizz[70][468] = 9'b111111111;
assign micromatrizz[70][469] = 9'b111111111;
assign micromatrizz[70][470] = 9'b111111111;
assign micromatrizz[70][471] = 9'b111111111;
assign micromatrizz[70][472] = 9'b111111111;
assign micromatrizz[70][473] = 9'b111111111;
assign micromatrizz[70][474] = 9'b111111111;
assign micromatrizz[70][475] = 9'b111111111;
assign micromatrizz[70][476] = 9'b111111111;
assign micromatrizz[70][477] = 9'b111111111;
assign micromatrizz[70][478] = 9'b111111111;
assign micromatrizz[70][479] = 9'b111111111;
assign micromatrizz[70][480] = 9'b111111111;
assign micromatrizz[70][481] = 9'b111111111;
assign micromatrizz[70][482] = 9'b111111111;
assign micromatrizz[70][483] = 9'b111111111;
assign micromatrizz[70][484] = 9'b111111111;
assign micromatrizz[70][485] = 9'b111111111;
assign micromatrizz[70][486] = 9'b111111111;
assign micromatrizz[70][487] = 9'b111111111;
assign micromatrizz[70][488] = 9'b111111111;
assign micromatrizz[70][489] = 9'b111111111;
assign micromatrizz[70][490] = 9'b111111111;
assign micromatrizz[70][491] = 9'b111111111;
assign micromatrizz[70][492] = 9'b111111111;
assign micromatrizz[70][493] = 9'b111111111;
assign micromatrizz[70][494] = 9'b111111111;
assign micromatrizz[70][495] = 9'b111111111;
assign micromatrizz[70][496] = 9'b111111111;
assign micromatrizz[70][497] = 9'b111111111;
assign micromatrizz[70][498] = 9'b111111111;
assign micromatrizz[70][499] = 9'b111111111;
assign micromatrizz[70][500] = 9'b111111111;
assign micromatrizz[70][501] = 9'b111111111;
assign micromatrizz[70][502] = 9'b111111111;
assign micromatrizz[70][503] = 9'b111111111;
assign micromatrizz[70][504] = 9'b111111111;
assign micromatrizz[70][505] = 9'b111111111;
assign micromatrizz[70][506] = 9'b111111111;
assign micromatrizz[70][507] = 9'b111111111;
assign micromatrizz[70][508] = 9'b111111111;
assign micromatrizz[70][509] = 9'b111111111;
assign micromatrizz[70][510] = 9'b111111111;
assign micromatrizz[70][511] = 9'b111111111;
assign micromatrizz[70][512] = 9'b111111111;
assign micromatrizz[70][513] = 9'b111111111;
assign micromatrizz[70][514] = 9'b111111111;
assign micromatrizz[70][515] = 9'b111111111;
assign micromatrizz[70][516] = 9'b111111111;
assign micromatrizz[70][517] = 9'b111111111;
assign micromatrizz[70][518] = 9'b111111111;
assign micromatrizz[70][519] = 9'b111111111;
assign micromatrizz[70][520] = 9'b111111111;
assign micromatrizz[70][521] = 9'b111111111;
assign micromatrizz[70][522] = 9'b111111111;
assign micromatrizz[70][523] = 9'b111111111;
assign micromatrizz[70][524] = 9'b111111111;
assign micromatrizz[70][525] = 9'b111111111;
assign micromatrizz[70][526] = 9'b111111111;
assign micromatrizz[70][527] = 9'b111111111;
assign micromatrizz[70][528] = 9'b111111111;
assign micromatrizz[70][529] = 9'b111111111;
assign micromatrizz[70][530] = 9'b111111111;
assign micromatrizz[70][531] = 9'b111111111;
assign micromatrizz[70][532] = 9'b111111111;
assign micromatrizz[70][533] = 9'b111111111;
assign micromatrizz[70][534] = 9'b111111111;
assign micromatrizz[70][535] = 9'b111111111;
assign micromatrizz[70][536] = 9'b111111111;
assign micromatrizz[70][537] = 9'b111111111;
assign micromatrizz[70][538] = 9'b111111111;
assign micromatrizz[70][539] = 9'b111111111;
assign micromatrizz[70][540] = 9'b111111111;
assign micromatrizz[70][541] = 9'b111111111;
assign micromatrizz[70][542] = 9'b111111111;
assign micromatrizz[70][543] = 9'b111111111;
assign micromatrizz[70][544] = 9'b111111111;
assign micromatrizz[70][545] = 9'b111111111;
assign micromatrizz[70][546] = 9'b111111111;
assign micromatrizz[70][547] = 9'b111111111;
assign micromatrizz[70][548] = 9'b111111111;
assign micromatrizz[70][549] = 9'b111111111;
assign micromatrizz[70][550] = 9'b111111111;
assign micromatrizz[70][551] = 9'b111111111;
assign micromatrizz[70][552] = 9'b111111111;
assign micromatrizz[70][553] = 9'b111111111;
assign micromatrizz[70][554] = 9'b111111111;
assign micromatrizz[70][555] = 9'b111111111;
assign micromatrizz[70][556] = 9'b111111111;
assign micromatrizz[70][557] = 9'b111111111;
assign micromatrizz[70][558] = 9'b111111111;
assign micromatrizz[70][559] = 9'b111111111;
assign micromatrizz[70][560] = 9'b111111111;
assign micromatrizz[70][561] = 9'b111111111;
assign micromatrizz[70][562] = 9'b111111111;
assign micromatrizz[70][563] = 9'b111111111;
assign micromatrizz[70][564] = 9'b111111111;
assign micromatrizz[70][565] = 9'b111111111;
assign micromatrizz[70][566] = 9'b111111111;
assign micromatrizz[70][567] = 9'b111111111;
assign micromatrizz[70][568] = 9'b111111111;
assign micromatrizz[70][569] = 9'b111111111;
assign micromatrizz[70][570] = 9'b111111111;
assign micromatrizz[70][571] = 9'b111111111;
assign micromatrizz[70][572] = 9'b111111111;
assign micromatrizz[70][573] = 9'b111111111;
assign micromatrizz[70][574] = 9'b111111111;
assign micromatrizz[70][575] = 9'b111111111;
assign micromatrizz[70][576] = 9'b111111111;
assign micromatrizz[70][577] = 9'b111111111;
assign micromatrizz[70][578] = 9'b111111111;
assign micromatrizz[70][579] = 9'b111111111;
assign micromatrizz[70][580] = 9'b111111111;
assign micromatrizz[70][581] = 9'b111111111;
assign micromatrizz[70][582] = 9'b111111111;
assign micromatrizz[70][583] = 9'b111111111;
assign micromatrizz[70][584] = 9'b111111111;
assign micromatrizz[70][585] = 9'b111111111;
assign micromatrizz[70][586] = 9'b111111111;
assign micromatrizz[70][587] = 9'b111111111;
assign micromatrizz[70][588] = 9'b111111111;
assign micromatrizz[70][589] = 9'b111111111;
assign micromatrizz[70][590] = 9'b111111111;
assign micromatrizz[70][591] = 9'b111111111;
assign micromatrizz[70][592] = 9'b111111111;
assign micromatrizz[70][593] = 9'b111111111;
assign micromatrizz[70][594] = 9'b111111111;
assign micromatrizz[70][595] = 9'b111111111;
assign micromatrizz[70][596] = 9'b111111111;
assign micromatrizz[70][597] = 9'b111111111;
assign micromatrizz[70][598] = 9'b111111111;
assign micromatrizz[70][599] = 9'b111111111;
assign micromatrizz[70][600] = 9'b111111111;
assign micromatrizz[70][601] = 9'b111111111;
assign micromatrizz[70][602] = 9'b111111111;
assign micromatrizz[70][603] = 9'b111111111;
assign micromatrizz[70][604] = 9'b111111111;
assign micromatrizz[70][605] = 9'b111111111;
assign micromatrizz[70][606] = 9'b111111111;
assign micromatrizz[70][607] = 9'b111111111;
assign micromatrizz[70][608] = 9'b111111111;
assign micromatrizz[70][609] = 9'b111111111;
assign micromatrizz[70][610] = 9'b111111111;
assign micromatrizz[70][611] = 9'b111111111;
assign micromatrizz[70][612] = 9'b111111111;
assign micromatrizz[70][613] = 9'b111111111;
assign micromatrizz[70][614] = 9'b111111111;
assign micromatrizz[70][615] = 9'b111111111;
assign micromatrizz[70][616] = 9'b111111111;
assign micromatrizz[70][617] = 9'b111111111;
assign micromatrizz[70][618] = 9'b111111111;
assign micromatrizz[70][619] = 9'b111111111;
assign micromatrizz[70][620] = 9'b111111111;
assign micromatrizz[70][621] = 9'b111111111;
assign micromatrizz[70][622] = 9'b111111111;
assign micromatrizz[70][623] = 9'b111111111;
assign micromatrizz[70][624] = 9'b111111111;
assign micromatrizz[70][625] = 9'b111111111;
assign micromatrizz[70][626] = 9'b111111111;
assign micromatrizz[70][627] = 9'b111111111;
assign micromatrizz[70][628] = 9'b111111111;
assign micromatrizz[70][629] = 9'b111111111;
assign micromatrizz[70][630] = 9'b111111111;
assign micromatrizz[70][631] = 9'b111111111;
assign micromatrizz[70][632] = 9'b111111111;
assign micromatrizz[70][633] = 9'b111111111;
assign micromatrizz[70][634] = 9'b111111111;
assign micromatrizz[70][635] = 9'b111111111;
assign micromatrizz[70][636] = 9'b111111111;
assign micromatrizz[70][637] = 9'b111111111;
assign micromatrizz[70][638] = 9'b111111111;
assign micromatrizz[70][639] = 9'b111111111;
assign micromatrizz[71][0] = 9'b111111111;
assign micromatrizz[71][1] = 9'b111111111;
assign micromatrizz[71][2] = 9'b111111111;
assign micromatrizz[71][3] = 9'b111111111;
assign micromatrizz[71][4] = 9'b111111111;
assign micromatrizz[71][5] = 9'b111111111;
assign micromatrizz[71][6] = 9'b111111111;
assign micromatrizz[71][7] = 9'b111111111;
assign micromatrizz[71][8] = 9'b111111111;
assign micromatrizz[71][9] = 9'b111111111;
assign micromatrizz[71][10] = 9'b111111111;
assign micromatrizz[71][11] = 9'b111111111;
assign micromatrizz[71][12] = 9'b111111111;
assign micromatrizz[71][13] = 9'b111111111;
assign micromatrizz[71][14] = 9'b111111111;
assign micromatrizz[71][15] = 9'b111111111;
assign micromatrizz[71][16] = 9'b111111111;
assign micromatrizz[71][17] = 9'b111111111;
assign micromatrizz[71][18] = 9'b111111111;
assign micromatrizz[71][19] = 9'b111111111;
assign micromatrizz[71][20] = 9'b111111111;
assign micromatrizz[71][21] = 9'b111111111;
assign micromatrizz[71][22] = 9'b111111111;
assign micromatrizz[71][23] = 9'b111111111;
assign micromatrizz[71][24] = 9'b111111111;
assign micromatrizz[71][25] = 9'b111111111;
assign micromatrizz[71][26] = 9'b111111111;
assign micromatrizz[71][27] = 9'b111111111;
assign micromatrizz[71][28] = 9'b111111111;
assign micromatrizz[71][29] = 9'b111111111;
assign micromatrizz[71][30] = 9'b111111111;
assign micromatrizz[71][31] = 9'b111111111;
assign micromatrizz[71][32] = 9'b111111111;
assign micromatrizz[71][33] = 9'b111111111;
assign micromatrizz[71][34] = 9'b111111111;
assign micromatrizz[71][35] = 9'b111111111;
assign micromatrizz[71][36] = 9'b111111111;
assign micromatrizz[71][37] = 9'b111111111;
assign micromatrizz[71][38] = 9'b111111111;
assign micromatrizz[71][39] = 9'b111111111;
assign micromatrizz[71][40] = 9'b111111111;
assign micromatrizz[71][41] = 9'b111111111;
assign micromatrizz[71][42] = 9'b111111111;
assign micromatrizz[71][43] = 9'b111111111;
assign micromatrizz[71][44] = 9'b111111111;
assign micromatrizz[71][45] = 9'b111111111;
assign micromatrizz[71][46] = 9'b111111111;
assign micromatrizz[71][47] = 9'b111111111;
assign micromatrizz[71][48] = 9'b111111111;
assign micromatrizz[71][49] = 9'b111111111;
assign micromatrizz[71][50] = 9'b111111111;
assign micromatrizz[71][51] = 9'b111111111;
assign micromatrizz[71][52] = 9'b111111111;
assign micromatrizz[71][53] = 9'b111111111;
assign micromatrizz[71][54] = 9'b111111111;
assign micromatrizz[71][55] = 9'b111111111;
assign micromatrizz[71][56] = 9'b111111111;
assign micromatrizz[71][57] = 9'b111111111;
assign micromatrizz[71][58] = 9'b111111111;
assign micromatrizz[71][59] = 9'b111111111;
assign micromatrizz[71][60] = 9'b111111111;
assign micromatrizz[71][61] = 9'b111111111;
assign micromatrizz[71][62] = 9'b111111111;
assign micromatrizz[71][63] = 9'b111111111;
assign micromatrizz[71][64] = 9'b111111111;
assign micromatrizz[71][65] = 9'b111111111;
assign micromatrizz[71][66] = 9'b111111111;
assign micromatrizz[71][67] = 9'b111111111;
assign micromatrizz[71][68] = 9'b111111111;
assign micromatrizz[71][69] = 9'b111111111;
assign micromatrizz[71][70] = 9'b111111111;
assign micromatrizz[71][71] = 9'b111111111;
assign micromatrizz[71][72] = 9'b111111111;
assign micromatrizz[71][73] = 9'b111111111;
assign micromatrizz[71][74] = 9'b111111111;
assign micromatrizz[71][75] = 9'b111111111;
assign micromatrizz[71][76] = 9'b111111111;
assign micromatrizz[71][77] = 9'b111111111;
assign micromatrizz[71][78] = 9'b111111111;
assign micromatrizz[71][79] = 9'b111111111;
assign micromatrizz[71][80] = 9'b111111111;
assign micromatrizz[71][81] = 9'b111111111;
assign micromatrizz[71][82] = 9'b111111111;
assign micromatrizz[71][83] = 9'b111111111;
assign micromatrizz[71][84] = 9'b111111111;
assign micromatrizz[71][85] = 9'b111111111;
assign micromatrizz[71][86] = 9'b111111111;
assign micromatrizz[71][87] = 9'b111111111;
assign micromatrizz[71][88] = 9'b111111111;
assign micromatrizz[71][89] = 9'b111111111;
assign micromatrizz[71][90] = 9'b111111111;
assign micromatrizz[71][91] = 9'b111111111;
assign micromatrizz[71][92] = 9'b111111111;
assign micromatrizz[71][93] = 9'b111111111;
assign micromatrizz[71][94] = 9'b111111111;
assign micromatrizz[71][95] = 9'b111111111;
assign micromatrizz[71][96] = 9'b111111111;
assign micromatrizz[71][97] = 9'b111111111;
assign micromatrizz[71][98] = 9'b111111111;
assign micromatrizz[71][99] = 9'b111111111;
assign micromatrizz[71][100] = 9'b111111111;
assign micromatrizz[71][101] = 9'b111111111;
assign micromatrizz[71][102] = 9'b111111111;
assign micromatrizz[71][103] = 9'b111111111;
assign micromatrizz[71][104] = 9'b111111111;
assign micromatrizz[71][105] = 9'b111111111;
assign micromatrizz[71][106] = 9'b111111111;
assign micromatrizz[71][107] = 9'b111111111;
assign micromatrizz[71][108] = 9'b111111111;
assign micromatrizz[71][109] = 9'b111111111;
assign micromatrizz[71][110] = 9'b111111111;
assign micromatrizz[71][111] = 9'b111111111;
assign micromatrizz[71][112] = 9'b111111111;
assign micromatrizz[71][113] = 9'b111111111;
assign micromatrizz[71][114] = 9'b111111111;
assign micromatrizz[71][115] = 9'b111111111;
assign micromatrizz[71][116] = 9'b111111111;
assign micromatrizz[71][117] = 9'b111111111;
assign micromatrizz[71][118] = 9'b111111111;
assign micromatrizz[71][119] = 9'b111111111;
assign micromatrizz[71][120] = 9'b111111111;
assign micromatrizz[71][121] = 9'b111111111;
assign micromatrizz[71][122] = 9'b111111111;
assign micromatrizz[71][123] = 9'b111111111;
assign micromatrizz[71][124] = 9'b111111111;
assign micromatrizz[71][125] = 9'b111111111;
assign micromatrizz[71][126] = 9'b111111111;
assign micromatrizz[71][127] = 9'b111111111;
assign micromatrizz[71][128] = 9'b111111111;
assign micromatrizz[71][129] = 9'b111111111;
assign micromatrizz[71][130] = 9'b111111111;
assign micromatrizz[71][131] = 9'b111111111;
assign micromatrizz[71][132] = 9'b111111111;
assign micromatrizz[71][133] = 9'b111111111;
assign micromatrizz[71][134] = 9'b111111111;
assign micromatrizz[71][135] = 9'b111111111;
assign micromatrizz[71][136] = 9'b111111111;
assign micromatrizz[71][137] = 9'b111111111;
assign micromatrizz[71][138] = 9'b111111111;
assign micromatrizz[71][139] = 9'b111111111;
assign micromatrizz[71][140] = 9'b111111111;
assign micromatrizz[71][141] = 9'b111111111;
assign micromatrizz[71][142] = 9'b111111111;
assign micromatrizz[71][143] = 9'b111111111;
assign micromatrizz[71][144] = 9'b111111111;
assign micromatrizz[71][145] = 9'b111111111;
assign micromatrizz[71][146] = 9'b111111111;
assign micromatrizz[71][147] = 9'b111111111;
assign micromatrizz[71][148] = 9'b111111111;
assign micromatrizz[71][149] = 9'b111111111;
assign micromatrizz[71][150] = 9'b111111111;
assign micromatrizz[71][151] = 9'b111111111;
assign micromatrizz[71][152] = 9'b111111111;
assign micromatrizz[71][153] = 9'b111111111;
assign micromatrizz[71][154] = 9'b111111111;
assign micromatrizz[71][155] = 9'b111111111;
assign micromatrizz[71][156] = 9'b111111111;
assign micromatrizz[71][157] = 9'b111111111;
assign micromatrizz[71][158] = 9'b111111111;
assign micromatrizz[71][159] = 9'b111111111;
assign micromatrizz[71][160] = 9'b111111111;
assign micromatrizz[71][161] = 9'b111111111;
assign micromatrizz[71][162] = 9'b111111111;
assign micromatrizz[71][163] = 9'b111111111;
assign micromatrizz[71][164] = 9'b111111111;
assign micromatrizz[71][165] = 9'b111111111;
assign micromatrizz[71][166] = 9'b111111111;
assign micromatrizz[71][167] = 9'b111111111;
assign micromatrizz[71][168] = 9'b111111111;
assign micromatrizz[71][169] = 9'b111111111;
assign micromatrizz[71][170] = 9'b111111111;
assign micromatrizz[71][171] = 9'b111111111;
assign micromatrizz[71][172] = 9'b111111111;
assign micromatrizz[71][173] = 9'b111111111;
assign micromatrizz[71][174] = 9'b111111111;
assign micromatrizz[71][175] = 9'b111111111;
assign micromatrizz[71][176] = 9'b111111111;
assign micromatrizz[71][177] = 9'b111111111;
assign micromatrizz[71][178] = 9'b111111111;
assign micromatrizz[71][179] = 9'b111111111;
assign micromatrizz[71][180] = 9'b111111111;
assign micromatrizz[71][181] = 9'b111111111;
assign micromatrizz[71][182] = 9'b111111111;
assign micromatrizz[71][183] = 9'b111111111;
assign micromatrizz[71][184] = 9'b111111111;
assign micromatrizz[71][185] = 9'b111111111;
assign micromatrizz[71][186] = 9'b111111111;
assign micromatrizz[71][187] = 9'b111111111;
assign micromatrizz[71][188] = 9'b111111111;
assign micromatrizz[71][189] = 9'b111111111;
assign micromatrizz[71][190] = 9'b111111111;
assign micromatrizz[71][191] = 9'b111111111;
assign micromatrizz[71][192] = 9'b111111111;
assign micromatrizz[71][193] = 9'b111111111;
assign micromatrizz[71][194] = 9'b111111111;
assign micromatrizz[71][195] = 9'b111111111;
assign micromatrizz[71][196] = 9'b111111111;
assign micromatrizz[71][197] = 9'b111111111;
assign micromatrizz[71][198] = 9'b111111111;
assign micromatrizz[71][199] = 9'b111111111;
assign micromatrizz[71][200] = 9'b111111111;
assign micromatrizz[71][201] = 9'b111111111;
assign micromatrizz[71][202] = 9'b111111111;
assign micromatrizz[71][203] = 9'b111111111;
assign micromatrizz[71][204] = 9'b111111111;
assign micromatrizz[71][205] = 9'b111111111;
assign micromatrizz[71][206] = 9'b111111111;
assign micromatrizz[71][207] = 9'b111111111;
assign micromatrizz[71][208] = 9'b111111111;
assign micromatrizz[71][209] = 9'b111111111;
assign micromatrizz[71][210] = 9'b111111111;
assign micromatrizz[71][211] = 9'b111111111;
assign micromatrizz[71][212] = 9'b111111111;
assign micromatrizz[71][213] = 9'b111111111;
assign micromatrizz[71][214] = 9'b111111111;
assign micromatrizz[71][215] = 9'b111111111;
assign micromatrizz[71][216] = 9'b111111111;
assign micromatrizz[71][217] = 9'b111111111;
assign micromatrizz[71][218] = 9'b111111111;
assign micromatrizz[71][219] = 9'b111111111;
assign micromatrizz[71][220] = 9'b111111111;
assign micromatrizz[71][221] = 9'b111111111;
assign micromatrizz[71][222] = 9'b111111111;
assign micromatrizz[71][223] = 9'b111111111;
assign micromatrizz[71][224] = 9'b111111111;
assign micromatrizz[71][225] = 9'b111111111;
assign micromatrizz[71][226] = 9'b111111111;
assign micromatrizz[71][227] = 9'b111111111;
assign micromatrizz[71][228] = 9'b111111111;
assign micromatrizz[71][229] = 9'b111111111;
assign micromatrizz[71][230] = 9'b111111111;
assign micromatrizz[71][231] = 9'b111111111;
assign micromatrizz[71][232] = 9'b111111111;
assign micromatrizz[71][233] = 9'b111111111;
assign micromatrizz[71][234] = 9'b111111111;
assign micromatrizz[71][235] = 9'b111111111;
assign micromatrizz[71][236] = 9'b111111111;
assign micromatrizz[71][237] = 9'b111111111;
assign micromatrizz[71][238] = 9'b111111111;
assign micromatrizz[71][239] = 9'b111111111;
assign micromatrizz[71][240] = 9'b111111111;
assign micromatrizz[71][241] = 9'b111111111;
assign micromatrizz[71][242] = 9'b111111111;
assign micromatrizz[71][243] = 9'b111111111;
assign micromatrizz[71][244] = 9'b111111111;
assign micromatrizz[71][245] = 9'b111111111;
assign micromatrizz[71][246] = 9'b111111111;
assign micromatrizz[71][247] = 9'b111111111;
assign micromatrizz[71][248] = 9'b111111111;
assign micromatrizz[71][249] = 9'b111111111;
assign micromatrizz[71][250] = 9'b111111111;
assign micromatrizz[71][251] = 9'b111111111;
assign micromatrizz[71][252] = 9'b111111111;
assign micromatrizz[71][253] = 9'b111111111;
assign micromatrizz[71][254] = 9'b111111111;
assign micromatrizz[71][255] = 9'b111111111;
assign micromatrizz[71][256] = 9'b111111111;
assign micromatrizz[71][257] = 9'b111111111;
assign micromatrizz[71][258] = 9'b111111111;
assign micromatrizz[71][259] = 9'b111111111;
assign micromatrizz[71][260] = 9'b111111111;
assign micromatrizz[71][261] = 9'b111111111;
assign micromatrizz[71][262] = 9'b111111111;
assign micromatrizz[71][263] = 9'b111111111;
assign micromatrizz[71][264] = 9'b111111111;
assign micromatrizz[71][265] = 9'b111111111;
assign micromatrizz[71][266] = 9'b111111111;
assign micromatrizz[71][267] = 9'b111111111;
assign micromatrizz[71][268] = 9'b111111111;
assign micromatrizz[71][269] = 9'b111111111;
assign micromatrizz[71][270] = 9'b111111111;
assign micromatrizz[71][271] = 9'b111111111;
assign micromatrizz[71][272] = 9'b111111111;
assign micromatrizz[71][273] = 9'b111111111;
assign micromatrizz[71][274] = 9'b111111111;
assign micromatrizz[71][275] = 9'b111111111;
assign micromatrizz[71][276] = 9'b111111111;
assign micromatrizz[71][277] = 9'b111111111;
assign micromatrizz[71][278] = 9'b111111111;
assign micromatrizz[71][279] = 9'b111111111;
assign micromatrizz[71][280] = 9'b111111111;
assign micromatrizz[71][281] = 9'b111111111;
assign micromatrizz[71][282] = 9'b111111111;
assign micromatrizz[71][283] = 9'b111111111;
assign micromatrizz[71][284] = 9'b111111111;
assign micromatrizz[71][285] = 9'b111111111;
assign micromatrizz[71][286] = 9'b111111111;
assign micromatrizz[71][287] = 9'b111111111;
assign micromatrizz[71][288] = 9'b111111111;
assign micromatrizz[71][289] = 9'b111111111;
assign micromatrizz[71][290] = 9'b111111111;
assign micromatrizz[71][291] = 9'b111111111;
assign micromatrizz[71][292] = 9'b111111111;
assign micromatrizz[71][293] = 9'b111111111;
assign micromatrizz[71][294] = 9'b111111111;
assign micromatrizz[71][295] = 9'b111111111;
assign micromatrizz[71][296] = 9'b111111111;
assign micromatrizz[71][297] = 9'b111111111;
assign micromatrizz[71][298] = 9'b111111111;
assign micromatrizz[71][299] = 9'b111111111;
assign micromatrizz[71][300] = 9'b111111111;
assign micromatrizz[71][301] = 9'b111111111;
assign micromatrizz[71][302] = 9'b111111111;
assign micromatrizz[71][303] = 9'b111111111;
assign micromatrizz[71][304] = 9'b111111111;
assign micromatrizz[71][305] = 9'b111111111;
assign micromatrizz[71][306] = 9'b111111111;
assign micromatrizz[71][307] = 9'b111111111;
assign micromatrizz[71][308] = 9'b111111111;
assign micromatrizz[71][309] = 9'b111111111;
assign micromatrizz[71][310] = 9'b111111111;
assign micromatrizz[71][311] = 9'b111111111;
assign micromatrizz[71][312] = 9'b111111111;
assign micromatrizz[71][313] = 9'b111111111;
assign micromatrizz[71][314] = 9'b111111111;
assign micromatrizz[71][315] = 9'b111111111;
assign micromatrizz[71][316] = 9'b111111111;
assign micromatrizz[71][317] = 9'b111111111;
assign micromatrizz[71][318] = 9'b111111111;
assign micromatrizz[71][319] = 9'b111111111;
assign micromatrizz[71][320] = 9'b111111111;
assign micromatrizz[71][321] = 9'b111111111;
assign micromatrizz[71][322] = 9'b111111111;
assign micromatrizz[71][323] = 9'b111111111;
assign micromatrizz[71][324] = 9'b111111111;
assign micromatrizz[71][325] = 9'b111111111;
assign micromatrizz[71][326] = 9'b111111111;
assign micromatrizz[71][327] = 9'b111111111;
assign micromatrizz[71][328] = 9'b111111111;
assign micromatrizz[71][329] = 9'b111111111;
assign micromatrizz[71][330] = 9'b111111111;
assign micromatrizz[71][331] = 9'b111111111;
assign micromatrizz[71][332] = 9'b111111111;
assign micromatrizz[71][333] = 9'b111111111;
assign micromatrizz[71][334] = 9'b111111111;
assign micromatrizz[71][335] = 9'b111111111;
assign micromatrizz[71][336] = 9'b111111111;
assign micromatrizz[71][337] = 9'b111111111;
assign micromatrizz[71][338] = 9'b111111111;
assign micromatrizz[71][339] = 9'b111111111;
assign micromatrizz[71][340] = 9'b111111111;
assign micromatrizz[71][341] = 9'b111111111;
assign micromatrizz[71][342] = 9'b111111111;
assign micromatrizz[71][343] = 9'b111111111;
assign micromatrizz[71][344] = 9'b111111111;
assign micromatrizz[71][345] = 9'b111111111;
assign micromatrizz[71][346] = 9'b111111111;
assign micromatrizz[71][347] = 9'b111111111;
assign micromatrizz[71][348] = 9'b111111111;
assign micromatrizz[71][349] = 9'b111111111;
assign micromatrizz[71][350] = 9'b111111111;
assign micromatrizz[71][351] = 9'b111111111;
assign micromatrizz[71][352] = 9'b111111111;
assign micromatrizz[71][353] = 9'b111111111;
assign micromatrizz[71][354] = 9'b111111111;
assign micromatrizz[71][355] = 9'b111111111;
assign micromatrizz[71][356] = 9'b111111111;
assign micromatrizz[71][357] = 9'b111111111;
assign micromatrizz[71][358] = 9'b111111111;
assign micromatrizz[71][359] = 9'b111111111;
assign micromatrizz[71][360] = 9'b111111111;
assign micromatrizz[71][361] = 9'b111111111;
assign micromatrizz[71][362] = 9'b111111111;
assign micromatrizz[71][363] = 9'b111111111;
assign micromatrizz[71][364] = 9'b111111111;
assign micromatrizz[71][365] = 9'b111111111;
assign micromatrizz[71][366] = 9'b111111111;
assign micromatrizz[71][367] = 9'b111111111;
assign micromatrizz[71][368] = 9'b111111111;
assign micromatrizz[71][369] = 9'b111111111;
assign micromatrizz[71][370] = 9'b111111111;
assign micromatrizz[71][371] = 9'b111111111;
assign micromatrizz[71][372] = 9'b111111111;
assign micromatrizz[71][373] = 9'b111111111;
assign micromatrizz[71][374] = 9'b111111111;
assign micromatrizz[71][375] = 9'b111111111;
assign micromatrizz[71][376] = 9'b111111111;
assign micromatrizz[71][377] = 9'b111111111;
assign micromatrizz[71][378] = 9'b111111111;
assign micromatrizz[71][379] = 9'b111111111;
assign micromatrizz[71][380] = 9'b111111111;
assign micromatrizz[71][381] = 9'b111111111;
assign micromatrizz[71][382] = 9'b111111111;
assign micromatrizz[71][383] = 9'b111111111;
assign micromatrizz[71][384] = 9'b111111111;
assign micromatrizz[71][385] = 9'b111111111;
assign micromatrizz[71][386] = 9'b111111111;
assign micromatrizz[71][387] = 9'b111111111;
assign micromatrizz[71][388] = 9'b111111111;
assign micromatrizz[71][389] = 9'b111111111;
assign micromatrizz[71][390] = 9'b111111111;
assign micromatrizz[71][391] = 9'b111111111;
assign micromatrizz[71][392] = 9'b111111111;
assign micromatrizz[71][393] = 9'b111111111;
assign micromatrizz[71][394] = 9'b111111111;
assign micromatrizz[71][395] = 9'b111111111;
assign micromatrizz[71][396] = 9'b111111111;
assign micromatrizz[71][397] = 9'b111111111;
assign micromatrizz[71][398] = 9'b111111111;
assign micromatrizz[71][399] = 9'b111111111;
assign micromatrizz[71][400] = 9'b111111111;
assign micromatrizz[71][401] = 9'b111111111;
assign micromatrizz[71][402] = 9'b111111111;
assign micromatrizz[71][403] = 9'b111111111;
assign micromatrizz[71][404] = 9'b111111111;
assign micromatrizz[71][405] = 9'b111111111;
assign micromatrizz[71][406] = 9'b111111111;
assign micromatrizz[71][407] = 9'b111111111;
assign micromatrizz[71][408] = 9'b111111111;
assign micromatrizz[71][409] = 9'b111111111;
assign micromatrizz[71][410] = 9'b111111111;
assign micromatrizz[71][411] = 9'b111111111;
assign micromatrizz[71][412] = 9'b111111111;
assign micromatrizz[71][413] = 9'b111111111;
assign micromatrizz[71][414] = 9'b111111111;
assign micromatrizz[71][415] = 9'b111111111;
assign micromatrizz[71][416] = 9'b111111111;
assign micromatrizz[71][417] = 9'b111111111;
assign micromatrizz[71][418] = 9'b111111111;
assign micromatrizz[71][419] = 9'b111111111;
assign micromatrizz[71][420] = 9'b111111111;
assign micromatrizz[71][421] = 9'b111111111;
assign micromatrizz[71][422] = 9'b111111111;
assign micromatrizz[71][423] = 9'b111111111;
assign micromatrizz[71][424] = 9'b111111111;
assign micromatrizz[71][425] = 9'b111111111;
assign micromatrizz[71][426] = 9'b111111111;
assign micromatrizz[71][427] = 9'b111111111;
assign micromatrizz[71][428] = 9'b111111111;
assign micromatrizz[71][429] = 9'b111111111;
assign micromatrizz[71][430] = 9'b111111111;
assign micromatrizz[71][431] = 9'b111111111;
assign micromatrizz[71][432] = 9'b111111111;
assign micromatrizz[71][433] = 9'b111111111;
assign micromatrizz[71][434] = 9'b111111111;
assign micromatrizz[71][435] = 9'b111111111;
assign micromatrizz[71][436] = 9'b111111111;
assign micromatrizz[71][437] = 9'b111111111;
assign micromatrizz[71][438] = 9'b111111111;
assign micromatrizz[71][439] = 9'b111111111;
assign micromatrizz[71][440] = 9'b111111111;
assign micromatrizz[71][441] = 9'b111111111;
assign micromatrizz[71][442] = 9'b111111111;
assign micromatrizz[71][443] = 9'b111111111;
assign micromatrizz[71][444] = 9'b111111111;
assign micromatrizz[71][445] = 9'b111111111;
assign micromatrizz[71][446] = 9'b111111111;
assign micromatrizz[71][447] = 9'b111111111;
assign micromatrizz[71][448] = 9'b111111111;
assign micromatrizz[71][449] = 9'b111111111;
assign micromatrizz[71][450] = 9'b111111111;
assign micromatrizz[71][451] = 9'b111111111;
assign micromatrizz[71][452] = 9'b111111111;
assign micromatrizz[71][453] = 9'b111111111;
assign micromatrizz[71][454] = 9'b111111111;
assign micromatrizz[71][455] = 9'b111111111;
assign micromatrizz[71][456] = 9'b111111111;
assign micromatrizz[71][457] = 9'b111111111;
assign micromatrizz[71][458] = 9'b111111111;
assign micromatrizz[71][459] = 9'b111111111;
assign micromatrizz[71][460] = 9'b111111111;
assign micromatrizz[71][461] = 9'b111111111;
assign micromatrizz[71][462] = 9'b111111111;
assign micromatrizz[71][463] = 9'b111111111;
assign micromatrizz[71][464] = 9'b111111111;
assign micromatrizz[71][465] = 9'b111111111;
assign micromatrizz[71][466] = 9'b111111111;
assign micromatrizz[71][467] = 9'b111111111;
assign micromatrizz[71][468] = 9'b111111111;
assign micromatrizz[71][469] = 9'b111111111;
assign micromatrizz[71][470] = 9'b111111111;
assign micromatrizz[71][471] = 9'b111111111;
assign micromatrizz[71][472] = 9'b111111111;
assign micromatrizz[71][473] = 9'b111111111;
assign micromatrizz[71][474] = 9'b111111111;
assign micromatrizz[71][475] = 9'b111111111;
assign micromatrizz[71][476] = 9'b111111111;
assign micromatrizz[71][477] = 9'b111111111;
assign micromatrizz[71][478] = 9'b111111111;
assign micromatrizz[71][479] = 9'b111111111;
assign micromatrizz[71][480] = 9'b111111111;
assign micromatrizz[71][481] = 9'b111111111;
assign micromatrizz[71][482] = 9'b111111111;
assign micromatrizz[71][483] = 9'b111111111;
assign micromatrizz[71][484] = 9'b111111111;
assign micromatrizz[71][485] = 9'b111111111;
assign micromatrizz[71][486] = 9'b111111111;
assign micromatrizz[71][487] = 9'b111111111;
assign micromatrizz[71][488] = 9'b111111111;
assign micromatrizz[71][489] = 9'b111111111;
assign micromatrizz[71][490] = 9'b111111111;
assign micromatrizz[71][491] = 9'b111111111;
assign micromatrizz[71][492] = 9'b111111111;
assign micromatrizz[71][493] = 9'b111111111;
assign micromatrizz[71][494] = 9'b111111111;
assign micromatrizz[71][495] = 9'b111111111;
assign micromatrizz[71][496] = 9'b111111111;
assign micromatrizz[71][497] = 9'b111111111;
assign micromatrizz[71][498] = 9'b111111111;
assign micromatrizz[71][499] = 9'b111111111;
assign micromatrizz[71][500] = 9'b111111111;
assign micromatrizz[71][501] = 9'b111111111;
assign micromatrizz[71][502] = 9'b111111111;
assign micromatrizz[71][503] = 9'b111111111;
assign micromatrizz[71][504] = 9'b111111111;
assign micromatrizz[71][505] = 9'b111111111;
assign micromatrizz[71][506] = 9'b111111111;
assign micromatrizz[71][507] = 9'b111111111;
assign micromatrizz[71][508] = 9'b111111111;
assign micromatrizz[71][509] = 9'b111111111;
assign micromatrizz[71][510] = 9'b111111111;
assign micromatrizz[71][511] = 9'b111111111;
assign micromatrizz[71][512] = 9'b111111111;
assign micromatrizz[71][513] = 9'b111111111;
assign micromatrizz[71][514] = 9'b111111111;
assign micromatrizz[71][515] = 9'b111111111;
assign micromatrizz[71][516] = 9'b111111111;
assign micromatrizz[71][517] = 9'b111111111;
assign micromatrizz[71][518] = 9'b111111111;
assign micromatrizz[71][519] = 9'b111111111;
assign micromatrizz[71][520] = 9'b111111111;
assign micromatrizz[71][521] = 9'b111111111;
assign micromatrizz[71][522] = 9'b111111111;
assign micromatrizz[71][523] = 9'b111111111;
assign micromatrizz[71][524] = 9'b111111111;
assign micromatrizz[71][525] = 9'b111111111;
assign micromatrizz[71][526] = 9'b111111111;
assign micromatrizz[71][527] = 9'b111111111;
assign micromatrizz[71][528] = 9'b111111111;
assign micromatrizz[71][529] = 9'b111111111;
assign micromatrizz[71][530] = 9'b111111111;
assign micromatrizz[71][531] = 9'b111111111;
assign micromatrizz[71][532] = 9'b111111111;
assign micromatrizz[71][533] = 9'b111111111;
assign micromatrizz[71][534] = 9'b111111111;
assign micromatrizz[71][535] = 9'b111111111;
assign micromatrizz[71][536] = 9'b111111111;
assign micromatrizz[71][537] = 9'b111111111;
assign micromatrizz[71][538] = 9'b111111111;
assign micromatrizz[71][539] = 9'b111111111;
assign micromatrizz[71][540] = 9'b111111111;
assign micromatrizz[71][541] = 9'b111111111;
assign micromatrizz[71][542] = 9'b111111111;
assign micromatrizz[71][543] = 9'b111111111;
assign micromatrizz[71][544] = 9'b111111111;
assign micromatrizz[71][545] = 9'b111111111;
assign micromatrizz[71][546] = 9'b111111111;
assign micromatrizz[71][547] = 9'b111111111;
assign micromatrizz[71][548] = 9'b111111111;
assign micromatrizz[71][549] = 9'b111111111;
assign micromatrizz[71][550] = 9'b111111111;
assign micromatrizz[71][551] = 9'b111111111;
assign micromatrizz[71][552] = 9'b111111111;
assign micromatrizz[71][553] = 9'b111111111;
assign micromatrizz[71][554] = 9'b111111111;
assign micromatrizz[71][555] = 9'b111111111;
assign micromatrizz[71][556] = 9'b111111111;
assign micromatrizz[71][557] = 9'b111111111;
assign micromatrizz[71][558] = 9'b111111111;
assign micromatrizz[71][559] = 9'b111111111;
assign micromatrizz[71][560] = 9'b111111111;
assign micromatrizz[71][561] = 9'b111111111;
assign micromatrizz[71][562] = 9'b111111111;
assign micromatrizz[71][563] = 9'b111111111;
assign micromatrizz[71][564] = 9'b111111111;
assign micromatrizz[71][565] = 9'b111111111;
assign micromatrizz[71][566] = 9'b111111111;
assign micromatrizz[71][567] = 9'b111111111;
assign micromatrizz[71][568] = 9'b111111111;
assign micromatrizz[71][569] = 9'b111111111;
assign micromatrizz[71][570] = 9'b111111111;
assign micromatrizz[71][571] = 9'b111111111;
assign micromatrizz[71][572] = 9'b111111111;
assign micromatrizz[71][573] = 9'b111111111;
assign micromatrizz[71][574] = 9'b111111111;
assign micromatrizz[71][575] = 9'b111111111;
assign micromatrizz[71][576] = 9'b111111111;
assign micromatrizz[71][577] = 9'b111111111;
assign micromatrizz[71][578] = 9'b111111111;
assign micromatrizz[71][579] = 9'b111111111;
assign micromatrizz[71][580] = 9'b111111111;
assign micromatrizz[71][581] = 9'b111111111;
assign micromatrizz[71][582] = 9'b111111111;
assign micromatrizz[71][583] = 9'b111111111;
assign micromatrizz[71][584] = 9'b111111111;
assign micromatrizz[71][585] = 9'b111111111;
assign micromatrizz[71][586] = 9'b111111111;
assign micromatrizz[71][587] = 9'b111111111;
assign micromatrizz[71][588] = 9'b111111111;
assign micromatrizz[71][589] = 9'b111111111;
assign micromatrizz[71][590] = 9'b111111111;
assign micromatrizz[71][591] = 9'b111111111;
assign micromatrizz[71][592] = 9'b111111111;
assign micromatrizz[71][593] = 9'b111111111;
assign micromatrizz[71][594] = 9'b111111111;
assign micromatrizz[71][595] = 9'b111111111;
assign micromatrizz[71][596] = 9'b111111111;
assign micromatrizz[71][597] = 9'b111111111;
assign micromatrizz[71][598] = 9'b111111111;
assign micromatrizz[71][599] = 9'b111111111;
assign micromatrizz[71][600] = 9'b111111111;
assign micromatrizz[71][601] = 9'b111111111;
assign micromatrizz[71][602] = 9'b111111111;
assign micromatrizz[71][603] = 9'b111111111;
assign micromatrizz[71][604] = 9'b111111111;
assign micromatrizz[71][605] = 9'b111111111;
assign micromatrizz[71][606] = 9'b111111111;
assign micromatrizz[71][607] = 9'b111111111;
assign micromatrizz[71][608] = 9'b111111111;
assign micromatrizz[71][609] = 9'b111111111;
assign micromatrizz[71][610] = 9'b111111111;
assign micromatrizz[71][611] = 9'b111111111;
assign micromatrizz[71][612] = 9'b111111111;
assign micromatrizz[71][613] = 9'b111111111;
assign micromatrizz[71][614] = 9'b111111111;
assign micromatrizz[71][615] = 9'b111111111;
assign micromatrizz[71][616] = 9'b111111111;
assign micromatrizz[71][617] = 9'b111111111;
assign micromatrizz[71][618] = 9'b111111111;
assign micromatrizz[71][619] = 9'b111111111;
assign micromatrizz[71][620] = 9'b111111111;
assign micromatrizz[71][621] = 9'b111111111;
assign micromatrizz[71][622] = 9'b111111111;
assign micromatrizz[71][623] = 9'b111111111;
assign micromatrizz[71][624] = 9'b111111111;
assign micromatrizz[71][625] = 9'b111111111;
assign micromatrizz[71][626] = 9'b111111111;
assign micromatrizz[71][627] = 9'b111111111;
assign micromatrizz[71][628] = 9'b111111111;
assign micromatrizz[71][629] = 9'b111111111;
assign micromatrizz[71][630] = 9'b111111111;
assign micromatrizz[71][631] = 9'b111111111;
assign micromatrizz[71][632] = 9'b111111111;
assign micromatrizz[71][633] = 9'b111111111;
assign micromatrizz[71][634] = 9'b111111111;
assign micromatrizz[71][635] = 9'b111111111;
assign micromatrizz[71][636] = 9'b111111111;
assign micromatrizz[71][637] = 9'b111111111;
assign micromatrizz[71][638] = 9'b111111111;
assign micromatrizz[71][639] = 9'b111111111;
assign micromatrizz[72][0] = 9'b111111111;
assign micromatrizz[72][1] = 9'b111111111;
assign micromatrizz[72][2] = 9'b111111111;
assign micromatrizz[72][3] = 9'b111111111;
assign micromatrizz[72][4] = 9'b111111111;
assign micromatrizz[72][5] = 9'b111111111;
assign micromatrizz[72][6] = 9'b111111111;
assign micromatrizz[72][7] = 9'b111111111;
assign micromatrizz[72][8] = 9'b111111111;
assign micromatrizz[72][9] = 9'b111111111;
assign micromatrizz[72][10] = 9'b111111111;
assign micromatrizz[72][11] = 9'b111111111;
assign micromatrizz[72][12] = 9'b111111111;
assign micromatrizz[72][13] = 9'b111111111;
assign micromatrizz[72][14] = 9'b111111111;
assign micromatrizz[72][15] = 9'b111111111;
assign micromatrizz[72][16] = 9'b111111111;
assign micromatrizz[72][17] = 9'b111111111;
assign micromatrizz[72][18] = 9'b111111111;
assign micromatrizz[72][19] = 9'b111111111;
assign micromatrizz[72][20] = 9'b111111111;
assign micromatrizz[72][21] = 9'b111111111;
assign micromatrizz[72][22] = 9'b111111111;
assign micromatrizz[72][23] = 9'b111111111;
assign micromatrizz[72][24] = 9'b111111111;
assign micromatrizz[72][25] = 9'b111111111;
assign micromatrizz[72][26] = 9'b111111111;
assign micromatrizz[72][27] = 9'b111111111;
assign micromatrizz[72][28] = 9'b111111111;
assign micromatrizz[72][29] = 9'b111111111;
assign micromatrizz[72][30] = 9'b111111111;
assign micromatrizz[72][31] = 9'b111111111;
assign micromatrizz[72][32] = 9'b111111111;
assign micromatrizz[72][33] = 9'b111111111;
assign micromatrizz[72][34] = 9'b111111111;
assign micromatrizz[72][35] = 9'b111111111;
assign micromatrizz[72][36] = 9'b111111111;
assign micromatrizz[72][37] = 9'b111111111;
assign micromatrizz[72][38] = 9'b111111111;
assign micromatrizz[72][39] = 9'b111111111;
assign micromatrizz[72][40] = 9'b111111111;
assign micromatrizz[72][41] = 9'b111111111;
assign micromatrizz[72][42] = 9'b111111111;
assign micromatrizz[72][43] = 9'b111111111;
assign micromatrizz[72][44] = 9'b111111111;
assign micromatrizz[72][45] = 9'b111111111;
assign micromatrizz[72][46] = 9'b111111111;
assign micromatrizz[72][47] = 9'b111111111;
assign micromatrizz[72][48] = 9'b111111111;
assign micromatrizz[72][49] = 9'b111111111;
assign micromatrizz[72][50] = 9'b111111111;
assign micromatrizz[72][51] = 9'b111111111;
assign micromatrizz[72][52] = 9'b111111111;
assign micromatrizz[72][53] = 9'b111111111;
assign micromatrizz[72][54] = 9'b111111111;
assign micromatrizz[72][55] = 9'b111111111;
assign micromatrizz[72][56] = 9'b111111111;
assign micromatrizz[72][57] = 9'b111111111;
assign micromatrizz[72][58] = 9'b111111111;
assign micromatrizz[72][59] = 9'b111111111;
assign micromatrizz[72][60] = 9'b111111111;
assign micromatrizz[72][61] = 9'b111111111;
assign micromatrizz[72][62] = 9'b111111111;
assign micromatrizz[72][63] = 9'b111111111;
assign micromatrizz[72][64] = 9'b111111111;
assign micromatrizz[72][65] = 9'b111111111;
assign micromatrizz[72][66] = 9'b111111111;
assign micromatrizz[72][67] = 9'b111111111;
assign micromatrizz[72][68] = 9'b111111111;
assign micromatrizz[72][69] = 9'b111111111;
assign micromatrizz[72][70] = 9'b111111111;
assign micromatrizz[72][71] = 9'b111111111;
assign micromatrizz[72][72] = 9'b111111111;
assign micromatrizz[72][73] = 9'b111111111;
assign micromatrizz[72][74] = 9'b111111111;
assign micromatrizz[72][75] = 9'b111111111;
assign micromatrizz[72][76] = 9'b111111111;
assign micromatrizz[72][77] = 9'b111111111;
assign micromatrizz[72][78] = 9'b111111111;
assign micromatrizz[72][79] = 9'b111111111;
assign micromatrizz[72][80] = 9'b111111111;
assign micromatrizz[72][81] = 9'b111111111;
assign micromatrizz[72][82] = 9'b111111111;
assign micromatrizz[72][83] = 9'b111111111;
assign micromatrizz[72][84] = 9'b111111111;
assign micromatrizz[72][85] = 9'b111111111;
assign micromatrizz[72][86] = 9'b111111111;
assign micromatrizz[72][87] = 9'b111111111;
assign micromatrizz[72][88] = 9'b111111111;
assign micromatrizz[72][89] = 9'b111111111;
assign micromatrizz[72][90] = 9'b111111111;
assign micromatrizz[72][91] = 9'b111111111;
assign micromatrizz[72][92] = 9'b111111111;
assign micromatrizz[72][93] = 9'b111111111;
assign micromatrizz[72][94] = 9'b111111111;
assign micromatrizz[72][95] = 9'b111111111;
assign micromatrizz[72][96] = 9'b111111111;
assign micromatrizz[72][97] = 9'b111111111;
assign micromatrizz[72][98] = 9'b111111111;
assign micromatrizz[72][99] = 9'b111111111;
assign micromatrizz[72][100] = 9'b111111111;
assign micromatrizz[72][101] = 9'b111111111;
assign micromatrizz[72][102] = 9'b111111111;
assign micromatrizz[72][103] = 9'b111111111;
assign micromatrizz[72][104] = 9'b111111111;
assign micromatrizz[72][105] = 9'b111111111;
assign micromatrizz[72][106] = 9'b111111111;
assign micromatrizz[72][107] = 9'b111111111;
assign micromatrizz[72][108] = 9'b111111111;
assign micromatrizz[72][109] = 9'b111111111;
assign micromatrizz[72][110] = 9'b111111111;
assign micromatrizz[72][111] = 9'b111111111;
assign micromatrizz[72][112] = 9'b111111111;
assign micromatrizz[72][113] = 9'b111111111;
assign micromatrizz[72][114] = 9'b111111111;
assign micromatrizz[72][115] = 9'b111111111;
assign micromatrizz[72][116] = 9'b111111111;
assign micromatrizz[72][117] = 9'b111111111;
assign micromatrizz[72][118] = 9'b111111111;
assign micromatrizz[72][119] = 9'b111111111;
assign micromatrizz[72][120] = 9'b111111111;
assign micromatrizz[72][121] = 9'b111111111;
assign micromatrizz[72][122] = 9'b111111111;
assign micromatrizz[72][123] = 9'b111111111;
assign micromatrizz[72][124] = 9'b111111111;
assign micromatrizz[72][125] = 9'b111111111;
assign micromatrizz[72][126] = 9'b111111111;
assign micromatrizz[72][127] = 9'b111111111;
assign micromatrizz[72][128] = 9'b111111111;
assign micromatrizz[72][129] = 9'b111111111;
assign micromatrizz[72][130] = 9'b111111111;
assign micromatrizz[72][131] = 9'b111111111;
assign micromatrizz[72][132] = 9'b111111111;
assign micromatrizz[72][133] = 9'b111111111;
assign micromatrizz[72][134] = 9'b111111111;
assign micromatrizz[72][135] = 9'b111111111;
assign micromatrizz[72][136] = 9'b111111111;
assign micromatrizz[72][137] = 9'b111111111;
assign micromatrizz[72][138] = 9'b111111111;
assign micromatrizz[72][139] = 9'b111111111;
assign micromatrizz[72][140] = 9'b111111111;
assign micromatrizz[72][141] = 9'b111111111;
assign micromatrizz[72][142] = 9'b111111111;
assign micromatrizz[72][143] = 9'b111111111;
assign micromatrizz[72][144] = 9'b111111111;
assign micromatrizz[72][145] = 9'b111111111;
assign micromatrizz[72][146] = 9'b111111111;
assign micromatrizz[72][147] = 9'b111111111;
assign micromatrizz[72][148] = 9'b111111111;
assign micromatrizz[72][149] = 9'b111111111;
assign micromatrizz[72][150] = 9'b111111111;
assign micromatrizz[72][151] = 9'b111111111;
assign micromatrizz[72][152] = 9'b111111111;
assign micromatrizz[72][153] = 9'b111111111;
assign micromatrizz[72][154] = 9'b111111111;
assign micromatrizz[72][155] = 9'b111111111;
assign micromatrizz[72][156] = 9'b111111111;
assign micromatrizz[72][157] = 9'b111111111;
assign micromatrizz[72][158] = 9'b111111111;
assign micromatrizz[72][159] = 9'b111111111;
assign micromatrizz[72][160] = 9'b111111111;
assign micromatrizz[72][161] = 9'b111111111;
assign micromatrizz[72][162] = 9'b111111111;
assign micromatrizz[72][163] = 9'b111111111;
assign micromatrizz[72][164] = 9'b111111111;
assign micromatrizz[72][165] = 9'b111111111;
assign micromatrizz[72][166] = 9'b111111111;
assign micromatrizz[72][167] = 9'b111111111;
assign micromatrizz[72][168] = 9'b111111111;
assign micromatrizz[72][169] = 9'b111111111;
assign micromatrizz[72][170] = 9'b111111111;
assign micromatrizz[72][171] = 9'b111111111;
assign micromatrizz[72][172] = 9'b111111111;
assign micromatrizz[72][173] = 9'b111111111;
assign micromatrizz[72][174] = 9'b111111111;
assign micromatrizz[72][175] = 9'b111111111;
assign micromatrizz[72][176] = 9'b111111111;
assign micromatrizz[72][177] = 9'b111111111;
assign micromatrizz[72][178] = 9'b111111111;
assign micromatrizz[72][179] = 9'b111111111;
assign micromatrizz[72][180] = 9'b111111111;
assign micromatrizz[72][181] = 9'b111111111;
assign micromatrizz[72][182] = 9'b111111111;
assign micromatrizz[72][183] = 9'b111111111;
assign micromatrizz[72][184] = 9'b111111111;
assign micromatrizz[72][185] = 9'b111111111;
assign micromatrizz[72][186] = 9'b111111111;
assign micromatrizz[72][187] = 9'b111111111;
assign micromatrizz[72][188] = 9'b111111111;
assign micromatrizz[72][189] = 9'b111111111;
assign micromatrizz[72][190] = 9'b111111111;
assign micromatrizz[72][191] = 9'b111111111;
assign micromatrizz[72][192] = 9'b111111111;
assign micromatrizz[72][193] = 9'b111111111;
assign micromatrizz[72][194] = 9'b111111111;
assign micromatrizz[72][195] = 9'b111111111;
assign micromatrizz[72][196] = 9'b111111111;
assign micromatrizz[72][197] = 9'b111111111;
assign micromatrizz[72][198] = 9'b111111111;
assign micromatrizz[72][199] = 9'b111111111;
assign micromatrizz[72][200] = 9'b111111111;
assign micromatrizz[72][201] = 9'b111111111;
assign micromatrizz[72][202] = 9'b111111111;
assign micromatrizz[72][203] = 9'b111111111;
assign micromatrizz[72][204] = 9'b111111111;
assign micromatrizz[72][205] = 9'b111111111;
assign micromatrizz[72][206] = 9'b111111111;
assign micromatrizz[72][207] = 9'b111111111;
assign micromatrizz[72][208] = 9'b111111111;
assign micromatrizz[72][209] = 9'b111111111;
assign micromatrizz[72][210] = 9'b111111111;
assign micromatrizz[72][211] = 9'b111111111;
assign micromatrizz[72][212] = 9'b111111111;
assign micromatrizz[72][213] = 9'b111111111;
assign micromatrizz[72][214] = 9'b111111111;
assign micromatrizz[72][215] = 9'b111111111;
assign micromatrizz[72][216] = 9'b111111111;
assign micromatrizz[72][217] = 9'b111111111;
assign micromatrizz[72][218] = 9'b111111111;
assign micromatrizz[72][219] = 9'b111111111;
assign micromatrizz[72][220] = 9'b111111111;
assign micromatrizz[72][221] = 9'b111111111;
assign micromatrizz[72][222] = 9'b111111111;
assign micromatrizz[72][223] = 9'b111111111;
assign micromatrizz[72][224] = 9'b111111111;
assign micromatrizz[72][225] = 9'b111111111;
assign micromatrizz[72][226] = 9'b111111111;
assign micromatrizz[72][227] = 9'b111111111;
assign micromatrizz[72][228] = 9'b111111111;
assign micromatrizz[72][229] = 9'b111111111;
assign micromatrizz[72][230] = 9'b111111111;
assign micromatrizz[72][231] = 9'b111111111;
assign micromatrizz[72][232] = 9'b111111111;
assign micromatrizz[72][233] = 9'b111111111;
assign micromatrizz[72][234] = 9'b111111111;
assign micromatrizz[72][235] = 9'b111111111;
assign micromatrizz[72][236] = 9'b111111111;
assign micromatrizz[72][237] = 9'b111111111;
assign micromatrizz[72][238] = 9'b111111111;
assign micromatrizz[72][239] = 9'b111111111;
assign micromatrizz[72][240] = 9'b111111111;
assign micromatrizz[72][241] = 9'b111111111;
assign micromatrizz[72][242] = 9'b111111111;
assign micromatrizz[72][243] = 9'b111111111;
assign micromatrizz[72][244] = 9'b111111111;
assign micromatrizz[72][245] = 9'b111111111;
assign micromatrizz[72][246] = 9'b111111111;
assign micromatrizz[72][247] = 9'b111111111;
assign micromatrizz[72][248] = 9'b111111111;
assign micromatrizz[72][249] = 9'b111111111;
assign micromatrizz[72][250] = 9'b111111111;
assign micromatrizz[72][251] = 9'b111111111;
assign micromatrizz[72][252] = 9'b111111111;
assign micromatrizz[72][253] = 9'b111111111;
assign micromatrizz[72][254] = 9'b111111111;
assign micromatrizz[72][255] = 9'b111111111;
assign micromatrizz[72][256] = 9'b111111111;
assign micromatrizz[72][257] = 9'b111111111;
assign micromatrizz[72][258] = 9'b111111111;
assign micromatrizz[72][259] = 9'b111111111;
assign micromatrizz[72][260] = 9'b111111111;
assign micromatrizz[72][261] = 9'b111111111;
assign micromatrizz[72][262] = 9'b111111111;
assign micromatrizz[72][263] = 9'b111111111;
assign micromatrizz[72][264] = 9'b111111111;
assign micromatrizz[72][265] = 9'b111111111;
assign micromatrizz[72][266] = 9'b111111111;
assign micromatrizz[72][267] = 9'b111111111;
assign micromatrizz[72][268] = 9'b111111111;
assign micromatrizz[72][269] = 9'b111111111;
assign micromatrizz[72][270] = 9'b111111111;
assign micromatrizz[72][271] = 9'b111111111;
assign micromatrizz[72][272] = 9'b111111111;
assign micromatrizz[72][273] = 9'b111111111;
assign micromatrizz[72][274] = 9'b111111111;
assign micromatrizz[72][275] = 9'b111111111;
assign micromatrizz[72][276] = 9'b111111111;
assign micromatrizz[72][277] = 9'b111111111;
assign micromatrizz[72][278] = 9'b111111111;
assign micromatrizz[72][279] = 9'b111111111;
assign micromatrizz[72][280] = 9'b111111111;
assign micromatrizz[72][281] = 9'b111111111;
assign micromatrizz[72][282] = 9'b111111111;
assign micromatrizz[72][283] = 9'b111111111;
assign micromatrizz[72][284] = 9'b111111111;
assign micromatrizz[72][285] = 9'b111111111;
assign micromatrizz[72][286] = 9'b111111111;
assign micromatrizz[72][287] = 9'b111111111;
assign micromatrizz[72][288] = 9'b111111111;
assign micromatrizz[72][289] = 9'b111111111;
assign micromatrizz[72][290] = 9'b111111111;
assign micromatrizz[72][291] = 9'b111111111;
assign micromatrizz[72][292] = 9'b111111111;
assign micromatrizz[72][293] = 9'b111111111;
assign micromatrizz[72][294] = 9'b111111111;
assign micromatrizz[72][295] = 9'b111111111;
assign micromatrizz[72][296] = 9'b111111111;
assign micromatrizz[72][297] = 9'b111111111;
assign micromatrizz[72][298] = 9'b111111111;
assign micromatrizz[72][299] = 9'b111111111;
assign micromatrizz[72][300] = 9'b111111111;
assign micromatrizz[72][301] = 9'b111111111;
assign micromatrizz[72][302] = 9'b111111111;
assign micromatrizz[72][303] = 9'b111111111;
assign micromatrizz[72][304] = 9'b111111111;
assign micromatrizz[72][305] = 9'b111111111;
assign micromatrizz[72][306] = 9'b111111111;
assign micromatrizz[72][307] = 9'b111111111;
assign micromatrizz[72][308] = 9'b111111111;
assign micromatrizz[72][309] = 9'b111111111;
assign micromatrizz[72][310] = 9'b111111111;
assign micromatrizz[72][311] = 9'b111111111;
assign micromatrizz[72][312] = 9'b111111111;
assign micromatrizz[72][313] = 9'b111111111;
assign micromatrizz[72][314] = 9'b111111111;
assign micromatrizz[72][315] = 9'b111111111;
assign micromatrizz[72][316] = 9'b111111111;
assign micromatrizz[72][317] = 9'b111111111;
assign micromatrizz[72][318] = 9'b111111111;
assign micromatrizz[72][319] = 9'b111111111;
assign micromatrizz[72][320] = 9'b111111111;
assign micromatrizz[72][321] = 9'b111111111;
assign micromatrizz[72][322] = 9'b111111111;
assign micromatrizz[72][323] = 9'b111111111;
assign micromatrizz[72][324] = 9'b111111111;
assign micromatrizz[72][325] = 9'b111111111;
assign micromatrizz[72][326] = 9'b111111111;
assign micromatrizz[72][327] = 9'b111111111;
assign micromatrizz[72][328] = 9'b111111111;
assign micromatrizz[72][329] = 9'b111111111;
assign micromatrizz[72][330] = 9'b111111111;
assign micromatrizz[72][331] = 9'b111111111;
assign micromatrizz[72][332] = 9'b111111111;
assign micromatrizz[72][333] = 9'b111111111;
assign micromatrizz[72][334] = 9'b111111111;
assign micromatrizz[72][335] = 9'b111111111;
assign micromatrizz[72][336] = 9'b111111111;
assign micromatrizz[72][337] = 9'b111111111;
assign micromatrizz[72][338] = 9'b111111111;
assign micromatrizz[72][339] = 9'b111111111;
assign micromatrizz[72][340] = 9'b111111111;
assign micromatrizz[72][341] = 9'b111111111;
assign micromatrizz[72][342] = 9'b111111111;
assign micromatrizz[72][343] = 9'b111111111;
assign micromatrizz[72][344] = 9'b111111111;
assign micromatrizz[72][345] = 9'b111111111;
assign micromatrizz[72][346] = 9'b111111111;
assign micromatrizz[72][347] = 9'b111111111;
assign micromatrizz[72][348] = 9'b111111111;
assign micromatrizz[72][349] = 9'b111111111;
assign micromatrizz[72][350] = 9'b111111111;
assign micromatrizz[72][351] = 9'b111111111;
assign micromatrizz[72][352] = 9'b111111111;
assign micromatrizz[72][353] = 9'b111111111;
assign micromatrizz[72][354] = 9'b111111111;
assign micromatrizz[72][355] = 9'b111111111;
assign micromatrizz[72][356] = 9'b111111111;
assign micromatrizz[72][357] = 9'b111111111;
assign micromatrizz[72][358] = 9'b111111111;
assign micromatrizz[72][359] = 9'b111111111;
assign micromatrizz[72][360] = 9'b111111111;
assign micromatrizz[72][361] = 9'b111111111;
assign micromatrizz[72][362] = 9'b111111111;
assign micromatrizz[72][363] = 9'b111111111;
assign micromatrizz[72][364] = 9'b111111111;
assign micromatrizz[72][365] = 9'b111111111;
assign micromatrizz[72][366] = 9'b111111111;
assign micromatrizz[72][367] = 9'b111111111;
assign micromatrizz[72][368] = 9'b111111111;
assign micromatrizz[72][369] = 9'b111111111;
assign micromatrizz[72][370] = 9'b111111111;
assign micromatrizz[72][371] = 9'b111111111;
assign micromatrizz[72][372] = 9'b111111111;
assign micromatrizz[72][373] = 9'b111111111;
assign micromatrizz[72][374] = 9'b111111111;
assign micromatrizz[72][375] = 9'b111111111;
assign micromatrizz[72][376] = 9'b111111111;
assign micromatrizz[72][377] = 9'b111111111;
assign micromatrizz[72][378] = 9'b111111111;
assign micromatrizz[72][379] = 9'b111111111;
assign micromatrizz[72][380] = 9'b111111111;
assign micromatrizz[72][381] = 9'b111111111;
assign micromatrizz[72][382] = 9'b111111111;
assign micromatrizz[72][383] = 9'b111111111;
assign micromatrizz[72][384] = 9'b111111111;
assign micromatrizz[72][385] = 9'b111111111;
assign micromatrizz[72][386] = 9'b111111111;
assign micromatrizz[72][387] = 9'b111111111;
assign micromatrizz[72][388] = 9'b111111111;
assign micromatrizz[72][389] = 9'b111111111;
assign micromatrizz[72][390] = 9'b111111111;
assign micromatrizz[72][391] = 9'b111111111;
assign micromatrizz[72][392] = 9'b111111111;
assign micromatrizz[72][393] = 9'b111111111;
assign micromatrizz[72][394] = 9'b111111111;
assign micromatrizz[72][395] = 9'b111111111;
assign micromatrizz[72][396] = 9'b111111111;
assign micromatrizz[72][397] = 9'b111111111;
assign micromatrizz[72][398] = 9'b111111111;
assign micromatrizz[72][399] = 9'b111111111;
assign micromatrizz[72][400] = 9'b111111111;
assign micromatrizz[72][401] = 9'b111111111;
assign micromatrizz[72][402] = 9'b111111111;
assign micromatrizz[72][403] = 9'b111111111;
assign micromatrizz[72][404] = 9'b111111111;
assign micromatrizz[72][405] = 9'b111111111;
assign micromatrizz[72][406] = 9'b111111111;
assign micromatrizz[72][407] = 9'b111111111;
assign micromatrizz[72][408] = 9'b111111111;
assign micromatrizz[72][409] = 9'b111111111;
assign micromatrizz[72][410] = 9'b111111111;
assign micromatrizz[72][411] = 9'b111111111;
assign micromatrizz[72][412] = 9'b111111111;
assign micromatrizz[72][413] = 9'b111111111;
assign micromatrizz[72][414] = 9'b111111111;
assign micromatrizz[72][415] = 9'b111111111;
assign micromatrizz[72][416] = 9'b111111111;
assign micromatrizz[72][417] = 9'b111111111;
assign micromatrizz[72][418] = 9'b111111111;
assign micromatrizz[72][419] = 9'b111111111;
assign micromatrizz[72][420] = 9'b111111111;
assign micromatrizz[72][421] = 9'b111111111;
assign micromatrizz[72][422] = 9'b111111111;
assign micromatrizz[72][423] = 9'b111111111;
assign micromatrizz[72][424] = 9'b111111111;
assign micromatrizz[72][425] = 9'b111111111;
assign micromatrizz[72][426] = 9'b111111111;
assign micromatrizz[72][427] = 9'b111111111;
assign micromatrizz[72][428] = 9'b111111111;
assign micromatrizz[72][429] = 9'b111111111;
assign micromatrizz[72][430] = 9'b111111111;
assign micromatrizz[72][431] = 9'b111111111;
assign micromatrizz[72][432] = 9'b111111111;
assign micromatrizz[72][433] = 9'b111111111;
assign micromatrizz[72][434] = 9'b111111111;
assign micromatrizz[72][435] = 9'b111111111;
assign micromatrizz[72][436] = 9'b111111111;
assign micromatrizz[72][437] = 9'b111111111;
assign micromatrizz[72][438] = 9'b111111111;
assign micromatrizz[72][439] = 9'b111111111;
assign micromatrizz[72][440] = 9'b111111111;
assign micromatrizz[72][441] = 9'b111111111;
assign micromatrizz[72][442] = 9'b111111111;
assign micromatrizz[72][443] = 9'b111111111;
assign micromatrizz[72][444] = 9'b111111111;
assign micromatrizz[72][445] = 9'b111111111;
assign micromatrizz[72][446] = 9'b111111111;
assign micromatrizz[72][447] = 9'b111111111;
assign micromatrizz[72][448] = 9'b111111111;
assign micromatrizz[72][449] = 9'b111111111;
assign micromatrizz[72][450] = 9'b111111111;
assign micromatrizz[72][451] = 9'b111111111;
assign micromatrizz[72][452] = 9'b111111111;
assign micromatrizz[72][453] = 9'b111111111;
assign micromatrizz[72][454] = 9'b111111111;
assign micromatrizz[72][455] = 9'b111111111;
assign micromatrizz[72][456] = 9'b111111111;
assign micromatrizz[72][457] = 9'b111111111;
assign micromatrizz[72][458] = 9'b111111111;
assign micromatrizz[72][459] = 9'b111111111;
assign micromatrizz[72][460] = 9'b111111111;
assign micromatrizz[72][461] = 9'b111111111;
assign micromatrizz[72][462] = 9'b111111111;
assign micromatrizz[72][463] = 9'b111111111;
assign micromatrizz[72][464] = 9'b111111111;
assign micromatrizz[72][465] = 9'b111111111;
assign micromatrizz[72][466] = 9'b111111111;
assign micromatrizz[72][467] = 9'b111111111;
assign micromatrizz[72][468] = 9'b111111111;
assign micromatrizz[72][469] = 9'b111111111;
assign micromatrizz[72][470] = 9'b111111111;
assign micromatrizz[72][471] = 9'b111111111;
assign micromatrizz[72][472] = 9'b111111111;
assign micromatrizz[72][473] = 9'b111111111;
assign micromatrizz[72][474] = 9'b111111111;
assign micromatrizz[72][475] = 9'b111111111;
assign micromatrizz[72][476] = 9'b111111111;
assign micromatrizz[72][477] = 9'b111111111;
assign micromatrizz[72][478] = 9'b111111111;
assign micromatrizz[72][479] = 9'b111111111;
assign micromatrizz[72][480] = 9'b111111111;
assign micromatrizz[72][481] = 9'b111111111;
assign micromatrizz[72][482] = 9'b111111111;
assign micromatrizz[72][483] = 9'b111111111;
assign micromatrizz[72][484] = 9'b111111111;
assign micromatrizz[72][485] = 9'b111111111;
assign micromatrizz[72][486] = 9'b111111111;
assign micromatrizz[72][487] = 9'b111111111;
assign micromatrizz[72][488] = 9'b111111111;
assign micromatrizz[72][489] = 9'b111111111;
assign micromatrizz[72][490] = 9'b111111111;
assign micromatrizz[72][491] = 9'b111111111;
assign micromatrizz[72][492] = 9'b111111111;
assign micromatrizz[72][493] = 9'b111111111;
assign micromatrizz[72][494] = 9'b111111111;
assign micromatrizz[72][495] = 9'b111111111;
assign micromatrizz[72][496] = 9'b111111111;
assign micromatrizz[72][497] = 9'b111111111;
assign micromatrizz[72][498] = 9'b111111111;
assign micromatrizz[72][499] = 9'b111111111;
assign micromatrizz[72][500] = 9'b111111111;
assign micromatrizz[72][501] = 9'b111111111;
assign micromatrizz[72][502] = 9'b111111111;
assign micromatrizz[72][503] = 9'b111111111;
assign micromatrizz[72][504] = 9'b111111111;
assign micromatrizz[72][505] = 9'b111111111;
assign micromatrizz[72][506] = 9'b111111111;
assign micromatrizz[72][507] = 9'b111111111;
assign micromatrizz[72][508] = 9'b111111111;
assign micromatrizz[72][509] = 9'b111111111;
assign micromatrizz[72][510] = 9'b111111111;
assign micromatrizz[72][511] = 9'b111111111;
assign micromatrizz[72][512] = 9'b111111111;
assign micromatrizz[72][513] = 9'b111111111;
assign micromatrizz[72][514] = 9'b111111111;
assign micromatrizz[72][515] = 9'b111111111;
assign micromatrizz[72][516] = 9'b111111111;
assign micromatrizz[72][517] = 9'b111111111;
assign micromatrizz[72][518] = 9'b111111111;
assign micromatrizz[72][519] = 9'b111111111;
assign micromatrizz[72][520] = 9'b111111111;
assign micromatrizz[72][521] = 9'b111111111;
assign micromatrizz[72][522] = 9'b111111111;
assign micromatrizz[72][523] = 9'b111111111;
assign micromatrizz[72][524] = 9'b111111111;
assign micromatrizz[72][525] = 9'b111111111;
assign micromatrizz[72][526] = 9'b111111111;
assign micromatrizz[72][527] = 9'b111111111;
assign micromatrizz[72][528] = 9'b111111111;
assign micromatrizz[72][529] = 9'b111111111;
assign micromatrizz[72][530] = 9'b111111111;
assign micromatrizz[72][531] = 9'b111111111;
assign micromatrizz[72][532] = 9'b111111111;
assign micromatrizz[72][533] = 9'b111111111;
assign micromatrizz[72][534] = 9'b111111111;
assign micromatrizz[72][535] = 9'b111111111;
assign micromatrizz[72][536] = 9'b111111111;
assign micromatrizz[72][537] = 9'b111111111;
assign micromatrizz[72][538] = 9'b111111111;
assign micromatrizz[72][539] = 9'b111111111;
assign micromatrizz[72][540] = 9'b111111111;
assign micromatrizz[72][541] = 9'b111111111;
assign micromatrizz[72][542] = 9'b111111111;
assign micromatrizz[72][543] = 9'b111111111;
assign micromatrizz[72][544] = 9'b111111111;
assign micromatrizz[72][545] = 9'b111111111;
assign micromatrizz[72][546] = 9'b111111111;
assign micromatrizz[72][547] = 9'b111111111;
assign micromatrizz[72][548] = 9'b111111111;
assign micromatrizz[72][549] = 9'b111111111;
assign micromatrizz[72][550] = 9'b111111111;
assign micromatrizz[72][551] = 9'b111111111;
assign micromatrizz[72][552] = 9'b111111111;
assign micromatrizz[72][553] = 9'b111111111;
assign micromatrizz[72][554] = 9'b111111111;
assign micromatrizz[72][555] = 9'b111111111;
assign micromatrizz[72][556] = 9'b111111111;
assign micromatrizz[72][557] = 9'b111111111;
assign micromatrizz[72][558] = 9'b111111111;
assign micromatrizz[72][559] = 9'b111111111;
assign micromatrizz[72][560] = 9'b111111111;
assign micromatrizz[72][561] = 9'b111111111;
assign micromatrizz[72][562] = 9'b111111111;
assign micromatrizz[72][563] = 9'b111111111;
assign micromatrizz[72][564] = 9'b111111111;
assign micromatrizz[72][565] = 9'b111111111;
assign micromatrizz[72][566] = 9'b111111111;
assign micromatrizz[72][567] = 9'b111111111;
assign micromatrizz[72][568] = 9'b111111111;
assign micromatrizz[72][569] = 9'b111111111;
assign micromatrizz[72][570] = 9'b111111111;
assign micromatrizz[72][571] = 9'b111111111;
assign micromatrizz[72][572] = 9'b111111111;
assign micromatrizz[72][573] = 9'b111111111;
assign micromatrizz[72][574] = 9'b111111111;
assign micromatrizz[72][575] = 9'b111111111;
assign micromatrizz[72][576] = 9'b111111111;
assign micromatrizz[72][577] = 9'b111111111;
assign micromatrizz[72][578] = 9'b111111111;
assign micromatrizz[72][579] = 9'b111111111;
assign micromatrizz[72][580] = 9'b111111111;
assign micromatrizz[72][581] = 9'b111111111;
assign micromatrizz[72][582] = 9'b111111111;
assign micromatrizz[72][583] = 9'b111111111;
assign micromatrizz[72][584] = 9'b111111111;
assign micromatrizz[72][585] = 9'b111111111;
assign micromatrizz[72][586] = 9'b111111111;
assign micromatrizz[72][587] = 9'b111111111;
assign micromatrizz[72][588] = 9'b111111111;
assign micromatrizz[72][589] = 9'b111111111;
assign micromatrizz[72][590] = 9'b111111111;
assign micromatrizz[72][591] = 9'b111111111;
assign micromatrizz[72][592] = 9'b111111111;
assign micromatrizz[72][593] = 9'b111111111;
assign micromatrizz[72][594] = 9'b111111111;
assign micromatrizz[72][595] = 9'b111111111;
assign micromatrizz[72][596] = 9'b111111111;
assign micromatrizz[72][597] = 9'b111111111;
assign micromatrizz[72][598] = 9'b111111111;
assign micromatrizz[72][599] = 9'b111111111;
assign micromatrizz[72][600] = 9'b111111111;
assign micromatrizz[72][601] = 9'b111111111;
assign micromatrizz[72][602] = 9'b111111111;
assign micromatrizz[72][603] = 9'b111111111;
assign micromatrizz[72][604] = 9'b111111111;
assign micromatrizz[72][605] = 9'b111111111;
assign micromatrizz[72][606] = 9'b111111111;
assign micromatrizz[72][607] = 9'b111111111;
assign micromatrizz[72][608] = 9'b111111111;
assign micromatrizz[72][609] = 9'b111111111;
assign micromatrizz[72][610] = 9'b111111111;
assign micromatrizz[72][611] = 9'b111111111;
assign micromatrizz[72][612] = 9'b111111111;
assign micromatrizz[72][613] = 9'b111111111;
assign micromatrizz[72][614] = 9'b111111111;
assign micromatrizz[72][615] = 9'b111111111;
assign micromatrizz[72][616] = 9'b111111111;
assign micromatrizz[72][617] = 9'b111111111;
assign micromatrizz[72][618] = 9'b111111111;
assign micromatrizz[72][619] = 9'b111111111;
assign micromatrizz[72][620] = 9'b111111111;
assign micromatrizz[72][621] = 9'b111111111;
assign micromatrizz[72][622] = 9'b111111111;
assign micromatrizz[72][623] = 9'b111111111;
assign micromatrizz[72][624] = 9'b111111111;
assign micromatrizz[72][625] = 9'b111111111;
assign micromatrizz[72][626] = 9'b111111111;
assign micromatrizz[72][627] = 9'b111111111;
assign micromatrizz[72][628] = 9'b111111111;
assign micromatrizz[72][629] = 9'b111111111;
assign micromatrizz[72][630] = 9'b111111111;
assign micromatrizz[72][631] = 9'b111111111;
assign micromatrizz[72][632] = 9'b111111111;
assign micromatrizz[72][633] = 9'b111111111;
assign micromatrizz[72][634] = 9'b111111111;
assign micromatrizz[72][635] = 9'b111111111;
assign micromatrizz[72][636] = 9'b111111111;
assign micromatrizz[72][637] = 9'b111111111;
assign micromatrizz[72][638] = 9'b111111111;
assign micromatrizz[72][639] = 9'b111111111;
assign micromatrizz[73][0] = 9'b111111111;
assign micromatrizz[73][1] = 9'b111111111;
assign micromatrizz[73][2] = 9'b111111111;
assign micromatrizz[73][3] = 9'b111111111;
assign micromatrizz[73][4] = 9'b111111111;
assign micromatrizz[73][5] = 9'b111111111;
assign micromatrizz[73][6] = 9'b111111111;
assign micromatrizz[73][7] = 9'b111111111;
assign micromatrizz[73][8] = 9'b111111111;
assign micromatrizz[73][9] = 9'b111111111;
assign micromatrizz[73][10] = 9'b111111111;
assign micromatrizz[73][11] = 9'b111111111;
assign micromatrizz[73][12] = 9'b111111111;
assign micromatrizz[73][13] = 9'b111111111;
assign micromatrizz[73][14] = 9'b111111111;
assign micromatrizz[73][15] = 9'b111111111;
assign micromatrizz[73][16] = 9'b111111111;
assign micromatrizz[73][17] = 9'b111111111;
assign micromatrizz[73][18] = 9'b111111111;
assign micromatrizz[73][19] = 9'b111111111;
assign micromatrizz[73][20] = 9'b111111111;
assign micromatrizz[73][21] = 9'b111111111;
assign micromatrizz[73][22] = 9'b111111111;
assign micromatrizz[73][23] = 9'b111111111;
assign micromatrizz[73][24] = 9'b111111111;
assign micromatrizz[73][25] = 9'b111111111;
assign micromatrizz[73][26] = 9'b111111111;
assign micromatrizz[73][27] = 9'b111111111;
assign micromatrizz[73][28] = 9'b111111111;
assign micromatrizz[73][29] = 9'b111111111;
assign micromatrizz[73][30] = 9'b111111111;
assign micromatrizz[73][31] = 9'b111111111;
assign micromatrizz[73][32] = 9'b111111111;
assign micromatrizz[73][33] = 9'b111111111;
assign micromatrizz[73][34] = 9'b111111111;
assign micromatrizz[73][35] = 9'b111111111;
assign micromatrizz[73][36] = 9'b111111111;
assign micromatrizz[73][37] = 9'b111111111;
assign micromatrizz[73][38] = 9'b111111111;
assign micromatrizz[73][39] = 9'b111111111;
assign micromatrizz[73][40] = 9'b111111111;
assign micromatrizz[73][41] = 9'b111111111;
assign micromatrizz[73][42] = 9'b111111111;
assign micromatrizz[73][43] = 9'b111111111;
assign micromatrizz[73][44] = 9'b111111111;
assign micromatrizz[73][45] = 9'b111111111;
assign micromatrizz[73][46] = 9'b111111111;
assign micromatrizz[73][47] = 9'b111111111;
assign micromatrizz[73][48] = 9'b111111111;
assign micromatrizz[73][49] = 9'b111111111;
assign micromatrizz[73][50] = 9'b111111111;
assign micromatrizz[73][51] = 9'b111111111;
assign micromatrizz[73][52] = 9'b111111111;
assign micromatrizz[73][53] = 9'b111111111;
assign micromatrizz[73][54] = 9'b111111111;
assign micromatrizz[73][55] = 9'b111111111;
assign micromatrizz[73][56] = 9'b111111111;
assign micromatrizz[73][57] = 9'b111111111;
assign micromatrizz[73][58] = 9'b111111111;
assign micromatrizz[73][59] = 9'b111111111;
assign micromatrizz[73][60] = 9'b111111111;
assign micromatrizz[73][61] = 9'b111111111;
assign micromatrizz[73][62] = 9'b111111111;
assign micromatrizz[73][63] = 9'b111111111;
assign micromatrizz[73][64] = 9'b111111111;
assign micromatrizz[73][65] = 9'b111111111;
assign micromatrizz[73][66] = 9'b111111111;
assign micromatrizz[73][67] = 9'b111111111;
assign micromatrizz[73][68] = 9'b111111111;
assign micromatrizz[73][69] = 9'b111111111;
assign micromatrizz[73][70] = 9'b111111111;
assign micromatrizz[73][71] = 9'b111111111;
assign micromatrizz[73][72] = 9'b111111111;
assign micromatrizz[73][73] = 9'b111111111;
assign micromatrizz[73][74] = 9'b111111111;
assign micromatrizz[73][75] = 9'b111111111;
assign micromatrizz[73][76] = 9'b111111111;
assign micromatrizz[73][77] = 9'b111111111;
assign micromatrizz[73][78] = 9'b111111111;
assign micromatrizz[73][79] = 9'b111111111;
assign micromatrizz[73][80] = 9'b111111111;
assign micromatrizz[73][81] = 9'b111111111;
assign micromatrizz[73][82] = 9'b111111111;
assign micromatrizz[73][83] = 9'b111111111;
assign micromatrizz[73][84] = 9'b111111111;
assign micromatrizz[73][85] = 9'b111111111;
assign micromatrizz[73][86] = 9'b111111111;
assign micromatrizz[73][87] = 9'b111111111;
assign micromatrizz[73][88] = 9'b111111111;
assign micromatrizz[73][89] = 9'b111111111;
assign micromatrizz[73][90] = 9'b111111111;
assign micromatrizz[73][91] = 9'b111111111;
assign micromatrizz[73][92] = 9'b111111111;
assign micromatrizz[73][93] = 9'b111111111;
assign micromatrizz[73][94] = 9'b111111111;
assign micromatrizz[73][95] = 9'b111111111;
assign micromatrizz[73][96] = 9'b111111111;
assign micromatrizz[73][97] = 9'b111111111;
assign micromatrizz[73][98] = 9'b111111111;
assign micromatrizz[73][99] = 9'b111111111;
assign micromatrizz[73][100] = 9'b111111111;
assign micromatrizz[73][101] = 9'b111111111;
assign micromatrizz[73][102] = 9'b111111111;
assign micromatrizz[73][103] = 9'b111111111;
assign micromatrizz[73][104] = 9'b111111111;
assign micromatrizz[73][105] = 9'b111111111;
assign micromatrizz[73][106] = 9'b111111111;
assign micromatrizz[73][107] = 9'b111111111;
assign micromatrizz[73][108] = 9'b111111111;
assign micromatrizz[73][109] = 9'b111111111;
assign micromatrizz[73][110] = 9'b111111111;
assign micromatrizz[73][111] = 9'b111111111;
assign micromatrizz[73][112] = 9'b111111111;
assign micromatrizz[73][113] = 9'b111111111;
assign micromatrizz[73][114] = 9'b111111111;
assign micromatrizz[73][115] = 9'b111111111;
assign micromatrizz[73][116] = 9'b111111111;
assign micromatrizz[73][117] = 9'b111111111;
assign micromatrizz[73][118] = 9'b111111111;
assign micromatrizz[73][119] = 9'b111111111;
assign micromatrizz[73][120] = 9'b111111111;
assign micromatrizz[73][121] = 9'b111111111;
assign micromatrizz[73][122] = 9'b111111111;
assign micromatrizz[73][123] = 9'b111111111;
assign micromatrizz[73][124] = 9'b111111111;
assign micromatrizz[73][125] = 9'b111111111;
assign micromatrizz[73][126] = 9'b111111111;
assign micromatrizz[73][127] = 9'b111111111;
assign micromatrizz[73][128] = 9'b111111111;
assign micromatrizz[73][129] = 9'b111111111;
assign micromatrizz[73][130] = 9'b111111111;
assign micromatrizz[73][131] = 9'b111111111;
assign micromatrizz[73][132] = 9'b111111111;
assign micromatrizz[73][133] = 9'b111111111;
assign micromatrizz[73][134] = 9'b111111111;
assign micromatrizz[73][135] = 9'b111111111;
assign micromatrizz[73][136] = 9'b111111111;
assign micromatrizz[73][137] = 9'b111111111;
assign micromatrizz[73][138] = 9'b111111111;
assign micromatrizz[73][139] = 9'b111111111;
assign micromatrizz[73][140] = 9'b111111111;
assign micromatrizz[73][141] = 9'b111111111;
assign micromatrizz[73][142] = 9'b111111111;
assign micromatrizz[73][143] = 9'b111111111;
assign micromatrizz[73][144] = 9'b111111111;
assign micromatrizz[73][145] = 9'b111111111;
assign micromatrizz[73][146] = 9'b111111111;
assign micromatrizz[73][147] = 9'b111111111;
assign micromatrizz[73][148] = 9'b111111111;
assign micromatrizz[73][149] = 9'b111111111;
assign micromatrizz[73][150] = 9'b111111111;
assign micromatrizz[73][151] = 9'b111111111;
assign micromatrizz[73][152] = 9'b111111111;
assign micromatrizz[73][153] = 9'b111111111;
assign micromatrizz[73][154] = 9'b111111111;
assign micromatrizz[73][155] = 9'b111111111;
assign micromatrizz[73][156] = 9'b111111111;
assign micromatrizz[73][157] = 9'b111111111;
assign micromatrizz[73][158] = 9'b111111111;
assign micromatrizz[73][159] = 9'b111111111;
assign micromatrizz[73][160] = 9'b111111111;
assign micromatrizz[73][161] = 9'b111111111;
assign micromatrizz[73][162] = 9'b111111111;
assign micromatrizz[73][163] = 9'b111111111;
assign micromatrizz[73][164] = 9'b111111111;
assign micromatrizz[73][165] = 9'b111111111;
assign micromatrizz[73][166] = 9'b111111111;
assign micromatrizz[73][167] = 9'b111111111;
assign micromatrizz[73][168] = 9'b111111111;
assign micromatrizz[73][169] = 9'b111111111;
assign micromatrizz[73][170] = 9'b111111111;
assign micromatrizz[73][171] = 9'b111111111;
assign micromatrizz[73][172] = 9'b111111111;
assign micromatrizz[73][173] = 9'b111111111;
assign micromatrizz[73][174] = 9'b111111111;
assign micromatrizz[73][175] = 9'b111111111;
assign micromatrizz[73][176] = 9'b111111111;
assign micromatrizz[73][177] = 9'b111111111;
assign micromatrizz[73][178] = 9'b111111111;
assign micromatrizz[73][179] = 9'b111111111;
assign micromatrizz[73][180] = 9'b111111111;
assign micromatrizz[73][181] = 9'b111111111;
assign micromatrizz[73][182] = 9'b111111111;
assign micromatrizz[73][183] = 9'b111111111;
assign micromatrizz[73][184] = 9'b111111111;
assign micromatrizz[73][185] = 9'b111111111;
assign micromatrizz[73][186] = 9'b111111111;
assign micromatrizz[73][187] = 9'b111111111;
assign micromatrizz[73][188] = 9'b111111111;
assign micromatrizz[73][189] = 9'b111111111;
assign micromatrizz[73][190] = 9'b111111111;
assign micromatrizz[73][191] = 9'b111111111;
assign micromatrizz[73][192] = 9'b111111111;
assign micromatrizz[73][193] = 9'b111111111;
assign micromatrizz[73][194] = 9'b111111111;
assign micromatrizz[73][195] = 9'b111111111;
assign micromatrizz[73][196] = 9'b111111111;
assign micromatrizz[73][197] = 9'b111111111;
assign micromatrizz[73][198] = 9'b111111111;
assign micromatrizz[73][199] = 9'b111111111;
assign micromatrizz[73][200] = 9'b111111111;
assign micromatrizz[73][201] = 9'b111111111;
assign micromatrizz[73][202] = 9'b111111111;
assign micromatrizz[73][203] = 9'b111111111;
assign micromatrizz[73][204] = 9'b111111111;
assign micromatrizz[73][205] = 9'b111111111;
assign micromatrizz[73][206] = 9'b111111111;
assign micromatrizz[73][207] = 9'b111111111;
assign micromatrizz[73][208] = 9'b111111111;
assign micromatrizz[73][209] = 9'b111111111;
assign micromatrizz[73][210] = 9'b111111111;
assign micromatrizz[73][211] = 9'b111111111;
assign micromatrizz[73][212] = 9'b111111111;
assign micromatrizz[73][213] = 9'b111111111;
assign micromatrizz[73][214] = 9'b111111111;
assign micromatrizz[73][215] = 9'b111111111;
assign micromatrizz[73][216] = 9'b111111111;
assign micromatrizz[73][217] = 9'b111111111;
assign micromatrizz[73][218] = 9'b111111111;
assign micromatrizz[73][219] = 9'b111111111;
assign micromatrizz[73][220] = 9'b111111111;
assign micromatrizz[73][221] = 9'b111111111;
assign micromatrizz[73][222] = 9'b111111111;
assign micromatrizz[73][223] = 9'b111111111;
assign micromatrizz[73][224] = 9'b111111111;
assign micromatrizz[73][225] = 9'b111111111;
assign micromatrizz[73][226] = 9'b111111111;
assign micromatrizz[73][227] = 9'b111111111;
assign micromatrizz[73][228] = 9'b111111111;
assign micromatrizz[73][229] = 9'b111111111;
assign micromatrizz[73][230] = 9'b111111111;
assign micromatrizz[73][231] = 9'b111111111;
assign micromatrizz[73][232] = 9'b111111111;
assign micromatrizz[73][233] = 9'b111111111;
assign micromatrizz[73][234] = 9'b111111111;
assign micromatrizz[73][235] = 9'b111111111;
assign micromatrizz[73][236] = 9'b111111111;
assign micromatrizz[73][237] = 9'b111111111;
assign micromatrizz[73][238] = 9'b111111111;
assign micromatrizz[73][239] = 9'b111111111;
assign micromatrizz[73][240] = 9'b111111111;
assign micromatrizz[73][241] = 9'b111111111;
assign micromatrizz[73][242] = 9'b111111111;
assign micromatrizz[73][243] = 9'b111111111;
assign micromatrizz[73][244] = 9'b111111111;
assign micromatrizz[73][245] = 9'b111111111;
assign micromatrizz[73][246] = 9'b111111111;
assign micromatrizz[73][247] = 9'b111111111;
assign micromatrizz[73][248] = 9'b111111111;
assign micromatrizz[73][249] = 9'b111111111;
assign micromatrizz[73][250] = 9'b111111111;
assign micromatrizz[73][251] = 9'b111111111;
assign micromatrizz[73][252] = 9'b111111111;
assign micromatrizz[73][253] = 9'b111111111;
assign micromatrizz[73][254] = 9'b111111111;
assign micromatrizz[73][255] = 9'b111111111;
assign micromatrizz[73][256] = 9'b111111111;
assign micromatrizz[73][257] = 9'b111111111;
assign micromatrizz[73][258] = 9'b111111111;
assign micromatrizz[73][259] = 9'b111111111;
assign micromatrizz[73][260] = 9'b111111111;
assign micromatrizz[73][261] = 9'b111111111;
assign micromatrizz[73][262] = 9'b111111111;
assign micromatrizz[73][263] = 9'b111111111;
assign micromatrizz[73][264] = 9'b111111111;
assign micromatrizz[73][265] = 9'b111111111;
assign micromatrizz[73][266] = 9'b111111111;
assign micromatrizz[73][267] = 9'b111111111;
assign micromatrizz[73][268] = 9'b111111111;
assign micromatrizz[73][269] = 9'b111111111;
assign micromatrizz[73][270] = 9'b111111111;
assign micromatrizz[73][271] = 9'b111111111;
assign micromatrizz[73][272] = 9'b111111111;
assign micromatrizz[73][273] = 9'b111111111;
assign micromatrizz[73][274] = 9'b111111111;
assign micromatrizz[73][275] = 9'b111111111;
assign micromatrizz[73][276] = 9'b111111111;
assign micromatrizz[73][277] = 9'b111111111;
assign micromatrizz[73][278] = 9'b111111111;
assign micromatrizz[73][279] = 9'b111111111;
assign micromatrizz[73][280] = 9'b111111111;
assign micromatrizz[73][281] = 9'b111111111;
assign micromatrizz[73][282] = 9'b111111111;
assign micromatrizz[73][283] = 9'b111111111;
assign micromatrizz[73][284] = 9'b111111111;
assign micromatrizz[73][285] = 9'b111111111;
assign micromatrizz[73][286] = 9'b111111111;
assign micromatrizz[73][287] = 9'b111111111;
assign micromatrizz[73][288] = 9'b111111111;
assign micromatrizz[73][289] = 9'b111111111;
assign micromatrizz[73][290] = 9'b111111111;
assign micromatrizz[73][291] = 9'b111111111;
assign micromatrizz[73][292] = 9'b111111111;
assign micromatrizz[73][293] = 9'b111111111;
assign micromatrizz[73][294] = 9'b111111111;
assign micromatrizz[73][295] = 9'b111111111;
assign micromatrizz[73][296] = 9'b111111111;
assign micromatrizz[73][297] = 9'b111111111;
assign micromatrizz[73][298] = 9'b111111111;
assign micromatrizz[73][299] = 9'b111111111;
assign micromatrizz[73][300] = 9'b111111111;
assign micromatrizz[73][301] = 9'b111111111;
assign micromatrizz[73][302] = 9'b111111111;
assign micromatrizz[73][303] = 9'b111111111;
assign micromatrizz[73][304] = 9'b111111111;
assign micromatrizz[73][305] = 9'b111111111;
assign micromatrizz[73][306] = 9'b111111111;
assign micromatrizz[73][307] = 9'b111111111;
assign micromatrizz[73][308] = 9'b111111111;
assign micromatrizz[73][309] = 9'b111111111;
assign micromatrizz[73][310] = 9'b111111111;
assign micromatrizz[73][311] = 9'b111111111;
assign micromatrizz[73][312] = 9'b111111111;
assign micromatrizz[73][313] = 9'b111111111;
assign micromatrizz[73][314] = 9'b111111111;
assign micromatrizz[73][315] = 9'b111111111;
assign micromatrizz[73][316] = 9'b111111111;
assign micromatrizz[73][317] = 9'b111111111;
assign micromatrizz[73][318] = 9'b111111111;
assign micromatrizz[73][319] = 9'b111111111;
assign micromatrizz[73][320] = 9'b111111111;
assign micromatrizz[73][321] = 9'b111111111;
assign micromatrizz[73][322] = 9'b111111111;
assign micromatrizz[73][323] = 9'b111111111;
assign micromatrizz[73][324] = 9'b111111111;
assign micromatrizz[73][325] = 9'b111111111;
assign micromatrizz[73][326] = 9'b111111111;
assign micromatrizz[73][327] = 9'b111111111;
assign micromatrizz[73][328] = 9'b111111111;
assign micromatrizz[73][329] = 9'b111111111;
assign micromatrizz[73][330] = 9'b111111111;
assign micromatrizz[73][331] = 9'b111111111;
assign micromatrizz[73][332] = 9'b111111111;
assign micromatrizz[73][333] = 9'b111111111;
assign micromatrizz[73][334] = 9'b111111111;
assign micromatrizz[73][335] = 9'b111111111;
assign micromatrizz[73][336] = 9'b111111111;
assign micromatrizz[73][337] = 9'b111111111;
assign micromatrizz[73][338] = 9'b111111111;
assign micromatrizz[73][339] = 9'b111111111;
assign micromatrizz[73][340] = 9'b111111111;
assign micromatrizz[73][341] = 9'b111111111;
assign micromatrizz[73][342] = 9'b111111111;
assign micromatrizz[73][343] = 9'b111111111;
assign micromatrizz[73][344] = 9'b111111111;
assign micromatrizz[73][345] = 9'b111111111;
assign micromatrizz[73][346] = 9'b111111111;
assign micromatrizz[73][347] = 9'b111111111;
assign micromatrizz[73][348] = 9'b111111111;
assign micromatrizz[73][349] = 9'b111111111;
assign micromatrizz[73][350] = 9'b111111111;
assign micromatrizz[73][351] = 9'b111111111;
assign micromatrizz[73][352] = 9'b111111111;
assign micromatrizz[73][353] = 9'b111111111;
assign micromatrizz[73][354] = 9'b111111111;
assign micromatrizz[73][355] = 9'b111111111;
assign micromatrizz[73][356] = 9'b111111111;
assign micromatrizz[73][357] = 9'b111111111;
assign micromatrizz[73][358] = 9'b111111111;
assign micromatrizz[73][359] = 9'b111111111;
assign micromatrizz[73][360] = 9'b111111111;
assign micromatrizz[73][361] = 9'b111111111;
assign micromatrizz[73][362] = 9'b111111111;
assign micromatrizz[73][363] = 9'b111111111;
assign micromatrizz[73][364] = 9'b111111111;
assign micromatrizz[73][365] = 9'b111111111;
assign micromatrizz[73][366] = 9'b111111111;
assign micromatrizz[73][367] = 9'b111111111;
assign micromatrizz[73][368] = 9'b111111111;
assign micromatrizz[73][369] = 9'b111111111;
assign micromatrizz[73][370] = 9'b111111111;
assign micromatrizz[73][371] = 9'b111111111;
assign micromatrizz[73][372] = 9'b111111111;
assign micromatrizz[73][373] = 9'b111111111;
assign micromatrizz[73][374] = 9'b111111111;
assign micromatrizz[73][375] = 9'b111111111;
assign micromatrizz[73][376] = 9'b111111111;
assign micromatrizz[73][377] = 9'b111111111;
assign micromatrizz[73][378] = 9'b111111111;
assign micromatrizz[73][379] = 9'b111111111;
assign micromatrizz[73][380] = 9'b111111111;
assign micromatrizz[73][381] = 9'b111111111;
assign micromatrizz[73][382] = 9'b111111111;
assign micromatrizz[73][383] = 9'b111111111;
assign micromatrizz[73][384] = 9'b111111111;
assign micromatrizz[73][385] = 9'b111111111;
assign micromatrizz[73][386] = 9'b111111111;
assign micromatrizz[73][387] = 9'b111111111;
assign micromatrizz[73][388] = 9'b111111111;
assign micromatrizz[73][389] = 9'b111111111;
assign micromatrizz[73][390] = 9'b111111111;
assign micromatrizz[73][391] = 9'b111111111;
assign micromatrizz[73][392] = 9'b111111111;
assign micromatrizz[73][393] = 9'b111111111;
assign micromatrizz[73][394] = 9'b111111111;
assign micromatrizz[73][395] = 9'b111111111;
assign micromatrizz[73][396] = 9'b111111111;
assign micromatrizz[73][397] = 9'b111111111;
assign micromatrizz[73][398] = 9'b111111111;
assign micromatrizz[73][399] = 9'b111111111;
assign micromatrizz[73][400] = 9'b111111111;
assign micromatrizz[73][401] = 9'b111111111;
assign micromatrizz[73][402] = 9'b111111111;
assign micromatrizz[73][403] = 9'b111111111;
assign micromatrizz[73][404] = 9'b111111111;
assign micromatrizz[73][405] = 9'b111111111;
assign micromatrizz[73][406] = 9'b111111111;
assign micromatrizz[73][407] = 9'b111111111;
assign micromatrizz[73][408] = 9'b111111111;
assign micromatrizz[73][409] = 9'b111111111;
assign micromatrizz[73][410] = 9'b111111111;
assign micromatrizz[73][411] = 9'b111111111;
assign micromatrizz[73][412] = 9'b111111111;
assign micromatrizz[73][413] = 9'b111111111;
assign micromatrizz[73][414] = 9'b111111111;
assign micromatrizz[73][415] = 9'b111111111;
assign micromatrizz[73][416] = 9'b111111111;
assign micromatrizz[73][417] = 9'b111111111;
assign micromatrizz[73][418] = 9'b111111111;
assign micromatrizz[73][419] = 9'b111111111;
assign micromatrizz[73][420] = 9'b111111111;
assign micromatrizz[73][421] = 9'b111111111;
assign micromatrizz[73][422] = 9'b111111111;
assign micromatrizz[73][423] = 9'b111111111;
assign micromatrizz[73][424] = 9'b111111111;
assign micromatrizz[73][425] = 9'b111111111;
assign micromatrizz[73][426] = 9'b111111111;
assign micromatrizz[73][427] = 9'b111111111;
assign micromatrizz[73][428] = 9'b111111111;
assign micromatrizz[73][429] = 9'b111111111;
assign micromatrizz[73][430] = 9'b111111111;
assign micromatrizz[73][431] = 9'b111111111;
assign micromatrizz[73][432] = 9'b111111111;
assign micromatrizz[73][433] = 9'b111111111;
assign micromatrizz[73][434] = 9'b111111111;
assign micromatrizz[73][435] = 9'b111111111;
assign micromatrizz[73][436] = 9'b111111111;
assign micromatrizz[73][437] = 9'b111111111;
assign micromatrizz[73][438] = 9'b111111111;
assign micromatrizz[73][439] = 9'b111111111;
assign micromatrizz[73][440] = 9'b111111111;
assign micromatrizz[73][441] = 9'b111111111;
assign micromatrizz[73][442] = 9'b111111111;
assign micromatrizz[73][443] = 9'b111111111;
assign micromatrizz[73][444] = 9'b111111111;
assign micromatrizz[73][445] = 9'b111111111;
assign micromatrizz[73][446] = 9'b111111111;
assign micromatrizz[73][447] = 9'b111111111;
assign micromatrizz[73][448] = 9'b111111111;
assign micromatrizz[73][449] = 9'b111111111;
assign micromatrizz[73][450] = 9'b111111111;
assign micromatrizz[73][451] = 9'b111111111;
assign micromatrizz[73][452] = 9'b111111111;
assign micromatrizz[73][453] = 9'b111111111;
assign micromatrizz[73][454] = 9'b111111111;
assign micromatrizz[73][455] = 9'b111111111;
assign micromatrizz[73][456] = 9'b111111111;
assign micromatrizz[73][457] = 9'b111111111;
assign micromatrizz[73][458] = 9'b111111111;
assign micromatrizz[73][459] = 9'b111111111;
assign micromatrizz[73][460] = 9'b111111111;
assign micromatrizz[73][461] = 9'b111111111;
assign micromatrizz[73][462] = 9'b111111111;
assign micromatrizz[73][463] = 9'b111111111;
assign micromatrizz[73][464] = 9'b111111111;
assign micromatrizz[73][465] = 9'b111111111;
assign micromatrizz[73][466] = 9'b111111111;
assign micromatrizz[73][467] = 9'b111111111;
assign micromatrizz[73][468] = 9'b111111111;
assign micromatrizz[73][469] = 9'b111111111;
assign micromatrizz[73][470] = 9'b111111111;
assign micromatrizz[73][471] = 9'b111111111;
assign micromatrizz[73][472] = 9'b111111111;
assign micromatrizz[73][473] = 9'b111111111;
assign micromatrizz[73][474] = 9'b111111111;
assign micromatrizz[73][475] = 9'b111111111;
assign micromatrizz[73][476] = 9'b111111111;
assign micromatrizz[73][477] = 9'b111111111;
assign micromatrizz[73][478] = 9'b111111111;
assign micromatrizz[73][479] = 9'b111111111;
assign micromatrizz[73][480] = 9'b111111111;
assign micromatrizz[73][481] = 9'b111111111;
assign micromatrizz[73][482] = 9'b111111111;
assign micromatrizz[73][483] = 9'b111111111;
assign micromatrizz[73][484] = 9'b111111111;
assign micromatrizz[73][485] = 9'b111111111;
assign micromatrizz[73][486] = 9'b111111111;
assign micromatrizz[73][487] = 9'b111111111;
assign micromatrizz[73][488] = 9'b111111111;
assign micromatrizz[73][489] = 9'b111111111;
assign micromatrizz[73][490] = 9'b111111111;
assign micromatrizz[73][491] = 9'b111111111;
assign micromatrizz[73][492] = 9'b111111111;
assign micromatrizz[73][493] = 9'b111111111;
assign micromatrizz[73][494] = 9'b111111111;
assign micromatrizz[73][495] = 9'b111111111;
assign micromatrizz[73][496] = 9'b111111111;
assign micromatrizz[73][497] = 9'b111111111;
assign micromatrizz[73][498] = 9'b111111111;
assign micromatrizz[73][499] = 9'b111111111;
assign micromatrizz[73][500] = 9'b111111111;
assign micromatrizz[73][501] = 9'b111111111;
assign micromatrizz[73][502] = 9'b111111111;
assign micromatrizz[73][503] = 9'b111111111;
assign micromatrizz[73][504] = 9'b111111111;
assign micromatrizz[73][505] = 9'b111111111;
assign micromatrizz[73][506] = 9'b111111111;
assign micromatrizz[73][507] = 9'b111111111;
assign micromatrizz[73][508] = 9'b111111111;
assign micromatrizz[73][509] = 9'b111111111;
assign micromatrizz[73][510] = 9'b111111111;
assign micromatrizz[73][511] = 9'b111111111;
assign micromatrizz[73][512] = 9'b111111111;
assign micromatrizz[73][513] = 9'b111111111;
assign micromatrizz[73][514] = 9'b111111111;
assign micromatrizz[73][515] = 9'b111111111;
assign micromatrizz[73][516] = 9'b111111111;
assign micromatrizz[73][517] = 9'b111111111;
assign micromatrizz[73][518] = 9'b111111111;
assign micromatrizz[73][519] = 9'b111111111;
assign micromatrizz[73][520] = 9'b111111111;
assign micromatrizz[73][521] = 9'b111111111;
assign micromatrizz[73][522] = 9'b111111111;
assign micromatrizz[73][523] = 9'b111111111;
assign micromatrizz[73][524] = 9'b111111111;
assign micromatrizz[73][525] = 9'b111111111;
assign micromatrizz[73][526] = 9'b111111111;
assign micromatrizz[73][527] = 9'b111111111;
assign micromatrizz[73][528] = 9'b111111111;
assign micromatrizz[73][529] = 9'b111111111;
assign micromatrizz[73][530] = 9'b111111111;
assign micromatrizz[73][531] = 9'b111111111;
assign micromatrizz[73][532] = 9'b111111111;
assign micromatrizz[73][533] = 9'b111111111;
assign micromatrizz[73][534] = 9'b111111111;
assign micromatrizz[73][535] = 9'b111111111;
assign micromatrizz[73][536] = 9'b111111111;
assign micromatrizz[73][537] = 9'b111111111;
assign micromatrizz[73][538] = 9'b111111111;
assign micromatrizz[73][539] = 9'b111111111;
assign micromatrizz[73][540] = 9'b111111111;
assign micromatrizz[73][541] = 9'b111111111;
assign micromatrizz[73][542] = 9'b111111111;
assign micromatrizz[73][543] = 9'b111111111;
assign micromatrizz[73][544] = 9'b111111111;
assign micromatrizz[73][545] = 9'b111111111;
assign micromatrizz[73][546] = 9'b111111111;
assign micromatrizz[73][547] = 9'b111111111;
assign micromatrizz[73][548] = 9'b111111111;
assign micromatrizz[73][549] = 9'b111111111;
assign micromatrizz[73][550] = 9'b111111111;
assign micromatrizz[73][551] = 9'b111111111;
assign micromatrizz[73][552] = 9'b111111111;
assign micromatrizz[73][553] = 9'b111111111;
assign micromatrizz[73][554] = 9'b111111111;
assign micromatrizz[73][555] = 9'b111111111;
assign micromatrizz[73][556] = 9'b111111111;
assign micromatrizz[73][557] = 9'b111111111;
assign micromatrizz[73][558] = 9'b111111111;
assign micromatrizz[73][559] = 9'b111111111;
assign micromatrizz[73][560] = 9'b111111111;
assign micromatrizz[73][561] = 9'b111111111;
assign micromatrizz[73][562] = 9'b111111111;
assign micromatrizz[73][563] = 9'b111111111;
assign micromatrizz[73][564] = 9'b111111111;
assign micromatrizz[73][565] = 9'b111111111;
assign micromatrizz[73][566] = 9'b111111111;
assign micromatrizz[73][567] = 9'b111111111;
assign micromatrizz[73][568] = 9'b111111111;
assign micromatrizz[73][569] = 9'b111111111;
assign micromatrizz[73][570] = 9'b111111111;
assign micromatrizz[73][571] = 9'b111111111;
assign micromatrizz[73][572] = 9'b111111111;
assign micromatrizz[73][573] = 9'b111111111;
assign micromatrizz[73][574] = 9'b111111111;
assign micromatrizz[73][575] = 9'b111111111;
assign micromatrizz[73][576] = 9'b111111111;
assign micromatrizz[73][577] = 9'b111111111;
assign micromatrizz[73][578] = 9'b111111111;
assign micromatrizz[73][579] = 9'b111111111;
assign micromatrizz[73][580] = 9'b111111111;
assign micromatrizz[73][581] = 9'b111111111;
assign micromatrizz[73][582] = 9'b111111111;
assign micromatrizz[73][583] = 9'b111111111;
assign micromatrizz[73][584] = 9'b111111111;
assign micromatrizz[73][585] = 9'b111111111;
assign micromatrizz[73][586] = 9'b111111111;
assign micromatrizz[73][587] = 9'b111111111;
assign micromatrizz[73][588] = 9'b111111111;
assign micromatrizz[73][589] = 9'b111111111;
assign micromatrizz[73][590] = 9'b111111111;
assign micromatrizz[73][591] = 9'b111111111;
assign micromatrizz[73][592] = 9'b111111111;
assign micromatrizz[73][593] = 9'b111111111;
assign micromatrizz[73][594] = 9'b111111111;
assign micromatrizz[73][595] = 9'b111111111;
assign micromatrizz[73][596] = 9'b111111111;
assign micromatrizz[73][597] = 9'b111111111;
assign micromatrizz[73][598] = 9'b111111111;
assign micromatrizz[73][599] = 9'b111111111;
assign micromatrizz[73][600] = 9'b111111111;
assign micromatrizz[73][601] = 9'b111111111;
assign micromatrizz[73][602] = 9'b111111111;
assign micromatrizz[73][603] = 9'b111111111;
assign micromatrizz[73][604] = 9'b111111111;
assign micromatrizz[73][605] = 9'b111111111;
assign micromatrizz[73][606] = 9'b111111111;
assign micromatrizz[73][607] = 9'b111111111;
assign micromatrizz[73][608] = 9'b111111111;
assign micromatrizz[73][609] = 9'b111111111;
assign micromatrizz[73][610] = 9'b111111111;
assign micromatrizz[73][611] = 9'b111111111;
assign micromatrizz[73][612] = 9'b111111111;
assign micromatrizz[73][613] = 9'b111111111;
assign micromatrizz[73][614] = 9'b111111111;
assign micromatrizz[73][615] = 9'b111111111;
assign micromatrizz[73][616] = 9'b111111111;
assign micromatrizz[73][617] = 9'b111111111;
assign micromatrizz[73][618] = 9'b111111111;
assign micromatrizz[73][619] = 9'b111111111;
assign micromatrizz[73][620] = 9'b111111111;
assign micromatrizz[73][621] = 9'b111111111;
assign micromatrizz[73][622] = 9'b111111111;
assign micromatrizz[73][623] = 9'b111111111;
assign micromatrizz[73][624] = 9'b111111111;
assign micromatrizz[73][625] = 9'b111111111;
assign micromatrizz[73][626] = 9'b111111111;
assign micromatrizz[73][627] = 9'b111111111;
assign micromatrizz[73][628] = 9'b111111111;
assign micromatrizz[73][629] = 9'b111111111;
assign micromatrizz[73][630] = 9'b111111111;
assign micromatrizz[73][631] = 9'b111111111;
assign micromatrizz[73][632] = 9'b111111111;
assign micromatrizz[73][633] = 9'b111111111;
assign micromatrizz[73][634] = 9'b111111111;
assign micromatrizz[73][635] = 9'b111111111;
assign micromatrizz[73][636] = 9'b111111111;
assign micromatrizz[73][637] = 9'b111111111;
assign micromatrizz[73][638] = 9'b111111111;
assign micromatrizz[73][639] = 9'b111111111;
assign micromatrizz[74][0] = 9'b111111111;
assign micromatrizz[74][1] = 9'b111111111;
assign micromatrizz[74][2] = 9'b111111111;
assign micromatrizz[74][3] = 9'b111111111;
assign micromatrizz[74][4] = 9'b111111111;
assign micromatrizz[74][5] = 9'b111111111;
assign micromatrizz[74][6] = 9'b111111111;
assign micromatrizz[74][7] = 9'b111111111;
assign micromatrizz[74][8] = 9'b111111111;
assign micromatrizz[74][9] = 9'b111111111;
assign micromatrizz[74][10] = 9'b111111111;
assign micromatrizz[74][11] = 9'b111111111;
assign micromatrizz[74][12] = 9'b111111111;
assign micromatrizz[74][13] = 9'b111111111;
assign micromatrizz[74][14] = 9'b111111111;
assign micromatrizz[74][15] = 9'b111111111;
assign micromatrizz[74][16] = 9'b111111111;
assign micromatrizz[74][17] = 9'b111111111;
assign micromatrizz[74][18] = 9'b111111111;
assign micromatrizz[74][19] = 9'b111111111;
assign micromatrizz[74][20] = 9'b111111111;
assign micromatrizz[74][21] = 9'b111111111;
assign micromatrizz[74][22] = 9'b111111111;
assign micromatrizz[74][23] = 9'b111111111;
assign micromatrizz[74][24] = 9'b111111111;
assign micromatrizz[74][25] = 9'b111111111;
assign micromatrizz[74][26] = 9'b111111111;
assign micromatrizz[74][27] = 9'b111111111;
assign micromatrizz[74][28] = 9'b111111111;
assign micromatrizz[74][29] = 9'b111111111;
assign micromatrizz[74][30] = 9'b111111111;
assign micromatrizz[74][31] = 9'b111111111;
assign micromatrizz[74][32] = 9'b111111111;
assign micromatrizz[74][33] = 9'b111111111;
assign micromatrizz[74][34] = 9'b111111111;
assign micromatrizz[74][35] = 9'b111111111;
assign micromatrizz[74][36] = 9'b111111111;
assign micromatrizz[74][37] = 9'b111111111;
assign micromatrizz[74][38] = 9'b111111111;
assign micromatrizz[74][39] = 9'b111111111;
assign micromatrizz[74][40] = 9'b111111111;
assign micromatrizz[74][41] = 9'b111111111;
assign micromatrizz[74][42] = 9'b111111111;
assign micromatrizz[74][43] = 9'b111111111;
assign micromatrizz[74][44] = 9'b111111111;
assign micromatrizz[74][45] = 9'b111111111;
assign micromatrizz[74][46] = 9'b111111111;
assign micromatrizz[74][47] = 9'b111111111;
assign micromatrizz[74][48] = 9'b111111111;
assign micromatrizz[74][49] = 9'b111111111;
assign micromatrizz[74][50] = 9'b111111111;
assign micromatrizz[74][51] = 9'b111111111;
assign micromatrizz[74][52] = 9'b111111111;
assign micromatrizz[74][53] = 9'b111111111;
assign micromatrizz[74][54] = 9'b111111111;
assign micromatrizz[74][55] = 9'b111111111;
assign micromatrizz[74][56] = 9'b111111111;
assign micromatrizz[74][57] = 9'b111111111;
assign micromatrizz[74][58] = 9'b111111111;
assign micromatrizz[74][59] = 9'b111111111;
assign micromatrizz[74][60] = 9'b111111111;
assign micromatrizz[74][61] = 9'b111111111;
assign micromatrizz[74][62] = 9'b111111111;
assign micromatrizz[74][63] = 9'b111111111;
assign micromatrizz[74][64] = 9'b111111111;
assign micromatrizz[74][65] = 9'b111111111;
assign micromatrizz[74][66] = 9'b111111111;
assign micromatrizz[74][67] = 9'b111111111;
assign micromatrizz[74][68] = 9'b111111111;
assign micromatrizz[74][69] = 9'b111111111;
assign micromatrizz[74][70] = 9'b111111111;
assign micromatrizz[74][71] = 9'b111111111;
assign micromatrizz[74][72] = 9'b111111111;
assign micromatrizz[74][73] = 9'b111111111;
assign micromatrizz[74][74] = 9'b111111111;
assign micromatrizz[74][75] = 9'b111111111;
assign micromatrizz[74][76] = 9'b111111111;
assign micromatrizz[74][77] = 9'b111111111;
assign micromatrizz[74][78] = 9'b111111111;
assign micromatrizz[74][79] = 9'b111111111;
assign micromatrizz[74][80] = 9'b111111111;
assign micromatrizz[74][81] = 9'b111111111;
assign micromatrizz[74][82] = 9'b111111111;
assign micromatrizz[74][83] = 9'b111111111;
assign micromatrizz[74][84] = 9'b111111111;
assign micromatrizz[74][85] = 9'b111111111;
assign micromatrizz[74][86] = 9'b111111111;
assign micromatrizz[74][87] = 9'b111111111;
assign micromatrizz[74][88] = 9'b111111111;
assign micromatrizz[74][89] = 9'b111111111;
assign micromatrizz[74][90] = 9'b111111111;
assign micromatrizz[74][91] = 9'b111111111;
assign micromatrizz[74][92] = 9'b111111111;
assign micromatrizz[74][93] = 9'b111111111;
assign micromatrizz[74][94] = 9'b111111111;
assign micromatrizz[74][95] = 9'b111111111;
assign micromatrizz[74][96] = 9'b111111111;
assign micromatrizz[74][97] = 9'b111111111;
assign micromatrizz[74][98] = 9'b111111111;
assign micromatrizz[74][99] = 9'b111111111;
assign micromatrizz[74][100] = 9'b111111111;
assign micromatrizz[74][101] = 9'b111111111;
assign micromatrizz[74][102] = 9'b111111111;
assign micromatrizz[74][103] = 9'b111111111;
assign micromatrizz[74][104] = 9'b111111111;
assign micromatrizz[74][105] = 9'b111111111;
assign micromatrizz[74][106] = 9'b111111111;
assign micromatrizz[74][107] = 9'b111111111;
assign micromatrizz[74][108] = 9'b111111111;
assign micromatrizz[74][109] = 9'b111111111;
assign micromatrizz[74][110] = 9'b111111111;
assign micromatrizz[74][111] = 9'b111111111;
assign micromatrizz[74][112] = 9'b111111111;
assign micromatrizz[74][113] = 9'b111111111;
assign micromatrizz[74][114] = 9'b111111111;
assign micromatrizz[74][115] = 9'b111111111;
assign micromatrizz[74][116] = 9'b111111111;
assign micromatrizz[74][117] = 9'b111111111;
assign micromatrizz[74][118] = 9'b111111111;
assign micromatrizz[74][119] = 9'b111111111;
assign micromatrizz[74][120] = 9'b111111111;
assign micromatrizz[74][121] = 9'b111111111;
assign micromatrizz[74][122] = 9'b111111111;
assign micromatrizz[74][123] = 9'b111111111;
assign micromatrizz[74][124] = 9'b111111111;
assign micromatrizz[74][125] = 9'b111111111;
assign micromatrizz[74][126] = 9'b111111111;
assign micromatrizz[74][127] = 9'b111111111;
assign micromatrizz[74][128] = 9'b111111111;
assign micromatrizz[74][129] = 9'b111111111;
assign micromatrizz[74][130] = 9'b111111111;
assign micromatrizz[74][131] = 9'b111111111;
assign micromatrizz[74][132] = 9'b111111111;
assign micromatrizz[74][133] = 9'b111111111;
assign micromatrizz[74][134] = 9'b111111111;
assign micromatrizz[74][135] = 9'b111111111;
assign micromatrizz[74][136] = 9'b111111111;
assign micromatrizz[74][137] = 9'b111111111;
assign micromatrizz[74][138] = 9'b111111111;
assign micromatrizz[74][139] = 9'b111111111;
assign micromatrizz[74][140] = 9'b111111111;
assign micromatrizz[74][141] = 9'b111111111;
assign micromatrizz[74][142] = 9'b111111111;
assign micromatrizz[74][143] = 9'b111111111;
assign micromatrizz[74][144] = 9'b111111111;
assign micromatrizz[74][145] = 9'b111111111;
assign micromatrizz[74][146] = 9'b111111111;
assign micromatrizz[74][147] = 9'b111111111;
assign micromatrizz[74][148] = 9'b111111111;
assign micromatrizz[74][149] = 9'b111111111;
assign micromatrizz[74][150] = 9'b111111111;
assign micromatrizz[74][151] = 9'b111111111;
assign micromatrizz[74][152] = 9'b111111111;
assign micromatrizz[74][153] = 9'b111111111;
assign micromatrizz[74][154] = 9'b111111111;
assign micromatrizz[74][155] = 9'b111111111;
assign micromatrizz[74][156] = 9'b111111111;
assign micromatrizz[74][157] = 9'b111111111;
assign micromatrizz[74][158] = 9'b111111111;
assign micromatrizz[74][159] = 9'b111111111;
assign micromatrizz[74][160] = 9'b111111111;
assign micromatrizz[74][161] = 9'b111111111;
assign micromatrizz[74][162] = 9'b111111111;
assign micromatrizz[74][163] = 9'b111111111;
assign micromatrizz[74][164] = 9'b111111111;
assign micromatrizz[74][165] = 9'b111111111;
assign micromatrizz[74][166] = 9'b111111111;
assign micromatrizz[74][167] = 9'b111111111;
assign micromatrizz[74][168] = 9'b111111111;
assign micromatrizz[74][169] = 9'b111111111;
assign micromatrizz[74][170] = 9'b111111111;
assign micromatrizz[74][171] = 9'b111111111;
assign micromatrizz[74][172] = 9'b111111111;
assign micromatrizz[74][173] = 9'b111111111;
assign micromatrizz[74][174] = 9'b111111111;
assign micromatrizz[74][175] = 9'b111111111;
assign micromatrizz[74][176] = 9'b111111111;
assign micromatrizz[74][177] = 9'b111111111;
assign micromatrizz[74][178] = 9'b111111111;
assign micromatrizz[74][179] = 9'b111111111;
assign micromatrizz[74][180] = 9'b111111111;
assign micromatrizz[74][181] = 9'b111111111;
assign micromatrizz[74][182] = 9'b111111111;
assign micromatrizz[74][183] = 9'b111111111;
assign micromatrizz[74][184] = 9'b111111111;
assign micromatrizz[74][185] = 9'b111111111;
assign micromatrizz[74][186] = 9'b111111111;
assign micromatrizz[74][187] = 9'b111111111;
assign micromatrizz[74][188] = 9'b111111111;
assign micromatrizz[74][189] = 9'b111111111;
assign micromatrizz[74][190] = 9'b111111111;
assign micromatrizz[74][191] = 9'b111111111;
assign micromatrizz[74][192] = 9'b111111111;
assign micromatrizz[74][193] = 9'b111111111;
assign micromatrizz[74][194] = 9'b111111111;
assign micromatrizz[74][195] = 9'b111111111;
assign micromatrizz[74][196] = 9'b111111111;
assign micromatrizz[74][197] = 9'b111111111;
assign micromatrizz[74][198] = 9'b111111111;
assign micromatrizz[74][199] = 9'b111111111;
assign micromatrizz[74][200] = 9'b111111111;
assign micromatrizz[74][201] = 9'b111111111;
assign micromatrizz[74][202] = 9'b111111111;
assign micromatrizz[74][203] = 9'b111111111;
assign micromatrizz[74][204] = 9'b111111111;
assign micromatrizz[74][205] = 9'b111111111;
assign micromatrizz[74][206] = 9'b111111111;
assign micromatrizz[74][207] = 9'b111111111;
assign micromatrizz[74][208] = 9'b111111111;
assign micromatrizz[74][209] = 9'b111111111;
assign micromatrizz[74][210] = 9'b111111111;
assign micromatrizz[74][211] = 9'b111111111;
assign micromatrizz[74][212] = 9'b111111111;
assign micromatrizz[74][213] = 9'b111111111;
assign micromatrizz[74][214] = 9'b111111111;
assign micromatrizz[74][215] = 9'b111111111;
assign micromatrizz[74][216] = 9'b111111111;
assign micromatrizz[74][217] = 9'b111111111;
assign micromatrizz[74][218] = 9'b111111111;
assign micromatrizz[74][219] = 9'b111111111;
assign micromatrizz[74][220] = 9'b111111111;
assign micromatrizz[74][221] = 9'b111111111;
assign micromatrizz[74][222] = 9'b111111111;
assign micromatrizz[74][223] = 9'b111111111;
assign micromatrizz[74][224] = 9'b111111111;
assign micromatrizz[74][225] = 9'b111111111;
assign micromatrizz[74][226] = 9'b111111111;
assign micromatrizz[74][227] = 9'b111111111;
assign micromatrizz[74][228] = 9'b111111111;
assign micromatrizz[74][229] = 9'b111111111;
assign micromatrizz[74][230] = 9'b111111111;
assign micromatrizz[74][231] = 9'b111111111;
assign micromatrizz[74][232] = 9'b111111111;
assign micromatrizz[74][233] = 9'b111111111;
assign micromatrizz[74][234] = 9'b111111111;
assign micromatrizz[74][235] = 9'b111111111;
assign micromatrizz[74][236] = 9'b111111111;
assign micromatrizz[74][237] = 9'b111111111;
assign micromatrizz[74][238] = 9'b111111111;
assign micromatrizz[74][239] = 9'b111111111;
assign micromatrizz[74][240] = 9'b111111111;
assign micromatrizz[74][241] = 9'b111111111;
assign micromatrizz[74][242] = 9'b111111111;
assign micromatrizz[74][243] = 9'b111111111;
assign micromatrizz[74][244] = 9'b111111111;
assign micromatrizz[74][245] = 9'b111111111;
assign micromatrizz[74][246] = 9'b111111111;
assign micromatrizz[74][247] = 9'b111111111;
assign micromatrizz[74][248] = 9'b111111111;
assign micromatrizz[74][249] = 9'b111111111;
assign micromatrizz[74][250] = 9'b111111111;
assign micromatrizz[74][251] = 9'b111111111;
assign micromatrizz[74][252] = 9'b111111111;
assign micromatrizz[74][253] = 9'b111111111;
assign micromatrizz[74][254] = 9'b111111111;
assign micromatrizz[74][255] = 9'b111111111;
assign micromatrizz[74][256] = 9'b111111111;
assign micromatrizz[74][257] = 9'b111111111;
assign micromatrizz[74][258] = 9'b111111111;
assign micromatrizz[74][259] = 9'b111111111;
assign micromatrizz[74][260] = 9'b111111111;
assign micromatrizz[74][261] = 9'b111111111;
assign micromatrizz[74][262] = 9'b111111111;
assign micromatrizz[74][263] = 9'b111111111;
assign micromatrizz[74][264] = 9'b111111111;
assign micromatrizz[74][265] = 9'b111111111;
assign micromatrizz[74][266] = 9'b111111111;
assign micromatrizz[74][267] = 9'b111111111;
assign micromatrizz[74][268] = 9'b111111111;
assign micromatrizz[74][269] = 9'b111111111;
assign micromatrizz[74][270] = 9'b111111111;
assign micromatrizz[74][271] = 9'b111111111;
assign micromatrizz[74][272] = 9'b111111111;
assign micromatrizz[74][273] = 9'b111111111;
assign micromatrizz[74][274] = 9'b111111111;
assign micromatrizz[74][275] = 9'b111111111;
assign micromatrizz[74][276] = 9'b111111111;
assign micromatrizz[74][277] = 9'b111111111;
assign micromatrizz[74][278] = 9'b111111111;
assign micromatrizz[74][279] = 9'b111111111;
assign micromatrizz[74][280] = 9'b111111111;
assign micromatrizz[74][281] = 9'b111111111;
assign micromatrizz[74][282] = 9'b111111111;
assign micromatrizz[74][283] = 9'b111111111;
assign micromatrizz[74][284] = 9'b111111111;
assign micromatrizz[74][285] = 9'b111111111;
assign micromatrizz[74][286] = 9'b111111111;
assign micromatrizz[74][287] = 9'b111111111;
assign micromatrizz[74][288] = 9'b111111111;
assign micromatrizz[74][289] = 9'b111111111;
assign micromatrizz[74][290] = 9'b111111111;
assign micromatrizz[74][291] = 9'b111111111;
assign micromatrizz[74][292] = 9'b111111111;
assign micromatrizz[74][293] = 9'b111111111;
assign micromatrizz[74][294] = 9'b111111111;
assign micromatrizz[74][295] = 9'b111111111;
assign micromatrizz[74][296] = 9'b111111111;
assign micromatrizz[74][297] = 9'b111111111;
assign micromatrizz[74][298] = 9'b111111111;
assign micromatrizz[74][299] = 9'b111111111;
assign micromatrizz[74][300] = 9'b111111111;
assign micromatrizz[74][301] = 9'b111111111;
assign micromatrizz[74][302] = 9'b111111111;
assign micromatrizz[74][303] = 9'b111111111;
assign micromatrizz[74][304] = 9'b111111111;
assign micromatrizz[74][305] = 9'b111111111;
assign micromatrizz[74][306] = 9'b111111111;
assign micromatrizz[74][307] = 9'b111111111;
assign micromatrizz[74][308] = 9'b111111111;
assign micromatrizz[74][309] = 9'b111111111;
assign micromatrizz[74][310] = 9'b111111111;
assign micromatrizz[74][311] = 9'b111111111;
assign micromatrizz[74][312] = 9'b111111111;
assign micromatrizz[74][313] = 9'b111111111;
assign micromatrizz[74][314] = 9'b111111111;
assign micromatrizz[74][315] = 9'b111111111;
assign micromatrizz[74][316] = 9'b111111111;
assign micromatrizz[74][317] = 9'b111111111;
assign micromatrizz[74][318] = 9'b111111111;
assign micromatrizz[74][319] = 9'b111111111;
assign micromatrizz[74][320] = 9'b111111111;
assign micromatrizz[74][321] = 9'b111111111;
assign micromatrizz[74][322] = 9'b111111111;
assign micromatrizz[74][323] = 9'b111111111;
assign micromatrizz[74][324] = 9'b111111111;
assign micromatrizz[74][325] = 9'b111111111;
assign micromatrizz[74][326] = 9'b111111111;
assign micromatrizz[74][327] = 9'b111111111;
assign micromatrizz[74][328] = 9'b111111111;
assign micromatrizz[74][329] = 9'b111111111;
assign micromatrizz[74][330] = 9'b111111111;
assign micromatrizz[74][331] = 9'b111111111;
assign micromatrizz[74][332] = 9'b111111111;
assign micromatrizz[74][333] = 9'b111111111;
assign micromatrizz[74][334] = 9'b111111111;
assign micromatrizz[74][335] = 9'b111111111;
assign micromatrizz[74][336] = 9'b111111111;
assign micromatrizz[74][337] = 9'b111111111;
assign micromatrizz[74][338] = 9'b111111111;
assign micromatrizz[74][339] = 9'b111111111;
assign micromatrizz[74][340] = 9'b111111111;
assign micromatrizz[74][341] = 9'b111111111;
assign micromatrizz[74][342] = 9'b111111111;
assign micromatrizz[74][343] = 9'b111111111;
assign micromatrizz[74][344] = 9'b111111111;
assign micromatrizz[74][345] = 9'b111111111;
assign micromatrizz[74][346] = 9'b111111111;
assign micromatrizz[74][347] = 9'b111111111;
assign micromatrizz[74][348] = 9'b111111111;
assign micromatrizz[74][349] = 9'b111111111;
assign micromatrizz[74][350] = 9'b111111111;
assign micromatrizz[74][351] = 9'b111111111;
assign micromatrizz[74][352] = 9'b111111111;
assign micromatrizz[74][353] = 9'b111111111;
assign micromatrizz[74][354] = 9'b111111111;
assign micromatrizz[74][355] = 9'b111111111;
assign micromatrizz[74][356] = 9'b111111111;
assign micromatrizz[74][357] = 9'b111111111;
assign micromatrizz[74][358] = 9'b111111111;
assign micromatrizz[74][359] = 9'b111111111;
assign micromatrizz[74][360] = 9'b111111111;
assign micromatrizz[74][361] = 9'b111111111;
assign micromatrizz[74][362] = 9'b111111111;
assign micromatrizz[74][363] = 9'b111111111;
assign micromatrizz[74][364] = 9'b111111111;
assign micromatrizz[74][365] = 9'b111111111;
assign micromatrizz[74][366] = 9'b111111111;
assign micromatrizz[74][367] = 9'b111111111;
assign micromatrizz[74][368] = 9'b111111111;
assign micromatrizz[74][369] = 9'b111111111;
assign micromatrizz[74][370] = 9'b111111111;
assign micromatrizz[74][371] = 9'b111111111;
assign micromatrizz[74][372] = 9'b111111111;
assign micromatrizz[74][373] = 9'b111111111;
assign micromatrizz[74][374] = 9'b111111111;
assign micromatrizz[74][375] = 9'b111111111;
assign micromatrizz[74][376] = 9'b111111111;
assign micromatrizz[74][377] = 9'b111111111;
assign micromatrizz[74][378] = 9'b111111111;
assign micromatrizz[74][379] = 9'b111111111;
assign micromatrizz[74][380] = 9'b111111111;
assign micromatrizz[74][381] = 9'b111111111;
assign micromatrizz[74][382] = 9'b111111111;
assign micromatrizz[74][383] = 9'b111111111;
assign micromatrizz[74][384] = 9'b111111111;
assign micromatrizz[74][385] = 9'b111111111;
assign micromatrizz[74][386] = 9'b111111111;
assign micromatrizz[74][387] = 9'b111111111;
assign micromatrizz[74][388] = 9'b111111111;
assign micromatrizz[74][389] = 9'b111111111;
assign micromatrizz[74][390] = 9'b111111111;
assign micromatrizz[74][391] = 9'b111111111;
assign micromatrizz[74][392] = 9'b111111111;
assign micromatrizz[74][393] = 9'b111111111;
assign micromatrizz[74][394] = 9'b111111111;
assign micromatrizz[74][395] = 9'b111111111;
assign micromatrizz[74][396] = 9'b111111111;
assign micromatrizz[74][397] = 9'b111111111;
assign micromatrizz[74][398] = 9'b111111111;
assign micromatrizz[74][399] = 9'b111111111;
assign micromatrizz[74][400] = 9'b111111111;
assign micromatrizz[74][401] = 9'b111111111;
assign micromatrizz[74][402] = 9'b111111111;
assign micromatrizz[74][403] = 9'b111111111;
assign micromatrizz[74][404] = 9'b111111111;
assign micromatrizz[74][405] = 9'b111111111;
assign micromatrizz[74][406] = 9'b111111111;
assign micromatrizz[74][407] = 9'b111111111;
assign micromatrizz[74][408] = 9'b111111111;
assign micromatrizz[74][409] = 9'b111111111;
assign micromatrizz[74][410] = 9'b111111111;
assign micromatrizz[74][411] = 9'b111111111;
assign micromatrizz[74][412] = 9'b111111111;
assign micromatrizz[74][413] = 9'b111111111;
assign micromatrizz[74][414] = 9'b111111111;
assign micromatrizz[74][415] = 9'b111111111;
assign micromatrizz[74][416] = 9'b111111111;
assign micromatrizz[74][417] = 9'b111111111;
assign micromatrizz[74][418] = 9'b111111111;
assign micromatrizz[74][419] = 9'b111111111;
assign micromatrizz[74][420] = 9'b111111111;
assign micromatrizz[74][421] = 9'b111111111;
assign micromatrizz[74][422] = 9'b111111111;
assign micromatrizz[74][423] = 9'b111111111;
assign micromatrizz[74][424] = 9'b111111111;
assign micromatrizz[74][425] = 9'b111111111;
assign micromatrizz[74][426] = 9'b111111111;
assign micromatrizz[74][427] = 9'b111111111;
assign micromatrizz[74][428] = 9'b111111111;
assign micromatrizz[74][429] = 9'b111111111;
assign micromatrizz[74][430] = 9'b111111111;
assign micromatrizz[74][431] = 9'b111111111;
assign micromatrizz[74][432] = 9'b111111111;
assign micromatrizz[74][433] = 9'b111111111;
assign micromatrizz[74][434] = 9'b111111111;
assign micromatrizz[74][435] = 9'b111111111;
assign micromatrizz[74][436] = 9'b111111111;
assign micromatrizz[74][437] = 9'b111111111;
assign micromatrizz[74][438] = 9'b111111111;
assign micromatrizz[74][439] = 9'b111111111;
assign micromatrizz[74][440] = 9'b111111111;
assign micromatrizz[74][441] = 9'b111111111;
assign micromatrizz[74][442] = 9'b111111111;
assign micromatrizz[74][443] = 9'b111111111;
assign micromatrizz[74][444] = 9'b111111111;
assign micromatrizz[74][445] = 9'b111111111;
assign micromatrizz[74][446] = 9'b111111111;
assign micromatrizz[74][447] = 9'b111111111;
assign micromatrizz[74][448] = 9'b111111111;
assign micromatrizz[74][449] = 9'b111111111;
assign micromatrizz[74][450] = 9'b111111111;
assign micromatrizz[74][451] = 9'b111111111;
assign micromatrizz[74][452] = 9'b111111111;
assign micromatrizz[74][453] = 9'b111111111;
assign micromatrizz[74][454] = 9'b111111111;
assign micromatrizz[74][455] = 9'b111111111;
assign micromatrizz[74][456] = 9'b111111111;
assign micromatrizz[74][457] = 9'b111111111;
assign micromatrizz[74][458] = 9'b111111111;
assign micromatrizz[74][459] = 9'b111111111;
assign micromatrizz[74][460] = 9'b111111111;
assign micromatrizz[74][461] = 9'b111111111;
assign micromatrizz[74][462] = 9'b111111111;
assign micromatrizz[74][463] = 9'b111111111;
assign micromatrizz[74][464] = 9'b111111111;
assign micromatrizz[74][465] = 9'b111111111;
assign micromatrizz[74][466] = 9'b111111111;
assign micromatrizz[74][467] = 9'b111111111;
assign micromatrizz[74][468] = 9'b111111111;
assign micromatrizz[74][469] = 9'b111111111;
assign micromatrizz[74][470] = 9'b111111111;
assign micromatrizz[74][471] = 9'b111111111;
assign micromatrizz[74][472] = 9'b111111111;
assign micromatrizz[74][473] = 9'b111111111;
assign micromatrizz[74][474] = 9'b111111111;
assign micromatrizz[74][475] = 9'b111111111;
assign micromatrizz[74][476] = 9'b111111111;
assign micromatrizz[74][477] = 9'b111111111;
assign micromatrizz[74][478] = 9'b111111111;
assign micromatrizz[74][479] = 9'b111111111;
assign micromatrizz[74][480] = 9'b111111111;
assign micromatrizz[74][481] = 9'b111111111;
assign micromatrizz[74][482] = 9'b111111111;
assign micromatrizz[74][483] = 9'b111111111;
assign micromatrizz[74][484] = 9'b111111111;
assign micromatrizz[74][485] = 9'b111111111;
assign micromatrizz[74][486] = 9'b111111111;
assign micromatrizz[74][487] = 9'b111111111;
assign micromatrizz[74][488] = 9'b111111111;
assign micromatrizz[74][489] = 9'b111111111;
assign micromatrizz[74][490] = 9'b111111111;
assign micromatrizz[74][491] = 9'b111111111;
assign micromatrizz[74][492] = 9'b111111111;
assign micromatrizz[74][493] = 9'b111111111;
assign micromatrizz[74][494] = 9'b111111111;
assign micromatrizz[74][495] = 9'b111111111;
assign micromatrizz[74][496] = 9'b111111111;
assign micromatrizz[74][497] = 9'b111111111;
assign micromatrizz[74][498] = 9'b111111111;
assign micromatrizz[74][499] = 9'b111111111;
assign micromatrizz[74][500] = 9'b111111111;
assign micromatrizz[74][501] = 9'b111111111;
assign micromatrizz[74][502] = 9'b111111111;
assign micromatrizz[74][503] = 9'b111111111;
assign micromatrizz[74][504] = 9'b111111111;
assign micromatrizz[74][505] = 9'b111111111;
assign micromatrizz[74][506] = 9'b111111111;
assign micromatrizz[74][507] = 9'b111111111;
assign micromatrizz[74][508] = 9'b111111111;
assign micromatrizz[74][509] = 9'b111111111;
assign micromatrizz[74][510] = 9'b111111111;
assign micromatrizz[74][511] = 9'b111111111;
assign micromatrizz[74][512] = 9'b111111111;
assign micromatrizz[74][513] = 9'b111111111;
assign micromatrizz[74][514] = 9'b111111111;
assign micromatrizz[74][515] = 9'b111111111;
assign micromatrizz[74][516] = 9'b111111111;
assign micromatrizz[74][517] = 9'b111111111;
assign micromatrizz[74][518] = 9'b111111111;
assign micromatrizz[74][519] = 9'b111111111;
assign micromatrizz[74][520] = 9'b111111111;
assign micromatrizz[74][521] = 9'b111111111;
assign micromatrizz[74][522] = 9'b111111111;
assign micromatrizz[74][523] = 9'b111111111;
assign micromatrizz[74][524] = 9'b111111111;
assign micromatrizz[74][525] = 9'b111111111;
assign micromatrizz[74][526] = 9'b111111111;
assign micromatrizz[74][527] = 9'b111111111;
assign micromatrizz[74][528] = 9'b111111111;
assign micromatrizz[74][529] = 9'b111111111;
assign micromatrizz[74][530] = 9'b111111111;
assign micromatrizz[74][531] = 9'b111111111;
assign micromatrizz[74][532] = 9'b111111111;
assign micromatrizz[74][533] = 9'b111111111;
assign micromatrizz[74][534] = 9'b111111111;
assign micromatrizz[74][535] = 9'b111111111;
assign micromatrizz[74][536] = 9'b111111111;
assign micromatrizz[74][537] = 9'b111111111;
assign micromatrizz[74][538] = 9'b111111111;
assign micromatrizz[74][539] = 9'b111111111;
assign micromatrizz[74][540] = 9'b111111111;
assign micromatrizz[74][541] = 9'b111111111;
assign micromatrizz[74][542] = 9'b111111111;
assign micromatrizz[74][543] = 9'b111111111;
assign micromatrizz[74][544] = 9'b111111111;
assign micromatrizz[74][545] = 9'b111111111;
assign micromatrizz[74][546] = 9'b111111111;
assign micromatrizz[74][547] = 9'b111111111;
assign micromatrizz[74][548] = 9'b111111111;
assign micromatrizz[74][549] = 9'b111111111;
assign micromatrizz[74][550] = 9'b111111111;
assign micromatrizz[74][551] = 9'b111111111;
assign micromatrizz[74][552] = 9'b111111111;
assign micromatrizz[74][553] = 9'b111111111;
assign micromatrizz[74][554] = 9'b111111111;
assign micromatrizz[74][555] = 9'b111111111;
assign micromatrizz[74][556] = 9'b111111111;
assign micromatrizz[74][557] = 9'b111111111;
assign micromatrizz[74][558] = 9'b111111111;
assign micromatrizz[74][559] = 9'b111111111;
assign micromatrizz[74][560] = 9'b111111111;
assign micromatrizz[74][561] = 9'b111111111;
assign micromatrizz[74][562] = 9'b111111111;
assign micromatrizz[74][563] = 9'b111111111;
assign micromatrizz[74][564] = 9'b111111111;
assign micromatrizz[74][565] = 9'b111111111;
assign micromatrizz[74][566] = 9'b111111111;
assign micromatrizz[74][567] = 9'b111111111;
assign micromatrizz[74][568] = 9'b111111111;
assign micromatrizz[74][569] = 9'b111111111;
assign micromatrizz[74][570] = 9'b111111111;
assign micromatrizz[74][571] = 9'b111111111;
assign micromatrizz[74][572] = 9'b111111111;
assign micromatrizz[74][573] = 9'b111111111;
assign micromatrizz[74][574] = 9'b111111111;
assign micromatrizz[74][575] = 9'b111111111;
assign micromatrizz[74][576] = 9'b111111111;
assign micromatrizz[74][577] = 9'b111111111;
assign micromatrizz[74][578] = 9'b111111111;
assign micromatrizz[74][579] = 9'b111111111;
assign micromatrizz[74][580] = 9'b111111111;
assign micromatrizz[74][581] = 9'b111111111;
assign micromatrizz[74][582] = 9'b111111111;
assign micromatrizz[74][583] = 9'b111111111;
assign micromatrizz[74][584] = 9'b111111111;
assign micromatrizz[74][585] = 9'b111111111;
assign micromatrizz[74][586] = 9'b111111111;
assign micromatrizz[74][587] = 9'b111111111;
assign micromatrizz[74][588] = 9'b111111111;
assign micromatrizz[74][589] = 9'b111111111;
assign micromatrizz[74][590] = 9'b111111111;
assign micromatrizz[74][591] = 9'b111111111;
assign micromatrizz[74][592] = 9'b111111111;
assign micromatrizz[74][593] = 9'b111111111;
assign micromatrizz[74][594] = 9'b111111111;
assign micromatrizz[74][595] = 9'b111111111;
assign micromatrizz[74][596] = 9'b111111111;
assign micromatrizz[74][597] = 9'b111111111;
assign micromatrizz[74][598] = 9'b111111111;
assign micromatrizz[74][599] = 9'b111111111;
assign micromatrizz[74][600] = 9'b111111111;
assign micromatrizz[74][601] = 9'b111111111;
assign micromatrizz[74][602] = 9'b111111111;
assign micromatrizz[74][603] = 9'b111111111;
assign micromatrizz[74][604] = 9'b111111111;
assign micromatrizz[74][605] = 9'b111111111;
assign micromatrizz[74][606] = 9'b111111111;
assign micromatrizz[74][607] = 9'b111111111;
assign micromatrizz[74][608] = 9'b111111111;
assign micromatrizz[74][609] = 9'b111111111;
assign micromatrizz[74][610] = 9'b111111111;
assign micromatrizz[74][611] = 9'b111111111;
assign micromatrizz[74][612] = 9'b111111111;
assign micromatrizz[74][613] = 9'b111111111;
assign micromatrizz[74][614] = 9'b111111111;
assign micromatrizz[74][615] = 9'b111111111;
assign micromatrizz[74][616] = 9'b111111111;
assign micromatrizz[74][617] = 9'b111111111;
assign micromatrizz[74][618] = 9'b111111111;
assign micromatrizz[74][619] = 9'b111111111;
assign micromatrizz[74][620] = 9'b111111111;
assign micromatrizz[74][621] = 9'b111111111;
assign micromatrizz[74][622] = 9'b111111111;
assign micromatrizz[74][623] = 9'b111111111;
assign micromatrizz[74][624] = 9'b111111111;
assign micromatrizz[74][625] = 9'b111111111;
assign micromatrizz[74][626] = 9'b111111111;
assign micromatrizz[74][627] = 9'b111111111;
assign micromatrizz[74][628] = 9'b111111111;
assign micromatrizz[74][629] = 9'b111111111;
assign micromatrizz[74][630] = 9'b111111111;
assign micromatrizz[74][631] = 9'b111111111;
assign micromatrizz[74][632] = 9'b111111111;
assign micromatrizz[74][633] = 9'b111111111;
assign micromatrizz[74][634] = 9'b111111111;
assign micromatrizz[74][635] = 9'b111111111;
assign micromatrizz[74][636] = 9'b111111111;
assign micromatrizz[74][637] = 9'b111111111;
assign micromatrizz[74][638] = 9'b111111111;
assign micromatrizz[74][639] = 9'b111111111;
assign micromatrizz[75][0] = 9'b111111111;
assign micromatrizz[75][1] = 9'b111111111;
assign micromatrizz[75][2] = 9'b111111111;
assign micromatrizz[75][3] = 9'b111111111;
assign micromatrizz[75][4] = 9'b111111111;
assign micromatrizz[75][5] = 9'b111111111;
assign micromatrizz[75][6] = 9'b111111111;
assign micromatrizz[75][7] = 9'b111111111;
assign micromatrizz[75][8] = 9'b111111111;
assign micromatrizz[75][9] = 9'b111111111;
assign micromatrizz[75][10] = 9'b111111111;
assign micromatrizz[75][11] = 9'b111111111;
assign micromatrizz[75][12] = 9'b111111111;
assign micromatrizz[75][13] = 9'b111111111;
assign micromatrizz[75][14] = 9'b111111111;
assign micromatrizz[75][15] = 9'b111111111;
assign micromatrizz[75][16] = 9'b111111111;
assign micromatrizz[75][17] = 9'b111111111;
assign micromatrizz[75][18] = 9'b111111111;
assign micromatrizz[75][19] = 9'b111111111;
assign micromatrizz[75][20] = 9'b111111111;
assign micromatrizz[75][21] = 9'b111111111;
assign micromatrizz[75][22] = 9'b111111111;
assign micromatrizz[75][23] = 9'b111111111;
assign micromatrizz[75][24] = 9'b111111111;
assign micromatrizz[75][25] = 9'b111111111;
assign micromatrizz[75][26] = 9'b111111111;
assign micromatrizz[75][27] = 9'b111111111;
assign micromatrizz[75][28] = 9'b111111111;
assign micromatrizz[75][29] = 9'b111111111;
assign micromatrizz[75][30] = 9'b111111111;
assign micromatrizz[75][31] = 9'b111111111;
assign micromatrizz[75][32] = 9'b111111111;
assign micromatrizz[75][33] = 9'b111111111;
assign micromatrizz[75][34] = 9'b111111111;
assign micromatrizz[75][35] = 9'b111111111;
assign micromatrizz[75][36] = 9'b111111111;
assign micromatrizz[75][37] = 9'b111111111;
assign micromatrizz[75][38] = 9'b111111111;
assign micromatrizz[75][39] = 9'b111111111;
assign micromatrizz[75][40] = 9'b111111111;
assign micromatrizz[75][41] = 9'b111111111;
assign micromatrizz[75][42] = 9'b111111111;
assign micromatrizz[75][43] = 9'b111111111;
assign micromatrizz[75][44] = 9'b111111111;
assign micromatrizz[75][45] = 9'b111111111;
assign micromatrizz[75][46] = 9'b111111111;
assign micromatrizz[75][47] = 9'b111111111;
assign micromatrizz[75][48] = 9'b111111111;
assign micromatrizz[75][49] = 9'b111111111;
assign micromatrizz[75][50] = 9'b111111111;
assign micromatrizz[75][51] = 9'b111111111;
assign micromatrizz[75][52] = 9'b111111111;
assign micromatrizz[75][53] = 9'b111111111;
assign micromatrizz[75][54] = 9'b111111111;
assign micromatrizz[75][55] = 9'b111111111;
assign micromatrizz[75][56] = 9'b111111111;
assign micromatrizz[75][57] = 9'b111111111;
assign micromatrizz[75][58] = 9'b111111111;
assign micromatrizz[75][59] = 9'b111111111;
assign micromatrizz[75][60] = 9'b111111111;
assign micromatrizz[75][61] = 9'b111111111;
assign micromatrizz[75][62] = 9'b111111111;
assign micromatrizz[75][63] = 9'b111111111;
assign micromatrizz[75][64] = 9'b111111111;
assign micromatrizz[75][65] = 9'b111111111;
assign micromatrizz[75][66] = 9'b111111111;
assign micromatrizz[75][67] = 9'b111111111;
assign micromatrizz[75][68] = 9'b111111111;
assign micromatrizz[75][69] = 9'b111111111;
assign micromatrizz[75][70] = 9'b111111111;
assign micromatrizz[75][71] = 9'b111111111;
assign micromatrizz[75][72] = 9'b111111111;
assign micromatrizz[75][73] = 9'b111111111;
assign micromatrizz[75][74] = 9'b111111111;
assign micromatrizz[75][75] = 9'b111111111;
assign micromatrizz[75][76] = 9'b111111111;
assign micromatrizz[75][77] = 9'b111111111;
assign micromatrizz[75][78] = 9'b111111111;
assign micromatrizz[75][79] = 9'b111111111;
assign micromatrizz[75][80] = 9'b111111111;
assign micromatrizz[75][81] = 9'b111111111;
assign micromatrizz[75][82] = 9'b111111111;
assign micromatrizz[75][83] = 9'b111111111;
assign micromatrizz[75][84] = 9'b111111111;
assign micromatrizz[75][85] = 9'b111111111;
assign micromatrizz[75][86] = 9'b111111111;
assign micromatrizz[75][87] = 9'b111111111;
assign micromatrizz[75][88] = 9'b111111111;
assign micromatrizz[75][89] = 9'b111111111;
assign micromatrizz[75][90] = 9'b111111111;
assign micromatrizz[75][91] = 9'b111111111;
assign micromatrizz[75][92] = 9'b111111111;
assign micromatrizz[75][93] = 9'b111111111;
assign micromatrizz[75][94] = 9'b111111111;
assign micromatrizz[75][95] = 9'b111111111;
assign micromatrizz[75][96] = 9'b111111111;
assign micromatrizz[75][97] = 9'b111111111;
assign micromatrizz[75][98] = 9'b111111111;
assign micromatrizz[75][99] = 9'b111111111;
assign micromatrizz[75][100] = 9'b111111111;
assign micromatrizz[75][101] = 9'b111111111;
assign micromatrizz[75][102] = 9'b111111111;
assign micromatrizz[75][103] = 9'b111111111;
assign micromatrizz[75][104] = 9'b111111111;
assign micromatrizz[75][105] = 9'b111111111;
assign micromatrizz[75][106] = 9'b111111111;
assign micromatrizz[75][107] = 9'b111111111;
assign micromatrizz[75][108] = 9'b111111111;
assign micromatrizz[75][109] = 9'b111111111;
assign micromatrizz[75][110] = 9'b111111111;
assign micromatrizz[75][111] = 9'b111111111;
assign micromatrizz[75][112] = 9'b111111111;
assign micromatrizz[75][113] = 9'b111111111;
assign micromatrizz[75][114] = 9'b111111111;
assign micromatrizz[75][115] = 9'b111111111;
assign micromatrizz[75][116] = 9'b111111111;
assign micromatrizz[75][117] = 9'b111111111;
assign micromatrizz[75][118] = 9'b111111111;
assign micromatrizz[75][119] = 9'b111111111;
assign micromatrizz[75][120] = 9'b111111111;
assign micromatrizz[75][121] = 9'b111111111;
assign micromatrizz[75][122] = 9'b111111111;
assign micromatrizz[75][123] = 9'b111111111;
assign micromatrizz[75][124] = 9'b111111111;
assign micromatrizz[75][125] = 9'b111111111;
assign micromatrizz[75][126] = 9'b111111111;
assign micromatrizz[75][127] = 9'b111111111;
assign micromatrizz[75][128] = 9'b111111111;
assign micromatrizz[75][129] = 9'b111111111;
assign micromatrizz[75][130] = 9'b111111111;
assign micromatrizz[75][131] = 9'b111111111;
assign micromatrizz[75][132] = 9'b111111111;
assign micromatrizz[75][133] = 9'b111111111;
assign micromatrizz[75][134] = 9'b111111111;
assign micromatrizz[75][135] = 9'b111111111;
assign micromatrizz[75][136] = 9'b111111111;
assign micromatrizz[75][137] = 9'b111111111;
assign micromatrizz[75][138] = 9'b111111111;
assign micromatrizz[75][139] = 9'b111111111;
assign micromatrizz[75][140] = 9'b111111111;
assign micromatrizz[75][141] = 9'b111111111;
assign micromatrizz[75][142] = 9'b111111111;
assign micromatrizz[75][143] = 9'b111111111;
assign micromatrizz[75][144] = 9'b111111111;
assign micromatrizz[75][145] = 9'b111111111;
assign micromatrizz[75][146] = 9'b111111111;
assign micromatrizz[75][147] = 9'b111111111;
assign micromatrizz[75][148] = 9'b111111111;
assign micromatrizz[75][149] = 9'b111111111;
assign micromatrizz[75][150] = 9'b111111111;
assign micromatrizz[75][151] = 9'b111111111;
assign micromatrizz[75][152] = 9'b111111111;
assign micromatrizz[75][153] = 9'b111111111;
assign micromatrizz[75][154] = 9'b111111111;
assign micromatrizz[75][155] = 9'b111111111;
assign micromatrizz[75][156] = 9'b111111111;
assign micromatrizz[75][157] = 9'b111111111;
assign micromatrizz[75][158] = 9'b111111111;
assign micromatrizz[75][159] = 9'b111111111;
assign micromatrizz[75][160] = 9'b111111111;
assign micromatrizz[75][161] = 9'b111111111;
assign micromatrizz[75][162] = 9'b111111111;
assign micromatrizz[75][163] = 9'b111111111;
assign micromatrizz[75][164] = 9'b111111111;
assign micromatrizz[75][165] = 9'b111111111;
assign micromatrizz[75][166] = 9'b111111111;
assign micromatrizz[75][167] = 9'b111111111;
assign micromatrizz[75][168] = 9'b111111111;
assign micromatrizz[75][169] = 9'b111111111;
assign micromatrizz[75][170] = 9'b111111111;
assign micromatrizz[75][171] = 9'b111111111;
assign micromatrizz[75][172] = 9'b111111111;
assign micromatrizz[75][173] = 9'b111111111;
assign micromatrizz[75][174] = 9'b111111111;
assign micromatrizz[75][175] = 9'b111111111;
assign micromatrizz[75][176] = 9'b111111111;
assign micromatrizz[75][177] = 9'b111111111;
assign micromatrizz[75][178] = 9'b111111111;
assign micromatrizz[75][179] = 9'b111111111;
assign micromatrizz[75][180] = 9'b111111111;
assign micromatrizz[75][181] = 9'b111111111;
assign micromatrizz[75][182] = 9'b111111111;
assign micromatrizz[75][183] = 9'b111111111;
assign micromatrizz[75][184] = 9'b111111111;
assign micromatrizz[75][185] = 9'b111111111;
assign micromatrizz[75][186] = 9'b111111111;
assign micromatrizz[75][187] = 9'b111111111;
assign micromatrizz[75][188] = 9'b111111111;
assign micromatrizz[75][189] = 9'b111111111;
assign micromatrizz[75][190] = 9'b111111111;
assign micromatrizz[75][191] = 9'b111111111;
assign micromatrizz[75][192] = 9'b111111111;
assign micromatrizz[75][193] = 9'b111111111;
assign micromatrizz[75][194] = 9'b111111111;
assign micromatrizz[75][195] = 9'b111111111;
assign micromatrizz[75][196] = 9'b111111111;
assign micromatrizz[75][197] = 9'b111111111;
assign micromatrizz[75][198] = 9'b111111111;
assign micromatrizz[75][199] = 9'b111111111;
assign micromatrizz[75][200] = 9'b111111111;
assign micromatrizz[75][201] = 9'b111111111;
assign micromatrizz[75][202] = 9'b111111111;
assign micromatrizz[75][203] = 9'b111111111;
assign micromatrizz[75][204] = 9'b111111111;
assign micromatrizz[75][205] = 9'b111111111;
assign micromatrizz[75][206] = 9'b111111111;
assign micromatrizz[75][207] = 9'b111111111;
assign micromatrizz[75][208] = 9'b111111111;
assign micromatrizz[75][209] = 9'b111111111;
assign micromatrizz[75][210] = 9'b111111111;
assign micromatrizz[75][211] = 9'b111111111;
assign micromatrizz[75][212] = 9'b111111111;
assign micromatrizz[75][213] = 9'b111111111;
assign micromatrizz[75][214] = 9'b111111111;
assign micromatrizz[75][215] = 9'b111111111;
assign micromatrizz[75][216] = 9'b111111111;
assign micromatrizz[75][217] = 9'b111111111;
assign micromatrizz[75][218] = 9'b111111111;
assign micromatrizz[75][219] = 9'b111111111;
assign micromatrizz[75][220] = 9'b111111111;
assign micromatrizz[75][221] = 9'b111111111;
assign micromatrizz[75][222] = 9'b111111111;
assign micromatrizz[75][223] = 9'b111111111;
assign micromatrizz[75][224] = 9'b111111111;
assign micromatrizz[75][225] = 9'b111111111;
assign micromatrizz[75][226] = 9'b111111111;
assign micromatrizz[75][227] = 9'b111111111;
assign micromatrizz[75][228] = 9'b111111111;
assign micromatrizz[75][229] = 9'b111111111;
assign micromatrizz[75][230] = 9'b111111111;
assign micromatrizz[75][231] = 9'b111111111;
assign micromatrizz[75][232] = 9'b111111111;
assign micromatrizz[75][233] = 9'b111111111;
assign micromatrizz[75][234] = 9'b111111111;
assign micromatrizz[75][235] = 9'b111111111;
assign micromatrizz[75][236] = 9'b111111111;
assign micromatrizz[75][237] = 9'b111111111;
assign micromatrizz[75][238] = 9'b111111111;
assign micromatrizz[75][239] = 9'b111111111;
assign micromatrizz[75][240] = 9'b111111111;
assign micromatrizz[75][241] = 9'b111111111;
assign micromatrizz[75][242] = 9'b111111111;
assign micromatrizz[75][243] = 9'b111111111;
assign micromatrizz[75][244] = 9'b111111111;
assign micromatrizz[75][245] = 9'b111111111;
assign micromatrizz[75][246] = 9'b111111111;
assign micromatrizz[75][247] = 9'b111111111;
assign micromatrizz[75][248] = 9'b111111111;
assign micromatrizz[75][249] = 9'b111111111;
assign micromatrizz[75][250] = 9'b111111111;
assign micromatrizz[75][251] = 9'b111111111;
assign micromatrizz[75][252] = 9'b111111111;
assign micromatrizz[75][253] = 9'b111111111;
assign micromatrizz[75][254] = 9'b111111111;
assign micromatrizz[75][255] = 9'b111111111;
assign micromatrizz[75][256] = 9'b111111111;
assign micromatrizz[75][257] = 9'b111111111;
assign micromatrizz[75][258] = 9'b111111111;
assign micromatrizz[75][259] = 9'b111111111;
assign micromatrizz[75][260] = 9'b111111111;
assign micromatrizz[75][261] = 9'b111111111;
assign micromatrizz[75][262] = 9'b111111111;
assign micromatrizz[75][263] = 9'b111111111;
assign micromatrizz[75][264] = 9'b111111111;
assign micromatrizz[75][265] = 9'b111111111;
assign micromatrizz[75][266] = 9'b111111111;
assign micromatrizz[75][267] = 9'b111111111;
assign micromatrizz[75][268] = 9'b111111111;
assign micromatrizz[75][269] = 9'b111111111;
assign micromatrizz[75][270] = 9'b111111111;
assign micromatrizz[75][271] = 9'b111111111;
assign micromatrizz[75][272] = 9'b111111111;
assign micromatrizz[75][273] = 9'b111111111;
assign micromatrizz[75][274] = 9'b111111111;
assign micromatrizz[75][275] = 9'b111111111;
assign micromatrizz[75][276] = 9'b111111111;
assign micromatrizz[75][277] = 9'b111111111;
assign micromatrizz[75][278] = 9'b111111111;
assign micromatrizz[75][279] = 9'b111111111;
assign micromatrizz[75][280] = 9'b111111111;
assign micromatrizz[75][281] = 9'b111111111;
assign micromatrizz[75][282] = 9'b111111111;
assign micromatrizz[75][283] = 9'b111111111;
assign micromatrizz[75][284] = 9'b111111111;
assign micromatrizz[75][285] = 9'b111111111;
assign micromatrizz[75][286] = 9'b111111111;
assign micromatrizz[75][287] = 9'b111111111;
assign micromatrizz[75][288] = 9'b111111111;
assign micromatrizz[75][289] = 9'b111111111;
assign micromatrizz[75][290] = 9'b111111111;
assign micromatrizz[75][291] = 9'b111111111;
assign micromatrizz[75][292] = 9'b111111111;
assign micromatrizz[75][293] = 9'b111111111;
assign micromatrizz[75][294] = 9'b111111111;
assign micromatrizz[75][295] = 9'b111111111;
assign micromatrizz[75][296] = 9'b111111111;
assign micromatrizz[75][297] = 9'b111111111;
assign micromatrizz[75][298] = 9'b111111111;
assign micromatrizz[75][299] = 9'b111111111;
assign micromatrizz[75][300] = 9'b111111111;
assign micromatrizz[75][301] = 9'b111111111;
assign micromatrizz[75][302] = 9'b111111111;
assign micromatrizz[75][303] = 9'b111111111;
assign micromatrizz[75][304] = 9'b111111111;
assign micromatrizz[75][305] = 9'b111111111;
assign micromatrizz[75][306] = 9'b111111111;
assign micromatrizz[75][307] = 9'b111111111;
assign micromatrizz[75][308] = 9'b111111111;
assign micromatrizz[75][309] = 9'b111111111;
assign micromatrizz[75][310] = 9'b111111111;
assign micromatrizz[75][311] = 9'b111111111;
assign micromatrizz[75][312] = 9'b111111111;
assign micromatrizz[75][313] = 9'b111111111;
assign micromatrizz[75][314] = 9'b111111111;
assign micromatrizz[75][315] = 9'b111111111;
assign micromatrizz[75][316] = 9'b111111111;
assign micromatrizz[75][317] = 9'b111111111;
assign micromatrizz[75][318] = 9'b111111111;
assign micromatrizz[75][319] = 9'b111111111;
assign micromatrizz[75][320] = 9'b111111111;
assign micromatrizz[75][321] = 9'b111111111;
assign micromatrizz[75][322] = 9'b111111111;
assign micromatrizz[75][323] = 9'b111111111;
assign micromatrizz[75][324] = 9'b111111111;
assign micromatrizz[75][325] = 9'b111111111;
assign micromatrizz[75][326] = 9'b111111111;
assign micromatrizz[75][327] = 9'b111111111;
assign micromatrizz[75][328] = 9'b111111111;
assign micromatrizz[75][329] = 9'b111111111;
assign micromatrizz[75][330] = 9'b111111111;
assign micromatrizz[75][331] = 9'b111111111;
assign micromatrizz[75][332] = 9'b111111111;
assign micromatrizz[75][333] = 9'b111111111;
assign micromatrizz[75][334] = 9'b111111111;
assign micromatrizz[75][335] = 9'b111111111;
assign micromatrizz[75][336] = 9'b111111111;
assign micromatrizz[75][337] = 9'b111111111;
assign micromatrizz[75][338] = 9'b111111111;
assign micromatrizz[75][339] = 9'b111111111;
assign micromatrizz[75][340] = 9'b111111111;
assign micromatrizz[75][341] = 9'b111111111;
assign micromatrizz[75][342] = 9'b111111111;
assign micromatrizz[75][343] = 9'b111111111;
assign micromatrizz[75][344] = 9'b111111111;
assign micromatrizz[75][345] = 9'b111111111;
assign micromatrizz[75][346] = 9'b111111111;
assign micromatrizz[75][347] = 9'b111111111;
assign micromatrizz[75][348] = 9'b111111111;
assign micromatrizz[75][349] = 9'b111111111;
assign micromatrizz[75][350] = 9'b111111111;
assign micromatrizz[75][351] = 9'b111111111;
assign micromatrizz[75][352] = 9'b111111111;
assign micromatrizz[75][353] = 9'b111111111;
assign micromatrizz[75][354] = 9'b111111111;
assign micromatrizz[75][355] = 9'b111111111;
assign micromatrizz[75][356] = 9'b111111111;
assign micromatrizz[75][357] = 9'b111111111;
assign micromatrizz[75][358] = 9'b111111111;
assign micromatrizz[75][359] = 9'b111111111;
assign micromatrizz[75][360] = 9'b111111111;
assign micromatrizz[75][361] = 9'b111111111;
assign micromatrizz[75][362] = 9'b111111111;
assign micromatrizz[75][363] = 9'b111111111;
assign micromatrizz[75][364] = 9'b111111111;
assign micromatrizz[75][365] = 9'b111111111;
assign micromatrizz[75][366] = 9'b111111111;
assign micromatrizz[75][367] = 9'b111111111;
assign micromatrizz[75][368] = 9'b111111111;
assign micromatrizz[75][369] = 9'b111111111;
assign micromatrizz[75][370] = 9'b111111111;
assign micromatrizz[75][371] = 9'b111111111;
assign micromatrizz[75][372] = 9'b111111111;
assign micromatrizz[75][373] = 9'b111111111;
assign micromatrizz[75][374] = 9'b111111111;
assign micromatrizz[75][375] = 9'b111111111;
assign micromatrizz[75][376] = 9'b111111111;
assign micromatrizz[75][377] = 9'b111111111;
assign micromatrizz[75][378] = 9'b111111111;
assign micromatrizz[75][379] = 9'b111111111;
assign micromatrizz[75][380] = 9'b111111111;
assign micromatrizz[75][381] = 9'b111111111;
assign micromatrizz[75][382] = 9'b111111111;
assign micromatrizz[75][383] = 9'b111111111;
assign micromatrizz[75][384] = 9'b111111111;
assign micromatrizz[75][385] = 9'b111111111;
assign micromatrizz[75][386] = 9'b111111111;
assign micromatrizz[75][387] = 9'b111111111;
assign micromatrizz[75][388] = 9'b111111111;
assign micromatrizz[75][389] = 9'b111111111;
assign micromatrizz[75][390] = 9'b111111111;
assign micromatrizz[75][391] = 9'b111111111;
assign micromatrizz[75][392] = 9'b111111111;
assign micromatrizz[75][393] = 9'b111111111;
assign micromatrizz[75][394] = 9'b111111111;
assign micromatrizz[75][395] = 9'b111111111;
assign micromatrizz[75][396] = 9'b111111111;
assign micromatrizz[75][397] = 9'b111111111;
assign micromatrizz[75][398] = 9'b111111111;
assign micromatrizz[75][399] = 9'b111111111;
assign micromatrizz[75][400] = 9'b111111111;
assign micromatrizz[75][401] = 9'b111111111;
assign micromatrizz[75][402] = 9'b111111111;
assign micromatrizz[75][403] = 9'b111111111;
assign micromatrizz[75][404] = 9'b111111111;
assign micromatrizz[75][405] = 9'b111111111;
assign micromatrizz[75][406] = 9'b111111111;
assign micromatrizz[75][407] = 9'b111111111;
assign micromatrizz[75][408] = 9'b111111111;
assign micromatrizz[75][409] = 9'b111111111;
assign micromatrizz[75][410] = 9'b111111111;
assign micromatrizz[75][411] = 9'b111111111;
assign micromatrizz[75][412] = 9'b111111111;
assign micromatrizz[75][413] = 9'b111111111;
assign micromatrizz[75][414] = 9'b111111111;
assign micromatrizz[75][415] = 9'b111111111;
assign micromatrizz[75][416] = 9'b111111111;
assign micromatrizz[75][417] = 9'b111111111;
assign micromatrizz[75][418] = 9'b111111111;
assign micromatrizz[75][419] = 9'b111111111;
assign micromatrizz[75][420] = 9'b111111111;
assign micromatrizz[75][421] = 9'b111111111;
assign micromatrizz[75][422] = 9'b111111111;
assign micromatrizz[75][423] = 9'b111111111;
assign micromatrizz[75][424] = 9'b111111111;
assign micromatrizz[75][425] = 9'b111111111;
assign micromatrizz[75][426] = 9'b111111111;
assign micromatrizz[75][427] = 9'b111111111;
assign micromatrizz[75][428] = 9'b111111111;
assign micromatrizz[75][429] = 9'b111111111;
assign micromatrizz[75][430] = 9'b111111111;
assign micromatrizz[75][431] = 9'b111111111;
assign micromatrizz[75][432] = 9'b111111111;
assign micromatrizz[75][433] = 9'b111111111;
assign micromatrizz[75][434] = 9'b111111111;
assign micromatrizz[75][435] = 9'b111111111;
assign micromatrizz[75][436] = 9'b111111111;
assign micromatrizz[75][437] = 9'b111111111;
assign micromatrizz[75][438] = 9'b111111111;
assign micromatrizz[75][439] = 9'b111111111;
assign micromatrizz[75][440] = 9'b111111111;
assign micromatrizz[75][441] = 9'b111111111;
assign micromatrizz[75][442] = 9'b111111111;
assign micromatrizz[75][443] = 9'b111111111;
assign micromatrizz[75][444] = 9'b111111111;
assign micromatrizz[75][445] = 9'b111111111;
assign micromatrizz[75][446] = 9'b111111111;
assign micromatrizz[75][447] = 9'b111111111;
assign micromatrizz[75][448] = 9'b111111111;
assign micromatrizz[75][449] = 9'b111111111;
assign micromatrizz[75][450] = 9'b111111111;
assign micromatrizz[75][451] = 9'b111111111;
assign micromatrizz[75][452] = 9'b111111111;
assign micromatrizz[75][453] = 9'b111111111;
assign micromatrizz[75][454] = 9'b111111111;
assign micromatrizz[75][455] = 9'b111111111;
assign micromatrizz[75][456] = 9'b111111111;
assign micromatrizz[75][457] = 9'b111111111;
assign micromatrizz[75][458] = 9'b111111111;
assign micromatrizz[75][459] = 9'b111111111;
assign micromatrizz[75][460] = 9'b111111111;
assign micromatrizz[75][461] = 9'b111111111;
assign micromatrizz[75][462] = 9'b111111111;
assign micromatrizz[75][463] = 9'b111111111;
assign micromatrizz[75][464] = 9'b111111111;
assign micromatrizz[75][465] = 9'b111111111;
assign micromatrizz[75][466] = 9'b111111111;
assign micromatrizz[75][467] = 9'b111111111;
assign micromatrizz[75][468] = 9'b111111111;
assign micromatrizz[75][469] = 9'b111111111;
assign micromatrizz[75][470] = 9'b111111111;
assign micromatrizz[75][471] = 9'b111111111;
assign micromatrizz[75][472] = 9'b111111111;
assign micromatrizz[75][473] = 9'b111111111;
assign micromatrizz[75][474] = 9'b111111111;
assign micromatrizz[75][475] = 9'b111111111;
assign micromatrizz[75][476] = 9'b111111111;
assign micromatrizz[75][477] = 9'b111111111;
assign micromatrizz[75][478] = 9'b111111111;
assign micromatrizz[75][479] = 9'b111111111;
assign micromatrizz[75][480] = 9'b111111111;
assign micromatrizz[75][481] = 9'b111111111;
assign micromatrizz[75][482] = 9'b111111111;
assign micromatrizz[75][483] = 9'b111111111;
assign micromatrizz[75][484] = 9'b111111111;
assign micromatrizz[75][485] = 9'b111111111;
assign micromatrizz[75][486] = 9'b111111111;
assign micromatrizz[75][487] = 9'b111111111;
assign micromatrizz[75][488] = 9'b111111111;
assign micromatrizz[75][489] = 9'b111111111;
assign micromatrizz[75][490] = 9'b111111111;
assign micromatrizz[75][491] = 9'b111111111;
assign micromatrizz[75][492] = 9'b111111111;
assign micromatrizz[75][493] = 9'b111111111;
assign micromatrizz[75][494] = 9'b111111111;
assign micromatrizz[75][495] = 9'b111111111;
assign micromatrizz[75][496] = 9'b111111111;
assign micromatrizz[75][497] = 9'b111111111;
assign micromatrizz[75][498] = 9'b111111111;
assign micromatrizz[75][499] = 9'b111111111;
assign micromatrizz[75][500] = 9'b111111111;
assign micromatrizz[75][501] = 9'b111111111;
assign micromatrizz[75][502] = 9'b111111111;
assign micromatrizz[75][503] = 9'b111111111;
assign micromatrizz[75][504] = 9'b111111111;
assign micromatrizz[75][505] = 9'b111111111;
assign micromatrizz[75][506] = 9'b111111111;
assign micromatrizz[75][507] = 9'b111111111;
assign micromatrizz[75][508] = 9'b111111111;
assign micromatrizz[75][509] = 9'b111111111;
assign micromatrizz[75][510] = 9'b111111111;
assign micromatrizz[75][511] = 9'b111111111;
assign micromatrizz[75][512] = 9'b111111111;
assign micromatrizz[75][513] = 9'b111111111;
assign micromatrizz[75][514] = 9'b111111111;
assign micromatrizz[75][515] = 9'b111111111;
assign micromatrizz[75][516] = 9'b111111111;
assign micromatrizz[75][517] = 9'b111111111;
assign micromatrizz[75][518] = 9'b111111111;
assign micromatrizz[75][519] = 9'b111111111;
assign micromatrizz[75][520] = 9'b111111111;
assign micromatrizz[75][521] = 9'b111111111;
assign micromatrizz[75][522] = 9'b111111111;
assign micromatrizz[75][523] = 9'b111111111;
assign micromatrizz[75][524] = 9'b111111111;
assign micromatrizz[75][525] = 9'b111111111;
assign micromatrizz[75][526] = 9'b111111111;
assign micromatrizz[75][527] = 9'b111111111;
assign micromatrizz[75][528] = 9'b111111111;
assign micromatrizz[75][529] = 9'b111111111;
assign micromatrizz[75][530] = 9'b111111111;
assign micromatrizz[75][531] = 9'b111111111;
assign micromatrizz[75][532] = 9'b111111111;
assign micromatrizz[75][533] = 9'b111111111;
assign micromatrizz[75][534] = 9'b111111111;
assign micromatrizz[75][535] = 9'b111111111;
assign micromatrizz[75][536] = 9'b111111111;
assign micromatrizz[75][537] = 9'b111111111;
assign micromatrizz[75][538] = 9'b111111111;
assign micromatrizz[75][539] = 9'b111111111;
assign micromatrizz[75][540] = 9'b111111111;
assign micromatrizz[75][541] = 9'b111111111;
assign micromatrizz[75][542] = 9'b111111111;
assign micromatrizz[75][543] = 9'b111111111;
assign micromatrizz[75][544] = 9'b111111111;
assign micromatrizz[75][545] = 9'b111111111;
assign micromatrizz[75][546] = 9'b111111111;
assign micromatrizz[75][547] = 9'b111111111;
assign micromatrizz[75][548] = 9'b111111111;
assign micromatrizz[75][549] = 9'b111111111;
assign micromatrizz[75][550] = 9'b111111111;
assign micromatrizz[75][551] = 9'b111111111;
assign micromatrizz[75][552] = 9'b111111111;
assign micromatrizz[75][553] = 9'b111111111;
assign micromatrizz[75][554] = 9'b111111111;
assign micromatrizz[75][555] = 9'b111111111;
assign micromatrizz[75][556] = 9'b111111111;
assign micromatrizz[75][557] = 9'b111111111;
assign micromatrizz[75][558] = 9'b111111111;
assign micromatrizz[75][559] = 9'b111111111;
assign micromatrizz[75][560] = 9'b111111111;
assign micromatrizz[75][561] = 9'b111111111;
assign micromatrizz[75][562] = 9'b111111111;
assign micromatrizz[75][563] = 9'b111111111;
assign micromatrizz[75][564] = 9'b111111111;
assign micromatrizz[75][565] = 9'b111111111;
assign micromatrizz[75][566] = 9'b111111111;
assign micromatrizz[75][567] = 9'b111111111;
assign micromatrizz[75][568] = 9'b111111111;
assign micromatrizz[75][569] = 9'b111111111;
assign micromatrizz[75][570] = 9'b111111111;
assign micromatrizz[75][571] = 9'b111111111;
assign micromatrizz[75][572] = 9'b111111111;
assign micromatrizz[75][573] = 9'b111111111;
assign micromatrizz[75][574] = 9'b111111111;
assign micromatrizz[75][575] = 9'b111111111;
assign micromatrizz[75][576] = 9'b111111111;
assign micromatrizz[75][577] = 9'b111111111;
assign micromatrizz[75][578] = 9'b111111111;
assign micromatrizz[75][579] = 9'b111111111;
assign micromatrizz[75][580] = 9'b111111111;
assign micromatrizz[75][581] = 9'b111111111;
assign micromatrizz[75][582] = 9'b111111111;
assign micromatrizz[75][583] = 9'b111111111;
assign micromatrizz[75][584] = 9'b111111111;
assign micromatrizz[75][585] = 9'b111111111;
assign micromatrizz[75][586] = 9'b111111111;
assign micromatrizz[75][587] = 9'b111111111;
assign micromatrizz[75][588] = 9'b111111111;
assign micromatrizz[75][589] = 9'b111111111;
assign micromatrizz[75][590] = 9'b111111111;
assign micromatrizz[75][591] = 9'b111111111;
assign micromatrizz[75][592] = 9'b111111111;
assign micromatrizz[75][593] = 9'b111111111;
assign micromatrizz[75][594] = 9'b111111111;
assign micromatrizz[75][595] = 9'b111111111;
assign micromatrizz[75][596] = 9'b111111111;
assign micromatrizz[75][597] = 9'b111111111;
assign micromatrizz[75][598] = 9'b111111111;
assign micromatrizz[75][599] = 9'b111111111;
assign micromatrizz[75][600] = 9'b111111111;
assign micromatrizz[75][601] = 9'b111111111;
assign micromatrizz[75][602] = 9'b111111111;
assign micromatrizz[75][603] = 9'b111111111;
assign micromatrizz[75][604] = 9'b111111111;
assign micromatrizz[75][605] = 9'b111111111;
assign micromatrizz[75][606] = 9'b111111111;
assign micromatrizz[75][607] = 9'b111111111;
assign micromatrizz[75][608] = 9'b111111111;
assign micromatrizz[75][609] = 9'b111111111;
assign micromatrizz[75][610] = 9'b111111111;
assign micromatrizz[75][611] = 9'b111111111;
assign micromatrizz[75][612] = 9'b111111111;
assign micromatrizz[75][613] = 9'b111111111;
assign micromatrizz[75][614] = 9'b111111111;
assign micromatrizz[75][615] = 9'b111111111;
assign micromatrizz[75][616] = 9'b111111111;
assign micromatrizz[75][617] = 9'b111111111;
assign micromatrizz[75][618] = 9'b111111111;
assign micromatrizz[75][619] = 9'b111111111;
assign micromatrizz[75][620] = 9'b111111111;
assign micromatrizz[75][621] = 9'b111111111;
assign micromatrizz[75][622] = 9'b111111111;
assign micromatrizz[75][623] = 9'b111111111;
assign micromatrizz[75][624] = 9'b111111111;
assign micromatrizz[75][625] = 9'b111111111;
assign micromatrizz[75][626] = 9'b111111111;
assign micromatrizz[75][627] = 9'b111111111;
assign micromatrizz[75][628] = 9'b111111111;
assign micromatrizz[75][629] = 9'b111111111;
assign micromatrizz[75][630] = 9'b111111111;
assign micromatrizz[75][631] = 9'b111111111;
assign micromatrizz[75][632] = 9'b111111111;
assign micromatrizz[75][633] = 9'b111111111;
assign micromatrizz[75][634] = 9'b111111111;
assign micromatrizz[75][635] = 9'b111111111;
assign micromatrizz[75][636] = 9'b111111111;
assign micromatrizz[75][637] = 9'b111111111;
assign micromatrizz[75][638] = 9'b111111111;
assign micromatrizz[75][639] = 9'b111111111;
assign micromatrizz[76][0] = 9'b111111111;
assign micromatrizz[76][1] = 9'b111111111;
assign micromatrizz[76][2] = 9'b111111111;
assign micromatrizz[76][3] = 9'b111111111;
assign micromatrizz[76][4] = 9'b111111111;
assign micromatrizz[76][5] = 9'b111111111;
assign micromatrizz[76][6] = 9'b111111111;
assign micromatrizz[76][7] = 9'b111111111;
assign micromatrizz[76][8] = 9'b111111111;
assign micromatrizz[76][9] = 9'b111111111;
assign micromatrizz[76][10] = 9'b111111111;
assign micromatrizz[76][11] = 9'b111111111;
assign micromatrizz[76][12] = 9'b111111111;
assign micromatrizz[76][13] = 9'b111111111;
assign micromatrizz[76][14] = 9'b111111111;
assign micromatrizz[76][15] = 9'b111111111;
assign micromatrizz[76][16] = 9'b111111111;
assign micromatrizz[76][17] = 9'b111111111;
assign micromatrizz[76][18] = 9'b111111111;
assign micromatrizz[76][19] = 9'b111111111;
assign micromatrizz[76][20] = 9'b111111111;
assign micromatrizz[76][21] = 9'b111111111;
assign micromatrizz[76][22] = 9'b111111111;
assign micromatrizz[76][23] = 9'b111111111;
assign micromatrizz[76][24] = 9'b111111111;
assign micromatrizz[76][25] = 9'b111111111;
assign micromatrizz[76][26] = 9'b111111111;
assign micromatrizz[76][27] = 9'b111111111;
assign micromatrizz[76][28] = 9'b111111111;
assign micromatrizz[76][29] = 9'b111111111;
assign micromatrizz[76][30] = 9'b111111111;
assign micromatrizz[76][31] = 9'b111111111;
assign micromatrizz[76][32] = 9'b111111111;
assign micromatrizz[76][33] = 9'b111111111;
assign micromatrizz[76][34] = 9'b111111111;
assign micromatrizz[76][35] = 9'b111111111;
assign micromatrizz[76][36] = 9'b111111111;
assign micromatrizz[76][37] = 9'b111111111;
assign micromatrizz[76][38] = 9'b111111111;
assign micromatrizz[76][39] = 9'b111111111;
assign micromatrizz[76][40] = 9'b111111111;
assign micromatrizz[76][41] = 9'b111111111;
assign micromatrizz[76][42] = 9'b111111111;
assign micromatrizz[76][43] = 9'b111111111;
assign micromatrizz[76][44] = 9'b111111111;
assign micromatrizz[76][45] = 9'b111111111;
assign micromatrizz[76][46] = 9'b111111111;
assign micromatrizz[76][47] = 9'b111111111;
assign micromatrizz[76][48] = 9'b111111111;
assign micromatrizz[76][49] = 9'b111111111;
assign micromatrizz[76][50] = 9'b111111111;
assign micromatrizz[76][51] = 9'b111111111;
assign micromatrizz[76][52] = 9'b111111111;
assign micromatrizz[76][53] = 9'b111111111;
assign micromatrizz[76][54] = 9'b111111111;
assign micromatrizz[76][55] = 9'b111111111;
assign micromatrizz[76][56] = 9'b111111111;
assign micromatrizz[76][57] = 9'b111111111;
assign micromatrizz[76][58] = 9'b111111111;
assign micromatrizz[76][59] = 9'b111111111;
assign micromatrizz[76][60] = 9'b111111111;
assign micromatrizz[76][61] = 9'b111111111;
assign micromatrizz[76][62] = 9'b111111111;
assign micromatrizz[76][63] = 9'b111111111;
assign micromatrizz[76][64] = 9'b111111111;
assign micromatrizz[76][65] = 9'b111111111;
assign micromatrizz[76][66] = 9'b111111111;
assign micromatrizz[76][67] = 9'b111111111;
assign micromatrizz[76][68] = 9'b111111111;
assign micromatrizz[76][69] = 9'b111111111;
assign micromatrizz[76][70] = 9'b111111111;
assign micromatrizz[76][71] = 9'b111111111;
assign micromatrizz[76][72] = 9'b111111111;
assign micromatrizz[76][73] = 9'b111111111;
assign micromatrizz[76][74] = 9'b111111111;
assign micromatrizz[76][75] = 9'b111111111;
assign micromatrizz[76][76] = 9'b111111111;
assign micromatrizz[76][77] = 9'b111111111;
assign micromatrizz[76][78] = 9'b111111111;
assign micromatrizz[76][79] = 9'b111111111;
assign micromatrizz[76][80] = 9'b111111111;
assign micromatrizz[76][81] = 9'b111111111;
assign micromatrizz[76][82] = 9'b111111111;
assign micromatrizz[76][83] = 9'b111111111;
assign micromatrizz[76][84] = 9'b111111111;
assign micromatrizz[76][85] = 9'b111111111;
assign micromatrizz[76][86] = 9'b111111111;
assign micromatrizz[76][87] = 9'b111111111;
assign micromatrizz[76][88] = 9'b111111111;
assign micromatrizz[76][89] = 9'b111111111;
assign micromatrizz[76][90] = 9'b111111111;
assign micromatrizz[76][91] = 9'b111111111;
assign micromatrizz[76][92] = 9'b111111111;
assign micromatrizz[76][93] = 9'b111111111;
assign micromatrizz[76][94] = 9'b111111111;
assign micromatrizz[76][95] = 9'b111111111;
assign micromatrizz[76][96] = 9'b111111111;
assign micromatrizz[76][97] = 9'b111111111;
assign micromatrizz[76][98] = 9'b111111111;
assign micromatrizz[76][99] = 9'b111111111;
assign micromatrizz[76][100] = 9'b111111111;
assign micromatrizz[76][101] = 9'b111111111;
assign micromatrizz[76][102] = 9'b111111111;
assign micromatrizz[76][103] = 9'b111111111;
assign micromatrizz[76][104] = 9'b111111111;
assign micromatrizz[76][105] = 9'b111111111;
assign micromatrizz[76][106] = 9'b111111111;
assign micromatrizz[76][107] = 9'b111111111;
assign micromatrizz[76][108] = 9'b111111111;
assign micromatrizz[76][109] = 9'b111111111;
assign micromatrizz[76][110] = 9'b111111111;
assign micromatrizz[76][111] = 9'b111111111;
assign micromatrizz[76][112] = 9'b111111111;
assign micromatrizz[76][113] = 9'b111111111;
assign micromatrizz[76][114] = 9'b111111111;
assign micromatrizz[76][115] = 9'b111111111;
assign micromatrizz[76][116] = 9'b111111111;
assign micromatrizz[76][117] = 9'b111111111;
assign micromatrizz[76][118] = 9'b111111111;
assign micromatrizz[76][119] = 9'b111111111;
assign micromatrizz[76][120] = 9'b111111111;
assign micromatrizz[76][121] = 9'b111111111;
assign micromatrizz[76][122] = 9'b111111111;
assign micromatrizz[76][123] = 9'b111111111;
assign micromatrizz[76][124] = 9'b111111111;
assign micromatrizz[76][125] = 9'b111111111;
assign micromatrizz[76][126] = 9'b111111111;
assign micromatrizz[76][127] = 9'b111111111;
assign micromatrizz[76][128] = 9'b111111111;
assign micromatrizz[76][129] = 9'b111111111;
assign micromatrizz[76][130] = 9'b111111111;
assign micromatrizz[76][131] = 9'b111111111;
assign micromatrizz[76][132] = 9'b111111111;
assign micromatrizz[76][133] = 9'b111111111;
assign micromatrizz[76][134] = 9'b111111111;
assign micromatrizz[76][135] = 9'b111111111;
assign micromatrizz[76][136] = 9'b111111111;
assign micromatrizz[76][137] = 9'b111111111;
assign micromatrizz[76][138] = 9'b111111111;
assign micromatrizz[76][139] = 9'b111111111;
assign micromatrizz[76][140] = 9'b111111111;
assign micromatrizz[76][141] = 9'b111111111;
assign micromatrizz[76][142] = 9'b111111111;
assign micromatrizz[76][143] = 9'b111111111;
assign micromatrizz[76][144] = 9'b111111111;
assign micromatrizz[76][145] = 9'b111111111;
assign micromatrizz[76][146] = 9'b111111111;
assign micromatrizz[76][147] = 9'b111111111;
assign micromatrizz[76][148] = 9'b111111111;
assign micromatrizz[76][149] = 9'b111111111;
assign micromatrizz[76][150] = 9'b111111111;
assign micromatrizz[76][151] = 9'b111111111;
assign micromatrizz[76][152] = 9'b111111111;
assign micromatrizz[76][153] = 9'b111111111;
assign micromatrizz[76][154] = 9'b111111111;
assign micromatrizz[76][155] = 9'b111111111;
assign micromatrizz[76][156] = 9'b111111111;
assign micromatrizz[76][157] = 9'b111111111;
assign micromatrizz[76][158] = 9'b111111111;
assign micromatrizz[76][159] = 9'b111111111;
assign micromatrizz[76][160] = 9'b111111111;
assign micromatrizz[76][161] = 9'b111111111;
assign micromatrizz[76][162] = 9'b111111111;
assign micromatrizz[76][163] = 9'b111111111;
assign micromatrizz[76][164] = 9'b111111111;
assign micromatrizz[76][165] = 9'b111111111;
assign micromatrizz[76][166] = 9'b111111111;
assign micromatrizz[76][167] = 9'b111111111;
assign micromatrizz[76][168] = 9'b111111111;
assign micromatrizz[76][169] = 9'b111111111;
assign micromatrizz[76][170] = 9'b111111111;
assign micromatrizz[76][171] = 9'b111111111;
assign micromatrizz[76][172] = 9'b111111111;
assign micromatrizz[76][173] = 9'b111111111;
assign micromatrizz[76][174] = 9'b111111111;
assign micromatrizz[76][175] = 9'b111111111;
assign micromatrizz[76][176] = 9'b111111111;
assign micromatrizz[76][177] = 9'b111111111;
assign micromatrizz[76][178] = 9'b111111111;
assign micromatrizz[76][179] = 9'b111111111;
assign micromatrizz[76][180] = 9'b111111111;
assign micromatrizz[76][181] = 9'b111111111;
assign micromatrizz[76][182] = 9'b111111111;
assign micromatrizz[76][183] = 9'b111111111;
assign micromatrizz[76][184] = 9'b111111111;
assign micromatrizz[76][185] = 9'b111111111;
assign micromatrizz[76][186] = 9'b111111111;
assign micromatrizz[76][187] = 9'b111111111;
assign micromatrizz[76][188] = 9'b111111111;
assign micromatrizz[76][189] = 9'b111111111;
assign micromatrizz[76][190] = 9'b111111111;
assign micromatrizz[76][191] = 9'b111111111;
assign micromatrizz[76][192] = 9'b111111111;
assign micromatrizz[76][193] = 9'b111111111;
assign micromatrizz[76][194] = 9'b111111111;
assign micromatrizz[76][195] = 9'b111111111;
assign micromatrizz[76][196] = 9'b111111111;
assign micromatrizz[76][197] = 9'b111111111;
assign micromatrizz[76][198] = 9'b111111111;
assign micromatrizz[76][199] = 9'b111111111;
assign micromatrizz[76][200] = 9'b111111111;
assign micromatrizz[76][201] = 9'b111111111;
assign micromatrizz[76][202] = 9'b111111111;
assign micromatrizz[76][203] = 9'b111111111;
assign micromatrizz[76][204] = 9'b111111111;
assign micromatrizz[76][205] = 9'b111111111;
assign micromatrizz[76][206] = 9'b111111111;
assign micromatrizz[76][207] = 9'b111111111;
assign micromatrizz[76][208] = 9'b111111111;
assign micromatrizz[76][209] = 9'b111111111;
assign micromatrizz[76][210] = 9'b111111111;
assign micromatrizz[76][211] = 9'b111111111;
assign micromatrizz[76][212] = 9'b111111111;
assign micromatrizz[76][213] = 9'b111111111;
assign micromatrizz[76][214] = 9'b111111111;
assign micromatrizz[76][215] = 9'b111111111;
assign micromatrizz[76][216] = 9'b111111111;
assign micromatrizz[76][217] = 9'b111111111;
assign micromatrizz[76][218] = 9'b111111111;
assign micromatrizz[76][219] = 9'b111111111;
assign micromatrizz[76][220] = 9'b111111111;
assign micromatrizz[76][221] = 9'b111111111;
assign micromatrizz[76][222] = 9'b111111111;
assign micromatrizz[76][223] = 9'b111111111;
assign micromatrizz[76][224] = 9'b111111111;
assign micromatrizz[76][225] = 9'b111111111;
assign micromatrizz[76][226] = 9'b111111111;
assign micromatrizz[76][227] = 9'b111111111;
assign micromatrizz[76][228] = 9'b111111111;
assign micromatrizz[76][229] = 9'b111111111;
assign micromatrizz[76][230] = 9'b111111111;
assign micromatrizz[76][231] = 9'b111111111;
assign micromatrizz[76][232] = 9'b111111111;
assign micromatrizz[76][233] = 9'b111111111;
assign micromatrizz[76][234] = 9'b111111111;
assign micromatrizz[76][235] = 9'b111111111;
assign micromatrizz[76][236] = 9'b111111111;
assign micromatrizz[76][237] = 9'b111111111;
assign micromatrizz[76][238] = 9'b111111111;
assign micromatrizz[76][239] = 9'b111111111;
assign micromatrizz[76][240] = 9'b111111111;
assign micromatrizz[76][241] = 9'b111111111;
assign micromatrizz[76][242] = 9'b111111111;
assign micromatrizz[76][243] = 9'b111111111;
assign micromatrizz[76][244] = 9'b111111111;
assign micromatrizz[76][245] = 9'b111111111;
assign micromatrizz[76][246] = 9'b111111111;
assign micromatrizz[76][247] = 9'b111111111;
assign micromatrizz[76][248] = 9'b111111111;
assign micromatrizz[76][249] = 9'b111111111;
assign micromatrizz[76][250] = 9'b111111111;
assign micromatrizz[76][251] = 9'b111111111;
assign micromatrizz[76][252] = 9'b111111111;
assign micromatrizz[76][253] = 9'b111111111;
assign micromatrizz[76][254] = 9'b111111111;
assign micromatrizz[76][255] = 9'b111111111;
assign micromatrizz[76][256] = 9'b111111111;
assign micromatrizz[76][257] = 9'b111111111;
assign micromatrizz[76][258] = 9'b111111111;
assign micromatrizz[76][259] = 9'b111111111;
assign micromatrizz[76][260] = 9'b111111111;
assign micromatrizz[76][261] = 9'b111111111;
assign micromatrizz[76][262] = 9'b111111111;
assign micromatrizz[76][263] = 9'b111111111;
assign micromatrizz[76][264] = 9'b111111111;
assign micromatrizz[76][265] = 9'b111111111;
assign micromatrizz[76][266] = 9'b111111111;
assign micromatrizz[76][267] = 9'b111111111;
assign micromatrizz[76][268] = 9'b111111111;
assign micromatrizz[76][269] = 9'b111111111;
assign micromatrizz[76][270] = 9'b111111111;
assign micromatrizz[76][271] = 9'b111111111;
assign micromatrizz[76][272] = 9'b111111111;
assign micromatrizz[76][273] = 9'b111111111;
assign micromatrizz[76][274] = 9'b111111111;
assign micromatrizz[76][275] = 9'b111111111;
assign micromatrizz[76][276] = 9'b111111111;
assign micromatrizz[76][277] = 9'b111111111;
assign micromatrizz[76][278] = 9'b111111111;
assign micromatrizz[76][279] = 9'b111111111;
assign micromatrizz[76][280] = 9'b111111111;
assign micromatrizz[76][281] = 9'b111111111;
assign micromatrizz[76][282] = 9'b111111111;
assign micromatrizz[76][283] = 9'b111111111;
assign micromatrizz[76][284] = 9'b111111111;
assign micromatrizz[76][285] = 9'b111111111;
assign micromatrizz[76][286] = 9'b111111111;
assign micromatrizz[76][287] = 9'b111111111;
assign micromatrizz[76][288] = 9'b111111111;
assign micromatrizz[76][289] = 9'b111111111;
assign micromatrizz[76][290] = 9'b111111111;
assign micromatrizz[76][291] = 9'b111111111;
assign micromatrizz[76][292] = 9'b111111111;
assign micromatrizz[76][293] = 9'b111111111;
assign micromatrizz[76][294] = 9'b111111111;
assign micromatrizz[76][295] = 9'b111111111;
assign micromatrizz[76][296] = 9'b111111111;
assign micromatrizz[76][297] = 9'b111111111;
assign micromatrizz[76][298] = 9'b111111111;
assign micromatrizz[76][299] = 9'b111111111;
assign micromatrizz[76][300] = 9'b111111111;
assign micromatrizz[76][301] = 9'b111111111;
assign micromatrizz[76][302] = 9'b111111111;
assign micromatrizz[76][303] = 9'b111111111;
assign micromatrizz[76][304] = 9'b111111111;
assign micromatrizz[76][305] = 9'b111111111;
assign micromatrizz[76][306] = 9'b111111111;
assign micromatrizz[76][307] = 9'b111111111;
assign micromatrizz[76][308] = 9'b111111111;
assign micromatrizz[76][309] = 9'b111111111;
assign micromatrizz[76][310] = 9'b111111111;
assign micromatrizz[76][311] = 9'b111111111;
assign micromatrizz[76][312] = 9'b111111111;
assign micromatrizz[76][313] = 9'b111111111;
assign micromatrizz[76][314] = 9'b111111111;
assign micromatrizz[76][315] = 9'b111111111;
assign micromatrizz[76][316] = 9'b111111111;
assign micromatrizz[76][317] = 9'b111111111;
assign micromatrizz[76][318] = 9'b111111111;
assign micromatrizz[76][319] = 9'b111111111;
assign micromatrizz[76][320] = 9'b111111111;
assign micromatrizz[76][321] = 9'b111111111;
assign micromatrizz[76][322] = 9'b111111111;
assign micromatrizz[76][323] = 9'b111111111;
assign micromatrizz[76][324] = 9'b111111111;
assign micromatrizz[76][325] = 9'b111111111;
assign micromatrizz[76][326] = 9'b111111111;
assign micromatrizz[76][327] = 9'b111111111;
assign micromatrizz[76][328] = 9'b111111111;
assign micromatrizz[76][329] = 9'b111111111;
assign micromatrizz[76][330] = 9'b111111111;
assign micromatrizz[76][331] = 9'b111111111;
assign micromatrizz[76][332] = 9'b111111111;
assign micromatrizz[76][333] = 9'b111111111;
assign micromatrizz[76][334] = 9'b111111111;
assign micromatrizz[76][335] = 9'b111111111;
assign micromatrizz[76][336] = 9'b111111111;
assign micromatrizz[76][337] = 9'b111111111;
assign micromatrizz[76][338] = 9'b111111111;
assign micromatrizz[76][339] = 9'b111111111;
assign micromatrizz[76][340] = 9'b111111111;
assign micromatrizz[76][341] = 9'b111111111;
assign micromatrizz[76][342] = 9'b111111111;
assign micromatrizz[76][343] = 9'b111111111;
assign micromatrizz[76][344] = 9'b111111111;
assign micromatrizz[76][345] = 9'b111111111;
assign micromatrizz[76][346] = 9'b111111111;
assign micromatrizz[76][347] = 9'b111111111;
assign micromatrizz[76][348] = 9'b111111111;
assign micromatrizz[76][349] = 9'b111111111;
assign micromatrizz[76][350] = 9'b111111111;
assign micromatrizz[76][351] = 9'b111111111;
assign micromatrizz[76][352] = 9'b111111111;
assign micromatrizz[76][353] = 9'b111111111;
assign micromatrizz[76][354] = 9'b111111111;
assign micromatrizz[76][355] = 9'b111111111;
assign micromatrizz[76][356] = 9'b111111111;
assign micromatrizz[76][357] = 9'b111111111;
assign micromatrizz[76][358] = 9'b111111111;
assign micromatrizz[76][359] = 9'b111111111;
assign micromatrizz[76][360] = 9'b111111111;
assign micromatrizz[76][361] = 9'b111111111;
assign micromatrizz[76][362] = 9'b111111111;
assign micromatrizz[76][363] = 9'b111111111;
assign micromatrizz[76][364] = 9'b111111111;
assign micromatrizz[76][365] = 9'b111111111;
assign micromatrizz[76][366] = 9'b111111111;
assign micromatrizz[76][367] = 9'b111111111;
assign micromatrizz[76][368] = 9'b111111111;
assign micromatrizz[76][369] = 9'b111111111;
assign micromatrizz[76][370] = 9'b111111111;
assign micromatrizz[76][371] = 9'b111111111;
assign micromatrizz[76][372] = 9'b111111111;
assign micromatrizz[76][373] = 9'b111111111;
assign micromatrizz[76][374] = 9'b111111111;
assign micromatrizz[76][375] = 9'b111111111;
assign micromatrizz[76][376] = 9'b111111111;
assign micromatrizz[76][377] = 9'b111111111;
assign micromatrizz[76][378] = 9'b111111111;
assign micromatrizz[76][379] = 9'b111111111;
assign micromatrizz[76][380] = 9'b111111111;
assign micromatrizz[76][381] = 9'b111111111;
assign micromatrizz[76][382] = 9'b111111111;
assign micromatrizz[76][383] = 9'b111111111;
assign micromatrizz[76][384] = 9'b111111111;
assign micromatrizz[76][385] = 9'b111111111;
assign micromatrizz[76][386] = 9'b111111111;
assign micromatrizz[76][387] = 9'b111111111;
assign micromatrizz[76][388] = 9'b111111111;
assign micromatrizz[76][389] = 9'b111111111;
assign micromatrizz[76][390] = 9'b111111111;
assign micromatrizz[76][391] = 9'b111111111;
assign micromatrizz[76][392] = 9'b111111111;
assign micromatrizz[76][393] = 9'b111111111;
assign micromatrizz[76][394] = 9'b111111111;
assign micromatrizz[76][395] = 9'b111111111;
assign micromatrizz[76][396] = 9'b111111111;
assign micromatrizz[76][397] = 9'b111111111;
assign micromatrizz[76][398] = 9'b111111111;
assign micromatrizz[76][399] = 9'b111111111;
assign micromatrizz[76][400] = 9'b111111111;
assign micromatrizz[76][401] = 9'b111111111;
assign micromatrizz[76][402] = 9'b111111111;
assign micromatrizz[76][403] = 9'b111111111;
assign micromatrizz[76][404] = 9'b111111111;
assign micromatrizz[76][405] = 9'b111111111;
assign micromatrizz[76][406] = 9'b111111111;
assign micromatrizz[76][407] = 9'b111111111;
assign micromatrizz[76][408] = 9'b111111111;
assign micromatrizz[76][409] = 9'b111111111;
assign micromatrizz[76][410] = 9'b111111111;
assign micromatrizz[76][411] = 9'b111111111;
assign micromatrizz[76][412] = 9'b111111111;
assign micromatrizz[76][413] = 9'b111111111;
assign micromatrizz[76][414] = 9'b111111111;
assign micromatrizz[76][415] = 9'b111111111;
assign micromatrizz[76][416] = 9'b111111111;
assign micromatrizz[76][417] = 9'b111111111;
assign micromatrizz[76][418] = 9'b111111111;
assign micromatrizz[76][419] = 9'b111111111;
assign micromatrizz[76][420] = 9'b111111111;
assign micromatrizz[76][421] = 9'b111111111;
assign micromatrizz[76][422] = 9'b111111111;
assign micromatrizz[76][423] = 9'b111111111;
assign micromatrizz[76][424] = 9'b111111111;
assign micromatrizz[76][425] = 9'b111111111;
assign micromatrizz[76][426] = 9'b111111111;
assign micromatrizz[76][427] = 9'b111111111;
assign micromatrizz[76][428] = 9'b111111111;
assign micromatrizz[76][429] = 9'b111111111;
assign micromatrizz[76][430] = 9'b111111111;
assign micromatrizz[76][431] = 9'b111111111;
assign micromatrizz[76][432] = 9'b111111111;
assign micromatrizz[76][433] = 9'b111111111;
assign micromatrizz[76][434] = 9'b111111111;
assign micromatrizz[76][435] = 9'b111111111;
assign micromatrizz[76][436] = 9'b111111111;
assign micromatrizz[76][437] = 9'b111111111;
assign micromatrizz[76][438] = 9'b111111111;
assign micromatrizz[76][439] = 9'b111111111;
assign micromatrizz[76][440] = 9'b111111111;
assign micromatrizz[76][441] = 9'b111111111;
assign micromatrizz[76][442] = 9'b111111111;
assign micromatrizz[76][443] = 9'b111111111;
assign micromatrizz[76][444] = 9'b111111111;
assign micromatrizz[76][445] = 9'b111111111;
assign micromatrizz[76][446] = 9'b111111111;
assign micromatrizz[76][447] = 9'b111111111;
assign micromatrizz[76][448] = 9'b111111111;
assign micromatrizz[76][449] = 9'b111111111;
assign micromatrizz[76][450] = 9'b111111111;
assign micromatrizz[76][451] = 9'b111111111;
assign micromatrizz[76][452] = 9'b111111111;
assign micromatrizz[76][453] = 9'b111111111;
assign micromatrizz[76][454] = 9'b111111111;
assign micromatrizz[76][455] = 9'b111111111;
assign micromatrizz[76][456] = 9'b111111111;
assign micromatrizz[76][457] = 9'b111111111;
assign micromatrizz[76][458] = 9'b111111111;
assign micromatrizz[76][459] = 9'b111111111;
assign micromatrizz[76][460] = 9'b111111111;
assign micromatrizz[76][461] = 9'b111111111;
assign micromatrizz[76][462] = 9'b111111111;
assign micromatrizz[76][463] = 9'b111111111;
assign micromatrizz[76][464] = 9'b111111111;
assign micromatrizz[76][465] = 9'b111111111;
assign micromatrizz[76][466] = 9'b111111111;
assign micromatrizz[76][467] = 9'b111111111;
assign micromatrizz[76][468] = 9'b111111111;
assign micromatrizz[76][469] = 9'b111111111;
assign micromatrizz[76][470] = 9'b111111111;
assign micromatrizz[76][471] = 9'b111111111;
assign micromatrizz[76][472] = 9'b111111111;
assign micromatrizz[76][473] = 9'b111111111;
assign micromatrizz[76][474] = 9'b111111111;
assign micromatrizz[76][475] = 9'b111111111;
assign micromatrizz[76][476] = 9'b111111111;
assign micromatrizz[76][477] = 9'b111111111;
assign micromatrizz[76][478] = 9'b111111111;
assign micromatrizz[76][479] = 9'b111111111;
assign micromatrizz[76][480] = 9'b111111111;
assign micromatrizz[76][481] = 9'b111111111;
assign micromatrizz[76][482] = 9'b111111111;
assign micromatrizz[76][483] = 9'b111111111;
assign micromatrizz[76][484] = 9'b111111111;
assign micromatrizz[76][485] = 9'b111111111;
assign micromatrizz[76][486] = 9'b111111111;
assign micromatrizz[76][487] = 9'b111111111;
assign micromatrizz[76][488] = 9'b111111111;
assign micromatrizz[76][489] = 9'b111111111;
assign micromatrizz[76][490] = 9'b111111111;
assign micromatrizz[76][491] = 9'b111111111;
assign micromatrizz[76][492] = 9'b111111111;
assign micromatrizz[76][493] = 9'b111111111;
assign micromatrizz[76][494] = 9'b111111111;
assign micromatrizz[76][495] = 9'b111111111;
assign micromatrizz[76][496] = 9'b111111111;
assign micromatrizz[76][497] = 9'b111111111;
assign micromatrizz[76][498] = 9'b111111111;
assign micromatrizz[76][499] = 9'b111111111;
assign micromatrizz[76][500] = 9'b111111111;
assign micromatrizz[76][501] = 9'b111111111;
assign micromatrizz[76][502] = 9'b111111111;
assign micromatrizz[76][503] = 9'b111111111;
assign micromatrizz[76][504] = 9'b111111111;
assign micromatrizz[76][505] = 9'b111111111;
assign micromatrizz[76][506] = 9'b111111111;
assign micromatrizz[76][507] = 9'b111111111;
assign micromatrizz[76][508] = 9'b111111111;
assign micromatrizz[76][509] = 9'b111111111;
assign micromatrizz[76][510] = 9'b111111111;
assign micromatrizz[76][511] = 9'b111111111;
assign micromatrizz[76][512] = 9'b111111111;
assign micromatrizz[76][513] = 9'b111111111;
assign micromatrizz[76][514] = 9'b111111111;
assign micromatrizz[76][515] = 9'b111111111;
assign micromatrizz[76][516] = 9'b111111111;
assign micromatrizz[76][517] = 9'b111111111;
assign micromatrizz[76][518] = 9'b111111111;
assign micromatrizz[76][519] = 9'b111111111;
assign micromatrizz[76][520] = 9'b111111111;
assign micromatrizz[76][521] = 9'b111111111;
assign micromatrizz[76][522] = 9'b111111111;
assign micromatrizz[76][523] = 9'b111111111;
assign micromatrizz[76][524] = 9'b111111111;
assign micromatrizz[76][525] = 9'b111111111;
assign micromatrizz[76][526] = 9'b111111111;
assign micromatrizz[76][527] = 9'b111111111;
assign micromatrizz[76][528] = 9'b111111111;
assign micromatrizz[76][529] = 9'b111111111;
assign micromatrizz[76][530] = 9'b111111111;
assign micromatrizz[76][531] = 9'b111111111;
assign micromatrizz[76][532] = 9'b111111111;
assign micromatrizz[76][533] = 9'b111111111;
assign micromatrizz[76][534] = 9'b111111111;
assign micromatrizz[76][535] = 9'b111111111;
assign micromatrizz[76][536] = 9'b111111111;
assign micromatrizz[76][537] = 9'b111111111;
assign micromatrizz[76][538] = 9'b111111111;
assign micromatrizz[76][539] = 9'b111111111;
assign micromatrizz[76][540] = 9'b111111111;
assign micromatrizz[76][541] = 9'b111111111;
assign micromatrizz[76][542] = 9'b111111111;
assign micromatrizz[76][543] = 9'b111111111;
assign micromatrizz[76][544] = 9'b111111111;
assign micromatrizz[76][545] = 9'b111111111;
assign micromatrizz[76][546] = 9'b111111111;
assign micromatrizz[76][547] = 9'b111111111;
assign micromatrizz[76][548] = 9'b111111111;
assign micromatrizz[76][549] = 9'b111111111;
assign micromatrizz[76][550] = 9'b111111111;
assign micromatrizz[76][551] = 9'b111111111;
assign micromatrizz[76][552] = 9'b111111111;
assign micromatrizz[76][553] = 9'b111111111;
assign micromatrizz[76][554] = 9'b111111111;
assign micromatrizz[76][555] = 9'b111111111;
assign micromatrizz[76][556] = 9'b111111111;
assign micromatrizz[76][557] = 9'b111111111;
assign micromatrizz[76][558] = 9'b111111111;
assign micromatrizz[76][559] = 9'b111111111;
assign micromatrizz[76][560] = 9'b111111111;
assign micromatrizz[76][561] = 9'b111111111;
assign micromatrizz[76][562] = 9'b111111111;
assign micromatrizz[76][563] = 9'b111111111;
assign micromatrizz[76][564] = 9'b111111111;
assign micromatrizz[76][565] = 9'b111111111;
assign micromatrizz[76][566] = 9'b111111111;
assign micromatrizz[76][567] = 9'b111111111;
assign micromatrizz[76][568] = 9'b111111111;
assign micromatrizz[76][569] = 9'b111111111;
assign micromatrizz[76][570] = 9'b111111111;
assign micromatrizz[76][571] = 9'b111111111;
assign micromatrizz[76][572] = 9'b111111111;
assign micromatrizz[76][573] = 9'b111111111;
assign micromatrizz[76][574] = 9'b111111111;
assign micromatrizz[76][575] = 9'b111111111;
assign micromatrizz[76][576] = 9'b111111111;
assign micromatrizz[76][577] = 9'b111111111;
assign micromatrizz[76][578] = 9'b111111111;
assign micromatrizz[76][579] = 9'b111111111;
assign micromatrizz[76][580] = 9'b111111111;
assign micromatrizz[76][581] = 9'b111111111;
assign micromatrizz[76][582] = 9'b111111111;
assign micromatrizz[76][583] = 9'b111111111;
assign micromatrizz[76][584] = 9'b111111111;
assign micromatrizz[76][585] = 9'b111111111;
assign micromatrizz[76][586] = 9'b111111111;
assign micromatrizz[76][587] = 9'b111111111;
assign micromatrizz[76][588] = 9'b111111111;
assign micromatrizz[76][589] = 9'b111111111;
assign micromatrizz[76][590] = 9'b111111111;
assign micromatrizz[76][591] = 9'b111111111;
assign micromatrizz[76][592] = 9'b111111111;
assign micromatrizz[76][593] = 9'b111111111;
assign micromatrizz[76][594] = 9'b111111111;
assign micromatrizz[76][595] = 9'b111111111;
assign micromatrizz[76][596] = 9'b111111111;
assign micromatrizz[76][597] = 9'b111111111;
assign micromatrizz[76][598] = 9'b111111111;
assign micromatrizz[76][599] = 9'b111111111;
assign micromatrizz[76][600] = 9'b111111111;
assign micromatrizz[76][601] = 9'b111111111;
assign micromatrizz[76][602] = 9'b111111111;
assign micromatrizz[76][603] = 9'b111111111;
assign micromatrizz[76][604] = 9'b111111111;
assign micromatrizz[76][605] = 9'b111111111;
assign micromatrizz[76][606] = 9'b111111111;
assign micromatrizz[76][607] = 9'b111111111;
assign micromatrizz[76][608] = 9'b111111111;
assign micromatrizz[76][609] = 9'b111111111;
assign micromatrizz[76][610] = 9'b111111111;
assign micromatrizz[76][611] = 9'b111111111;
assign micromatrizz[76][612] = 9'b111111111;
assign micromatrizz[76][613] = 9'b111111111;
assign micromatrizz[76][614] = 9'b111111111;
assign micromatrizz[76][615] = 9'b111111111;
assign micromatrizz[76][616] = 9'b111111111;
assign micromatrizz[76][617] = 9'b111111111;
assign micromatrizz[76][618] = 9'b111111111;
assign micromatrizz[76][619] = 9'b111111111;
assign micromatrizz[76][620] = 9'b111111111;
assign micromatrizz[76][621] = 9'b111111111;
assign micromatrizz[76][622] = 9'b111111111;
assign micromatrizz[76][623] = 9'b111111111;
assign micromatrizz[76][624] = 9'b111111111;
assign micromatrizz[76][625] = 9'b111111111;
assign micromatrizz[76][626] = 9'b111111111;
assign micromatrizz[76][627] = 9'b111111111;
assign micromatrizz[76][628] = 9'b111111111;
assign micromatrizz[76][629] = 9'b111111111;
assign micromatrizz[76][630] = 9'b111111111;
assign micromatrizz[76][631] = 9'b111111111;
assign micromatrizz[76][632] = 9'b111111111;
assign micromatrizz[76][633] = 9'b111111111;
assign micromatrizz[76][634] = 9'b111111111;
assign micromatrizz[76][635] = 9'b111111111;
assign micromatrizz[76][636] = 9'b111111111;
assign micromatrizz[76][637] = 9'b111111111;
assign micromatrizz[76][638] = 9'b111111111;
assign micromatrizz[76][639] = 9'b111111111;
assign micromatrizz[77][0] = 9'b111111111;
assign micromatrizz[77][1] = 9'b111111111;
assign micromatrizz[77][2] = 9'b111111111;
assign micromatrizz[77][3] = 9'b111111111;
assign micromatrizz[77][4] = 9'b111111111;
assign micromatrizz[77][5] = 9'b111111111;
assign micromatrizz[77][6] = 9'b111111111;
assign micromatrizz[77][7] = 9'b111111111;
assign micromatrizz[77][8] = 9'b111111111;
assign micromatrizz[77][9] = 9'b111111111;
assign micromatrizz[77][10] = 9'b111111111;
assign micromatrizz[77][11] = 9'b111111111;
assign micromatrizz[77][12] = 9'b111111111;
assign micromatrizz[77][13] = 9'b111111111;
assign micromatrizz[77][14] = 9'b111111111;
assign micromatrizz[77][15] = 9'b111111111;
assign micromatrizz[77][16] = 9'b111111111;
assign micromatrizz[77][17] = 9'b111111111;
assign micromatrizz[77][18] = 9'b111111111;
assign micromatrizz[77][19] = 9'b111111111;
assign micromatrizz[77][20] = 9'b111111111;
assign micromatrizz[77][21] = 9'b111111111;
assign micromatrizz[77][22] = 9'b111111111;
assign micromatrizz[77][23] = 9'b111111111;
assign micromatrizz[77][24] = 9'b111111111;
assign micromatrizz[77][25] = 9'b111111111;
assign micromatrizz[77][26] = 9'b111111111;
assign micromatrizz[77][27] = 9'b111111111;
assign micromatrizz[77][28] = 9'b111111111;
assign micromatrizz[77][29] = 9'b111111111;
assign micromatrizz[77][30] = 9'b111111111;
assign micromatrizz[77][31] = 9'b111111111;
assign micromatrizz[77][32] = 9'b111111111;
assign micromatrizz[77][33] = 9'b111111111;
assign micromatrizz[77][34] = 9'b111111111;
assign micromatrizz[77][35] = 9'b111111111;
assign micromatrizz[77][36] = 9'b111111111;
assign micromatrizz[77][37] = 9'b111111111;
assign micromatrizz[77][38] = 9'b111111111;
assign micromatrizz[77][39] = 9'b111111111;
assign micromatrizz[77][40] = 9'b111111111;
assign micromatrizz[77][41] = 9'b111111111;
assign micromatrizz[77][42] = 9'b111111111;
assign micromatrizz[77][43] = 9'b111111111;
assign micromatrizz[77][44] = 9'b111111111;
assign micromatrizz[77][45] = 9'b111111111;
assign micromatrizz[77][46] = 9'b111111111;
assign micromatrizz[77][47] = 9'b111111111;
assign micromatrizz[77][48] = 9'b111111111;
assign micromatrizz[77][49] = 9'b111111111;
assign micromatrizz[77][50] = 9'b111111111;
assign micromatrizz[77][51] = 9'b111111111;
assign micromatrizz[77][52] = 9'b111111111;
assign micromatrizz[77][53] = 9'b111111111;
assign micromatrizz[77][54] = 9'b111111111;
assign micromatrizz[77][55] = 9'b111111111;
assign micromatrizz[77][56] = 9'b111111111;
assign micromatrizz[77][57] = 9'b111111111;
assign micromatrizz[77][58] = 9'b111111111;
assign micromatrizz[77][59] = 9'b111111111;
assign micromatrizz[77][60] = 9'b111111111;
assign micromatrizz[77][61] = 9'b111111111;
assign micromatrizz[77][62] = 9'b111111111;
assign micromatrizz[77][63] = 9'b111111111;
assign micromatrizz[77][64] = 9'b111111111;
assign micromatrizz[77][65] = 9'b111111111;
assign micromatrizz[77][66] = 9'b111111111;
assign micromatrizz[77][67] = 9'b111111111;
assign micromatrizz[77][68] = 9'b111111111;
assign micromatrizz[77][69] = 9'b111111111;
assign micromatrizz[77][70] = 9'b111111111;
assign micromatrizz[77][71] = 9'b111111111;
assign micromatrizz[77][72] = 9'b111111111;
assign micromatrizz[77][73] = 9'b111111111;
assign micromatrizz[77][74] = 9'b111111111;
assign micromatrizz[77][75] = 9'b111111111;
assign micromatrizz[77][76] = 9'b111111111;
assign micromatrizz[77][77] = 9'b111111111;
assign micromatrizz[77][78] = 9'b111111111;
assign micromatrizz[77][79] = 9'b111111111;
assign micromatrizz[77][80] = 9'b111111111;
assign micromatrizz[77][81] = 9'b111111111;
assign micromatrizz[77][82] = 9'b111111111;
assign micromatrizz[77][83] = 9'b111111111;
assign micromatrizz[77][84] = 9'b111111111;
assign micromatrizz[77][85] = 9'b111111111;
assign micromatrizz[77][86] = 9'b111111111;
assign micromatrizz[77][87] = 9'b111111111;
assign micromatrizz[77][88] = 9'b111111111;
assign micromatrizz[77][89] = 9'b111111111;
assign micromatrizz[77][90] = 9'b111111111;
assign micromatrizz[77][91] = 9'b111111111;
assign micromatrizz[77][92] = 9'b111111111;
assign micromatrizz[77][93] = 9'b111111111;
assign micromatrizz[77][94] = 9'b111111111;
assign micromatrizz[77][95] = 9'b111111111;
assign micromatrizz[77][96] = 9'b111111111;
assign micromatrizz[77][97] = 9'b111111111;
assign micromatrizz[77][98] = 9'b111111111;
assign micromatrizz[77][99] = 9'b111111111;
assign micromatrizz[77][100] = 9'b111111111;
assign micromatrizz[77][101] = 9'b111111111;
assign micromatrizz[77][102] = 9'b111111111;
assign micromatrizz[77][103] = 9'b111111111;
assign micromatrizz[77][104] = 9'b111111111;
assign micromatrizz[77][105] = 9'b111111111;
assign micromatrizz[77][106] = 9'b111111111;
assign micromatrizz[77][107] = 9'b111111111;
assign micromatrizz[77][108] = 9'b111111111;
assign micromatrizz[77][109] = 9'b111111111;
assign micromatrizz[77][110] = 9'b111111111;
assign micromatrizz[77][111] = 9'b111111111;
assign micromatrizz[77][112] = 9'b111111111;
assign micromatrizz[77][113] = 9'b111111111;
assign micromatrizz[77][114] = 9'b111111111;
assign micromatrizz[77][115] = 9'b111111111;
assign micromatrizz[77][116] = 9'b111111111;
assign micromatrizz[77][117] = 9'b111111111;
assign micromatrizz[77][118] = 9'b111111111;
assign micromatrizz[77][119] = 9'b111111111;
assign micromatrizz[77][120] = 9'b111111111;
assign micromatrizz[77][121] = 9'b111111111;
assign micromatrizz[77][122] = 9'b111111111;
assign micromatrizz[77][123] = 9'b111111111;
assign micromatrizz[77][124] = 9'b111111111;
assign micromatrizz[77][125] = 9'b111111111;
assign micromatrizz[77][126] = 9'b111111111;
assign micromatrizz[77][127] = 9'b111111111;
assign micromatrizz[77][128] = 9'b111111111;
assign micromatrizz[77][129] = 9'b111111111;
assign micromatrizz[77][130] = 9'b111111111;
assign micromatrizz[77][131] = 9'b111111111;
assign micromatrizz[77][132] = 9'b111111111;
assign micromatrizz[77][133] = 9'b111111111;
assign micromatrizz[77][134] = 9'b111111111;
assign micromatrizz[77][135] = 9'b111111111;
assign micromatrizz[77][136] = 9'b111111111;
assign micromatrizz[77][137] = 9'b111111111;
assign micromatrizz[77][138] = 9'b111111111;
assign micromatrizz[77][139] = 9'b111111111;
assign micromatrizz[77][140] = 9'b111111111;
assign micromatrizz[77][141] = 9'b111111111;
assign micromatrizz[77][142] = 9'b111111111;
assign micromatrizz[77][143] = 9'b111111111;
assign micromatrizz[77][144] = 9'b111111111;
assign micromatrizz[77][145] = 9'b111111111;
assign micromatrizz[77][146] = 9'b111111111;
assign micromatrizz[77][147] = 9'b111111111;
assign micromatrizz[77][148] = 9'b111111111;
assign micromatrizz[77][149] = 9'b111111111;
assign micromatrizz[77][150] = 9'b111111111;
assign micromatrizz[77][151] = 9'b111111111;
assign micromatrizz[77][152] = 9'b111111111;
assign micromatrizz[77][153] = 9'b111111111;
assign micromatrizz[77][154] = 9'b111111111;
assign micromatrizz[77][155] = 9'b111111111;
assign micromatrizz[77][156] = 9'b111111111;
assign micromatrizz[77][157] = 9'b111111111;
assign micromatrizz[77][158] = 9'b111111111;
assign micromatrizz[77][159] = 9'b111111111;
assign micromatrizz[77][160] = 9'b111111111;
assign micromatrizz[77][161] = 9'b111111111;
assign micromatrizz[77][162] = 9'b111111111;
assign micromatrizz[77][163] = 9'b111111111;
assign micromatrizz[77][164] = 9'b111111111;
assign micromatrizz[77][165] = 9'b111111111;
assign micromatrizz[77][166] = 9'b111111111;
assign micromatrizz[77][167] = 9'b111111111;
assign micromatrizz[77][168] = 9'b111111111;
assign micromatrizz[77][169] = 9'b111111111;
assign micromatrizz[77][170] = 9'b111111111;
assign micromatrizz[77][171] = 9'b111111111;
assign micromatrizz[77][172] = 9'b111111111;
assign micromatrizz[77][173] = 9'b111111111;
assign micromatrizz[77][174] = 9'b111111111;
assign micromatrizz[77][175] = 9'b111111111;
assign micromatrizz[77][176] = 9'b111111111;
assign micromatrizz[77][177] = 9'b111111111;
assign micromatrizz[77][178] = 9'b111111111;
assign micromatrizz[77][179] = 9'b111111111;
assign micromatrizz[77][180] = 9'b111111111;
assign micromatrizz[77][181] = 9'b111111111;
assign micromatrizz[77][182] = 9'b111111111;
assign micromatrizz[77][183] = 9'b111111111;
assign micromatrizz[77][184] = 9'b111111111;
assign micromatrizz[77][185] = 9'b111111111;
assign micromatrizz[77][186] = 9'b111111111;
assign micromatrizz[77][187] = 9'b111111111;
assign micromatrizz[77][188] = 9'b111111111;
assign micromatrizz[77][189] = 9'b111111111;
assign micromatrizz[77][190] = 9'b111111111;
assign micromatrizz[77][191] = 9'b111111111;
assign micromatrizz[77][192] = 9'b111111111;
assign micromatrizz[77][193] = 9'b111111111;
assign micromatrizz[77][194] = 9'b111111111;
assign micromatrizz[77][195] = 9'b111111111;
assign micromatrizz[77][196] = 9'b111111111;
assign micromatrizz[77][197] = 9'b111111111;
assign micromatrizz[77][198] = 9'b111111111;
assign micromatrizz[77][199] = 9'b111111111;
assign micromatrizz[77][200] = 9'b111111111;
assign micromatrizz[77][201] = 9'b111111111;
assign micromatrizz[77][202] = 9'b111111111;
assign micromatrizz[77][203] = 9'b111111111;
assign micromatrizz[77][204] = 9'b111111111;
assign micromatrizz[77][205] = 9'b111111111;
assign micromatrizz[77][206] = 9'b111111111;
assign micromatrizz[77][207] = 9'b111111111;
assign micromatrizz[77][208] = 9'b111111111;
assign micromatrizz[77][209] = 9'b111111111;
assign micromatrizz[77][210] = 9'b111111111;
assign micromatrizz[77][211] = 9'b111111111;
assign micromatrizz[77][212] = 9'b111111111;
assign micromatrizz[77][213] = 9'b111111111;
assign micromatrizz[77][214] = 9'b111111111;
assign micromatrizz[77][215] = 9'b111111111;
assign micromatrizz[77][216] = 9'b111111111;
assign micromatrizz[77][217] = 9'b111111111;
assign micromatrizz[77][218] = 9'b111111111;
assign micromatrizz[77][219] = 9'b111111111;
assign micromatrizz[77][220] = 9'b111111111;
assign micromatrizz[77][221] = 9'b111111111;
assign micromatrizz[77][222] = 9'b111111111;
assign micromatrizz[77][223] = 9'b111111111;
assign micromatrizz[77][224] = 9'b111111111;
assign micromatrizz[77][225] = 9'b111111111;
assign micromatrizz[77][226] = 9'b111111111;
assign micromatrizz[77][227] = 9'b111111111;
assign micromatrizz[77][228] = 9'b111111111;
assign micromatrizz[77][229] = 9'b111111111;
assign micromatrizz[77][230] = 9'b111111111;
assign micromatrizz[77][231] = 9'b111111111;
assign micromatrizz[77][232] = 9'b111111111;
assign micromatrizz[77][233] = 9'b111111111;
assign micromatrizz[77][234] = 9'b111111111;
assign micromatrizz[77][235] = 9'b111111111;
assign micromatrizz[77][236] = 9'b111111111;
assign micromatrizz[77][237] = 9'b111111111;
assign micromatrizz[77][238] = 9'b111111111;
assign micromatrizz[77][239] = 9'b111111111;
assign micromatrizz[77][240] = 9'b111111111;
assign micromatrizz[77][241] = 9'b111111111;
assign micromatrizz[77][242] = 9'b111111111;
assign micromatrizz[77][243] = 9'b111111111;
assign micromatrizz[77][244] = 9'b111111111;
assign micromatrizz[77][245] = 9'b111111111;
assign micromatrizz[77][246] = 9'b111111111;
assign micromatrizz[77][247] = 9'b111111111;
assign micromatrizz[77][248] = 9'b111111111;
assign micromatrizz[77][249] = 9'b111111111;
assign micromatrizz[77][250] = 9'b111111111;
assign micromatrizz[77][251] = 9'b111111111;
assign micromatrizz[77][252] = 9'b111111111;
assign micromatrizz[77][253] = 9'b111111111;
assign micromatrizz[77][254] = 9'b111111111;
assign micromatrizz[77][255] = 9'b111111111;
assign micromatrizz[77][256] = 9'b111111111;
assign micromatrizz[77][257] = 9'b111111111;
assign micromatrizz[77][258] = 9'b111111111;
assign micromatrizz[77][259] = 9'b111111111;
assign micromatrizz[77][260] = 9'b111111111;
assign micromatrizz[77][261] = 9'b111111111;
assign micromatrizz[77][262] = 9'b111111111;
assign micromatrizz[77][263] = 9'b111111111;
assign micromatrizz[77][264] = 9'b111111111;
assign micromatrizz[77][265] = 9'b111111111;
assign micromatrizz[77][266] = 9'b111111111;
assign micromatrizz[77][267] = 9'b111111111;
assign micromatrizz[77][268] = 9'b111111111;
assign micromatrizz[77][269] = 9'b111111111;
assign micromatrizz[77][270] = 9'b111111111;
assign micromatrizz[77][271] = 9'b111111111;
assign micromatrizz[77][272] = 9'b111111111;
assign micromatrizz[77][273] = 9'b111111111;
assign micromatrizz[77][274] = 9'b111111111;
assign micromatrizz[77][275] = 9'b111111111;
assign micromatrizz[77][276] = 9'b111111111;
assign micromatrizz[77][277] = 9'b111111111;
assign micromatrizz[77][278] = 9'b111111111;
assign micromatrizz[77][279] = 9'b111111111;
assign micromatrizz[77][280] = 9'b111111111;
assign micromatrizz[77][281] = 9'b111111111;
assign micromatrizz[77][282] = 9'b111111111;
assign micromatrizz[77][283] = 9'b111111111;
assign micromatrizz[77][284] = 9'b111111111;
assign micromatrizz[77][285] = 9'b111111111;
assign micromatrizz[77][286] = 9'b111111111;
assign micromatrizz[77][287] = 9'b111111111;
assign micromatrizz[77][288] = 9'b111111111;
assign micromatrizz[77][289] = 9'b111111111;
assign micromatrizz[77][290] = 9'b111111111;
assign micromatrizz[77][291] = 9'b111111111;
assign micromatrizz[77][292] = 9'b111111111;
assign micromatrizz[77][293] = 9'b111111111;
assign micromatrizz[77][294] = 9'b111111111;
assign micromatrizz[77][295] = 9'b111111111;
assign micromatrizz[77][296] = 9'b111111111;
assign micromatrizz[77][297] = 9'b111111111;
assign micromatrizz[77][298] = 9'b111111111;
assign micromatrizz[77][299] = 9'b111111111;
assign micromatrizz[77][300] = 9'b111111111;
assign micromatrizz[77][301] = 9'b111111111;
assign micromatrizz[77][302] = 9'b111111111;
assign micromatrizz[77][303] = 9'b111111111;
assign micromatrizz[77][304] = 9'b111111111;
assign micromatrizz[77][305] = 9'b111111111;
assign micromatrizz[77][306] = 9'b111111111;
assign micromatrizz[77][307] = 9'b111111111;
assign micromatrizz[77][308] = 9'b111111111;
assign micromatrizz[77][309] = 9'b111111111;
assign micromatrizz[77][310] = 9'b111111111;
assign micromatrizz[77][311] = 9'b111111111;
assign micromatrizz[77][312] = 9'b111111111;
assign micromatrizz[77][313] = 9'b111111111;
assign micromatrizz[77][314] = 9'b111111111;
assign micromatrizz[77][315] = 9'b111111111;
assign micromatrizz[77][316] = 9'b111111111;
assign micromatrizz[77][317] = 9'b111111111;
assign micromatrizz[77][318] = 9'b111111111;
assign micromatrizz[77][319] = 9'b111111111;
assign micromatrizz[77][320] = 9'b111111111;
assign micromatrizz[77][321] = 9'b111111111;
assign micromatrizz[77][322] = 9'b111111111;
assign micromatrizz[77][323] = 9'b111111111;
assign micromatrizz[77][324] = 9'b111111111;
assign micromatrizz[77][325] = 9'b111111111;
assign micromatrizz[77][326] = 9'b111111111;
assign micromatrizz[77][327] = 9'b111111111;
assign micromatrizz[77][328] = 9'b111111111;
assign micromatrizz[77][329] = 9'b111111111;
assign micromatrizz[77][330] = 9'b111111111;
assign micromatrizz[77][331] = 9'b111111111;
assign micromatrizz[77][332] = 9'b111111111;
assign micromatrizz[77][333] = 9'b111111111;
assign micromatrizz[77][334] = 9'b111111111;
assign micromatrizz[77][335] = 9'b111111111;
assign micromatrizz[77][336] = 9'b111111111;
assign micromatrizz[77][337] = 9'b111111111;
assign micromatrizz[77][338] = 9'b111111111;
assign micromatrizz[77][339] = 9'b111111111;
assign micromatrizz[77][340] = 9'b111111111;
assign micromatrizz[77][341] = 9'b111111111;
assign micromatrizz[77][342] = 9'b111111111;
assign micromatrizz[77][343] = 9'b111111111;
assign micromatrizz[77][344] = 9'b111111111;
assign micromatrizz[77][345] = 9'b111111111;
assign micromatrizz[77][346] = 9'b111111111;
assign micromatrizz[77][347] = 9'b111111111;
assign micromatrizz[77][348] = 9'b111111111;
assign micromatrizz[77][349] = 9'b111111111;
assign micromatrizz[77][350] = 9'b111111111;
assign micromatrizz[77][351] = 9'b111111111;
assign micromatrizz[77][352] = 9'b111111111;
assign micromatrizz[77][353] = 9'b111111111;
assign micromatrizz[77][354] = 9'b111111111;
assign micromatrizz[77][355] = 9'b111111111;
assign micromatrizz[77][356] = 9'b111111111;
assign micromatrizz[77][357] = 9'b111111111;
assign micromatrizz[77][358] = 9'b111111111;
assign micromatrizz[77][359] = 9'b111111111;
assign micromatrizz[77][360] = 9'b111111111;
assign micromatrizz[77][361] = 9'b111111111;
assign micromatrizz[77][362] = 9'b111111111;
assign micromatrizz[77][363] = 9'b111111111;
assign micromatrizz[77][364] = 9'b111111111;
assign micromatrizz[77][365] = 9'b111111111;
assign micromatrizz[77][366] = 9'b111111111;
assign micromatrizz[77][367] = 9'b111111111;
assign micromatrizz[77][368] = 9'b111111111;
assign micromatrizz[77][369] = 9'b111111111;
assign micromatrizz[77][370] = 9'b111111111;
assign micromatrizz[77][371] = 9'b111111111;
assign micromatrizz[77][372] = 9'b111111111;
assign micromatrizz[77][373] = 9'b111111111;
assign micromatrizz[77][374] = 9'b111111111;
assign micromatrizz[77][375] = 9'b111111111;
assign micromatrizz[77][376] = 9'b111111111;
assign micromatrizz[77][377] = 9'b111111111;
assign micromatrizz[77][378] = 9'b111111111;
assign micromatrizz[77][379] = 9'b111111111;
assign micromatrizz[77][380] = 9'b111111111;
assign micromatrizz[77][381] = 9'b111111111;
assign micromatrizz[77][382] = 9'b111111111;
assign micromatrizz[77][383] = 9'b111111111;
assign micromatrizz[77][384] = 9'b111111111;
assign micromatrizz[77][385] = 9'b111111111;
assign micromatrizz[77][386] = 9'b111111111;
assign micromatrizz[77][387] = 9'b111111111;
assign micromatrizz[77][388] = 9'b111111111;
assign micromatrizz[77][389] = 9'b111111111;
assign micromatrizz[77][390] = 9'b111111111;
assign micromatrizz[77][391] = 9'b111111111;
assign micromatrizz[77][392] = 9'b111111111;
assign micromatrizz[77][393] = 9'b111111111;
assign micromatrizz[77][394] = 9'b111111111;
assign micromatrizz[77][395] = 9'b111111111;
assign micromatrizz[77][396] = 9'b111111111;
assign micromatrizz[77][397] = 9'b111111111;
assign micromatrizz[77][398] = 9'b111111111;
assign micromatrizz[77][399] = 9'b111111111;
assign micromatrizz[77][400] = 9'b111111111;
assign micromatrizz[77][401] = 9'b111111111;
assign micromatrizz[77][402] = 9'b111111111;
assign micromatrizz[77][403] = 9'b111111111;
assign micromatrizz[77][404] = 9'b111111111;
assign micromatrizz[77][405] = 9'b111111111;
assign micromatrizz[77][406] = 9'b111111111;
assign micromatrizz[77][407] = 9'b111111111;
assign micromatrizz[77][408] = 9'b111111111;
assign micromatrizz[77][409] = 9'b111111111;
assign micromatrizz[77][410] = 9'b111111111;
assign micromatrizz[77][411] = 9'b111111111;
assign micromatrizz[77][412] = 9'b111111111;
assign micromatrizz[77][413] = 9'b111111111;
assign micromatrizz[77][414] = 9'b111111111;
assign micromatrizz[77][415] = 9'b111111111;
assign micromatrizz[77][416] = 9'b111111111;
assign micromatrizz[77][417] = 9'b111111111;
assign micromatrizz[77][418] = 9'b111111111;
assign micromatrizz[77][419] = 9'b111111111;
assign micromatrizz[77][420] = 9'b111111111;
assign micromatrizz[77][421] = 9'b111111111;
assign micromatrizz[77][422] = 9'b111111111;
assign micromatrizz[77][423] = 9'b111111111;
assign micromatrizz[77][424] = 9'b111111111;
assign micromatrizz[77][425] = 9'b111111111;
assign micromatrizz[77][426] = 9'b111111111;
assign micromatrizz[77][427] = 9'b111111111;
assign micromatrizz[77][428] = 9'b111111111;
assign micromatrizz[77][429] = 9'b111111111;
assign micromatrizz[77][430] = 9'b111111111;
assign micromatrizz[77][431] = 9'b111111111;
assign micromatrizz[77][432] = 9'b111111111;
assign micromatrizz[77][433] = 9'b111111111;
assign micromatrizz[77][434] = 9'b111111111;
assign micromatrizz[77][435] = 9'b111111111;
assign micromatrizz[77][436] = 9'b111111111;
assign micromatrizz[77][437] = 9'b111111111;
assign micromatrizz[77][438] = 9'b111111111;
assign micromatrizz[77][439] = 9'b111111111;
assign micromatrizz[77][440] = 9'b111111111;
assign micromatrizz[77][441] = 9'b111111111;
assign micromatrizz[77][442] = 9'b111111111;
assign micromatrizz[77][443] = 9'b111111111;
assign micromatrizz[77][444] = 9'b111111111;
assign micromatrizz[77][445] = 9'b111111111;
assign micromatrizz[77][446] = 9'b111111111;
assign micromatrizz[77][447] = 9'b111111111;
assign micromatrizz[77][448] = 9'b111111111;
assign micromatrizz[77][449] = 9'b111111111;
assign micromatrizz[77][450] = 9'b111111111;
assign micromatrizz[77][451] = 9'b111111111;
assign micromatrizz[77][452] = 9'b111111111;
assign micromatrizz[77][453] = 9'b111111111;
assign micromatrizz[77][454] = 9'b111111111;
assign micromatrizz[77][455] = 9'b111111111;
assign micromatrizz[77][456] = 9'b111111111;
assign micromatrizz[77][457] = 9'b111111111;
assign micromatrizz[77][458] = 9'b111111111;
assign micromatrizz[77][459] = 9'b111111111;
assign micromatrizz[77][460] = 9'b111111111;
assign micromatrizz[77][461] = 9'b111111111;
assign micromatrizz[77][462] = 9'b111111111;
assign micromatrizz[77][463] = 9'b111111111;
assign micromatrizz[77][464] = 9'b111111111;
assign micromatrizz[77][465] = 9'b111111111;
assign micromatrizz[77][466] = 9'b111111111;
assign micromatrizz[77][467] = 9'b111111111;
assign micromatrizz[77][468] = 9'b111111111;
assign micromatrizz[77][469] = 9'b111111111;
assign micromatrizz[77][470] = 9'b111111111;
assign micromatrizz[77][471] = 9'b111111111;
assign micromatrizz[77][472] = 9'b111111111;
assign micromatrizz[77][473] = 9'b111111111;
assign micromatrizz[77][474] = 9'b111111111;
assign micromatrizz[77][475] = 9'b111111111;
assign micromatrizz[77][476] = 9'b111111111;
assign micromatrizz[77][477] = 9'b111111111;
assign micromatrizz[77][478] = 9'b111111111;
assign micromatrizz[77][479] = 9'b111111111;
assign micromatrizz[77][480] = 9'b111111111;
assign micromatrizz[77][481] = 9'b111111111;
assign micromatrizz[77][482] = 9'b111111111;
assign micromatrizz[77][483] = 9'b111111111;
assign micromatrizz[77][484] = 9'b111111111;
assign micromatrizz[77][485] = 9'b111111111;
assign micromatrizz[77][486] = 9'b111111111;
assign micromatrizz[77][487] = 9'b111111111;
assign micromatrizz[77][488] = 9'b111111111;
assign micromatrizz[77][489] = 9'b111111111;
assign micromatrizz[77][490] = 9'b111111111;
assign micromatrizz[77][491] = 9'b111111111;
assign micromatrizz[77][492] = 9'b111111111;
assign micromatrizz[77][493] = 9'b111111111;
assign micromatrizz[77][494] = 9'b111111111;
assign micromatrizz[77][495] = 9'b111111111;
assign micromatrizz[77][496] = 9'b111111111;
assign micromatrizz[77][497] = 9'b111111111;
assign micromatrizz[77][498] = 9'b111111111;
assign micromatrizz[77][499] = 9'b111111111;
assign micromatrizz[77][500] = 9'b111111111;
assign micromatrizz[77][501] = 9'b111111111;
assign micromatrizz[77][502] = 9'b111111111;
assign micromatrizz[77][503] = 9'b111111111;
assign micromatrizz[77][504] = 9'b111111111;
assign micromatrizz[77][505] = 9'b111111111;
assign micromatrizz[77][506] = 9'b111111111;
assign micromatrizz[77][507] = 9'b111111111;
assign micromatrizz[77][508] = 9'b111111111;
assign micromatrizz[77][509] = 9'b111111111;
assign micromatrizz[77][510] = 9'b111111111;
assign micromatrizz[77][511] = 9'b111111111;
assign micromatrizz[77][512] = 9'b111111111;
assign micromatrizz[77][513] = 9'b111111111;
assign micromatrizz[77][514] = 9'b111111111;
assign micromatrizz[77][515] = 9'b111111111;
assign micromatrizz[77][516] = 9'b111111111;
assign micromatrizz[77][517] = 9'b111111111;
assign micromatrizz[77][518] = 9'b111111111;
assign micromatrizz[77][519] = 9'b111111111;
assign micromatrizz[77][520] = 9'b111111111;
assign micromatrizz[77][521] = 9'b111111111;
assign micromatrizz[77][522] = 9'b111111111;
assign micromatrizz[77][523] = 9'b111111111;
assign micromatrizz[77][524] = 9'b111111111;
assign micromatrizz[77][525] = 9'b111111111;
assign micromatrizz[77][526] = 9'b111111111;
assign micromatrizz[77][527] = 9'b111111111;
assign micromatrizz[77][528] = 9'b111111111;
assign micromatrizz[77][529] = 9'b111111111;
assign micromatrizz[77][530] = 9'b111111111;
assign micromatrizz[77][531] = 9'b111111111;
assign micromatrizz[77][532] = 9'b111111111;
assign micromatrizz[77][533] = 9'b111111111;
assign micromatrizz[77][534] = 9'b111111111;
assign micromatrizz[77][535] = 9'b111111111;
assign micromatrizz[77][536] = 9'b111111111;
assign micromatrizz[77][537] = 9'b111111111;
assign micromatrizz[77][538] = 9'b111111111;
assign micromatrizz[77][539] = 9'b111111111;
assign micromatrizz[77][540] = 9'b111111111;
assign micromatrizz[77][541] = 9'b111111111;
assign micromatrizz[77][542] = 9'b111111111;
assign micromatrizz[77][543] = 9'b111111111;
assign micromatrizz[77][544] = 9'b111111111;
assign micromatrizz[77][545] = 9'b111111111;
assign micromatrizz[77][546] = 9'b111111111;
assign micromatrizz[77][547] = 9'b111111111;
assign micromatrizz[77][548] = 9'b111111111;
assign micromatrizz[77][549] = 9'b111111111;
assign micromatrizz[77][550] = 9'b111111111;
assign micromatrizz[77][551] = 9'b111111111;
assign micromatrizz[77][552] = 9'b111111111;
assign micromatrizz[77][553] = 9'b111111111;
assign micromatrizz[77][554] = 9'b111111111;
assign micromatrizz[77][555] = 9'b111111111;
assign micromatrizz[77][556] = 9'b111111111;
assign micromatrizz[77][557] = 9'b111111111;
assign micromatrizz[77][558] = 9'b111111111;
assign micromatrizz[77][559] = 9'b111111111;
assign micromatrizz[77][560] = 9'b111111111;
assign micromatrizz[77][561] = 9'b111111111;
assign micromatrizz[77][562] = 9'b111111111;
assign micromatrizz[77][563] = 9'b111111111;
assign micromatrizz[77][564] = 9'b111111111;
assign micromatrizz[77][565] = 9'b111111111;
assign micromatrizz[77][566] = 9'b111111111;
assign micromatrizz[77][567] = 9'b111111111;
assign micromatrizz[77][568] = 9'b111111111;
assign micromatrizz[77][569] = 9'b111111111;
assign micromatrizz[77][570] = 9'b111111111;
assign micromatrizz[77][571] = 9'b111111111;
assign micromatrizz[77][572] = 9'b111111111;
assign micromatrizz[77][573] = 9'b111111111;
assign micromatrizz[77][574] = 9'b111111111;
assign micromatrizz[77][575] = 9'b111111111;
assign micromatrizz[77][576] = 9'b111111111;
assign micromatrizz[77][577] = 9'b111111111;
assign micromatrizz[77][578] = 9'b111111111;
assign micromatrizz[77][579] = 9'b111111111;
assign micromatrizz[77][580] = 9'b111111111;
assign micromatrizz[77][581] = 9'b111111111;
assign micromatrizz[77][582] = 9'b111111111;
assign micromatrizz[77][583] = 9'b111111111;
assign micromatrizz[77][584] = 9'b111111111;
assign micromatrizz[77][585] = 9'b111111111;
assign micromatrizz[77][586] = 9'b111111111;
assign micromatrizz[77][587] = 9'b111111111;
assign micromatrizz[77][588] = 9'b111111111;
assign micromatrizz[77][589] = 9'b111111111;
assign micromatrizz[77][590] = 9'b111111111;
assign micromatrizz[77][591] = 9'b111111111;
assign micromatrizz[77][592] = 9'b111111111;
assign micromatrizz[77][593] = 9'b111111111;
assign micromatrizz[77][594] = 9'b111111111;
assign micromatrizz[77][595] = 9'b111111111;
assign micromatrizz[77][596] = 9'b111111111;
assign micromatrizz[77][597] = 9'b111111111;
assign micromatrizz[77][598] = 9'b111111111;
assign micromatrizz[77][599] = 9'b111111111;
assign micromatrizz[77][600] = 9'b111111111;
assign micromatrizz[77][601] = 9'b111111111;
assign micromatrizz[77][602] = 9'b111111111;
assign micromatrizz[77][603] = 9'b111111111;
assign micromatrizz[77][604] = 9'b111111111;
assign micromatrizz[77][605] = 9'b111111111;
assign micromatrizz[77][606] = 9'b111111111;
assign micromatrizz[77][607] = 9'b111111111;
assign micromatrizz[77][608] = 9'b111111111;
assign micromatrizz[77][609] = 9'b111111111;
assign micromatrizz[77][610] = 9'b111111111;
assign micromatrizz[77][611] = 9'b111111111;
assign micromatrizz[77][612] = 9'b111111111;
assign micromatrizz[77][613] = 9'b111111111;
assign micromatrizz[77][614] = 9'b111111111;
assign micromatrizz[77][615] = 9'b111111111;
assign micromatrizz[77][616] = 9'b111111111;
assign micromatrizz[77][617] = 9'b111111111;
assign micromatrizz[77][618] = 9'b111111111;
assign micromatrizz[77][619] = 9'b111111111;
assign micromatrizz[77][620] = 9'b111111111;
assign micromatrizz[77][621] = 9'b111111111;
assign micromatrizz[77][622] = 9'b111111111;
assign micromatrizz[77][623] = 9'b111111111;
assign micromatrizz[77][624] = 9'b111111111;
assign micromatrizz[77][625] = 9'b111111111;
assign micromatrizz[77][626] = 9'b111111111;
assign micromatrizz[77][627] = 9'b111111111;
assign micromatrizz[77][628] = 9'b111111111;
assign micromatrizz[77][629] = 9'b111111111;
assign micromatrizz[77][630] = 9'b111111111;
assign micromatrizz[77][631] = 9'b111111111;
assign micromatrizz[77][632] = 9'b111111111;
assign micromatrizz[77][633] = 9'b111111111;
assign micromatrizz[77][634] = 9'b111111111;
assign micromatrizz[77][635] = 9'b111111111;
assign micromatrizz[77][636] = 9'b111111111;
assign micromatrizz[77][637] = 9'b111111111;
assign micromatrizz[77][638] = 9'b111111111;
assign micromatrizz[77][639] = 9'b111111111;
assign micromatrizz[78][0] = 9'b111111111;
assign micromatrizz[78][1] = 9'b111111111;
assign micromatrizz[78][2] = 9'b111111111;
assign micromatrizz[78][3] = 9'b111111111;
assign micromatrizz[78][4] = 9'b111111111;
assign micromatrizz[78][5] = 9'b111111111;
assign micromatrizz[78][6] = 9'b111111111;
assign micromatrizz[78][7] = 9'b111111111;
assign micromatrizz[78][8] = 9'b111111111;
assign micromatrizz[78][9] = 9'b111111111;
assign micromatrizz[78][10] = 9'b111111111;
assign micromatrizz[78][11] = 9'b111111111;
assign micromatrizz[78][12] = 9'b111111111;
assign micromatrizz[78][13] = 9'b111111111;
assign micromatrizz[78][14] = 9'b111111111;
assign micromatrizz[78][15] = 9'b111111111;
assign micromatrizz[78][16] = 9'b111111111;
assign micromatrizz[78][17] = 9'b111111111;
assign micromatrizz[78][18] = 9'b111111111;
assign micromatrizz[78][19] = 9'b111111111;
assign micromatrizz[78][20] = 9'b111111111;
assign micromatrizz[78][21] = 9'b111111111;
assign micromatrizz[78][22] = 9'b111111111;
assign micromatrizz[78][23] = 9'b111111111;
assign micromatrizz[78][24] = 9'b111111111;
assign micromatrizz[78][25] = 9'b111111111;
assign micromatrizz[78][26] = 9'b111111111;
assign micromatrizz[78][27] = 9'b111111111;
assign micromatrizz[78][28] = 9'b111111111;
assign micromatrizz[78][29] = 9'b111111111;
assign micromatrizz[78][30] = 9'b111111111;
assign micromatrizz[78][31] = 9'b111111111;
assign micromatrizz[78][32] = 9'b111111111;
assign micromatrizz[78][33] = 9'b111111111;
assign micromatrizz[78][34] = 9'b111111111;
assign micromatrizz[78][35] = 9'b111111111;
assign micromatrizz[78][36] = 9'b111111111;
assign micromatrizz[78][37] = 9'b111111111;
assign micromatrizz[78][38] = 9'b111111111;
assign micromatrizz[78][39] = 9'b111111111;
assign micromatrizz[78][40] = 9'b111111111;
assign micromatrizz[78][41] = 9'b111111111;
assign micromatrizz[78][42] = 9'b111111111;
assign micromatrizz[78][43] = 9'b111111111;
assign micromatrizz[78][44] = 9'b111111111;
assign micromatrizz[78][45] = 9'b111111111;
assign micromatrizz[78][46] = 9'b111111111;
assign micromatrizz[78][47] = 9'b111111111;
assign micromatrizz[78][48] = 9'b111111111;
assign micromatrizz[78][49] = 9'b111111111;
assign micromatrizz[78][50] = 9'b111111111;
assign micromatrizz[78][51] = 9'b111111111;
assign micromatrizz[78][52] = 9'b111111111;
assign micromatrizz[78][53] = 9'b111111111;
assign micromatrizz[78][54] = 9'b111111111;
assign micromatrizz[78][55] = 9'b111111111;
assign micromatrizz[78][56] = 9'b111111111;
assign micromatrizz[78][57] = 9'b111111111;
assign micromatrizz[78][58] = 9'b111111111;
assign micromatrizz[78][59] = 9'b111111111;
assign micromatrizz[78][60] = 9'b111111111;
assign micromatrizz[78][61] = 9'b111111111;
assign micromatrizz[78][62] = 9'b111111111;
assign micromatrizz[78][63] = 9'b111111111;
assign micromatrizz[78][64] = 9'b111111111;
assign micromatrizz[78][65] = 9'b111111111;
assign micromatrizz[78][66] = 9'b111111111;
assign micromatrizz[78][67] = 9'b111111111;
assign micromatrizz[78][68] = 9'b111111111;
assign micromatrizz[78][69] = 9'b111111111;
assign micromatrizz[78][70] = 9'b111111111;
assign micromatrizz[78][71] = 9'b111111111;
assign micromatrizz[78][72] = 9'b111111111;
assign micromatrizz[78][73] = 9'b111111111;
assign micromatrizz[78][74] = 9'b111111111;
assign micromatrizz[78][75] = 9'b111111111;
assign micromatrizz[78][76] = 9'b111111111;
assign micromatrizz[78][77] = 9'b111111111;
assign micromatrizz[78][78] = 9'b111111111;
assign micromatrizz[78][79] = 9'b111111111;
assign micromatrizz[78][80] = 9'b111111111;
assign micromatrizz[78][81] = 9'b111111111;
assign micromatrizz[78][82] = 9'b111111111;
assign micromatrizz[78][83] = 9'b111111111;
assign micromatrizz[78][84] = 9'b111111111;
assign micromatrizz[78][85] = 9'b111111111;
assign micromatrizz[78][86] = 9'b111111111;
assign micromatrizz[78][87] = 9'b111111111;
assign micromatrizz[78][88] = 9'b111111111;
assign micromatrizz[78][89] = 9'b111111111;
assign micromatrizz[78][90] = 9'b111111111;
assign micromatrizz[78][91] = 9'b111111111;
assign micromatrizz[78][92] = 9'b111111111;
assign micromatrizz[78][93] = 9'b111111111;
assign micromatrizz[78][94] = 9'b111111111;
assign micromatrizz[78][95] = 9'b111111111;
assign micromatrizz[78][96] = 9'b111111111;
assign micromatrizz[78][97] = 9'b111111111;
assign micromatrizz[78][98] = 9'b111111111;
assign micromatrizz[78][99] = 9'b111111111;
assign micromatrizz[78][100] = 9'b111111111;
assign micromatrizz[78][101] = 9'b111111111;
assign micromatrizz[78][102] = 9'b111111111;
assign micromatrizz[78][103] = 9'b111111111;
assign micromatrizz[78][104] = 9'b111111111;
assign micromatrizz[78][105] = 9'b111111111;
assign micromatrizz[78][106] = 9'b111111111;
assign micromatrizz[78][107] = 9'b111111111;
assign micromatrizz[78][108] = 9'b111111111;
assign micromatrizz[78][109] = 9'b111111111;
assign micromatrizz[78][110] = 9'b111111111;
assign micromatrizz[78][111] = 9'b111111111;
assign micromatrizz[78][112] = 9'b111111111;
assign micromatrizz[78][113] = 9'b111111111;
assign micromatrizz[78][114] = 9'b111111111;
assign micromatrizz[78][115] = 9'b111111111;
assign micromatrizz[78][116] = 9'b111111111;
assign micromatrizz[78][117] = 9'b111111111;
assign micromatrizz[78][118] = 9'b111111111;
assign micromatrizz[78][119] = 9'b111111111;
assign micromatrizz[78][120] = 9'b111111111;
assign micromatrizz[78][121] = 9'b111111111;
assign micromatrizz[78][122] = 9'b111111111;
assign micromatrizz[78][123] = 9'b111111111;
assign micromatrizz[78][124] = 9'b111111111;
assign micromatrizz[78][125] = 9'b111111111;
assign micromatrizz[78][126] = 9'b111111111;
assign micromatrizz[78][127] = 9'b111111111;
assign micromatrizz[78][128] = 9'b111111111;
assign micromatrizz[78][129] = 9'b111111111;
assign micromatrizz[78][130] = 9'b111111111;
assign micromatrizz[78][131] = 9'b111111111;
assign micromatrizz[78][132] = 9'b111111111;
assign micromatrizz[78][133] = 9'b111111111;
assign micromatrizz[78][134] = 9'b111111111;
assign micromatrizz[78][135] = 9'b111111111;
assign micromatrizz[78][136] = 9'b111111111;
assign micromatrizz[78][137] = 9'b111111111;
assign micromatrizz[78][138] = 9'b111111111;
assign micromatrizz[78][139] = 9'b111111111;
assign micromatrizz[78][140] = 9'b111111111;
assign micromatrizz[78][141] = 9'b111111111;
assign micromatrizz[78][142] = 9'b111111111;
assign micromatrizz[78][143] = 9'b111111111;
assign micromatrizz[78][144] = 9'b111111111;
assign micromatrizz[78][145] = 9'b111111111;
assign micromatrizz[78][146] = 9'b111111111;
assign micromatrizz[78][147] = 9'b111111111;
assign micromatrizz[78][148] = 9'b111111111;
assign micromatrizz[78][149] = 9'b111111111;
assign micromatrizz[78][150] = 9'b111111111;
assign micromatrizz[78][151] = 9'b111111111;
assign micromatrizz[78][152] = 9'b111111111;
assign micromatrizz[78][153] = 9'b111111111;
assign micromatrizz[78][154] = 9'b111111111;
assign micromatrizz[78][155] = 9'b111111111;
assign micromatrizz[78][156] = 9'b111111111;
assign micromatrizz[78][157] = 9'b111111111;
assign micromatrizz[78][158] = 9'b111111111;
assign micromatrizz[78][159] = 9'b111111111;
assign micromatrizz[78][160] = 9'b111111111;
assign micromatrizz[78][161] = 9'b111111111;
assign micromatrizz[78][162] = 9'b111111111;
assign micromatrizz[78][163] = 9'b111111111;
assign micromatrizz[78][164] = 9'b111111111;
assign micromatrizz[78][165] = 9'b111111111;
assign micromatrizz[78][166] = 9'b111111111;
assign micromatrizz[78][167] = 9'b111111111;
assign micromatrizz[78][168] = 9'b111111111;
assign micromatrizz[78][169] = 9'b111111111;
assign micromatrizz[78][170] = 9'b111111111;
assign micromatrizz[78][171] = 9'b111111111;
assign micromatrizz[78][172] = 9'b111111111;
assign micromatrizz[78][173] = 9'b111111111;
assign micromatrizz[78][174] = 9'b111111111;
assign micromatrizz[78][175] = 9'b111111111;
assign micromatrizz[78][176] = 9'b111111111;
assign micromatrizz[78][177] = 9'b111111111;
assign micromatrizz[78][178] = 9'b111111111;
assign micromatrizz[78][179] = 9'b111111111;
assign micromatrizz[78][180] = 9'b111111111;
assign micromatrizz[78][181] = 9'b111111111;
assign micromatrizz[78][182] = 9'b111111111;
assign micromatrizz[78][183] = 9'b111111111;
assign micromatrizz[78][184] = 9'b111111111;
assign micromatrizz[78][185] = 9'b111111111;
assign micromatrizz[78][186] = 9'b111111111;
assign micromatrizz[78][187] = 9'b111111111;
assign micromatrizz[78][188] = 9'b111111111;
assign micromatrizz[78][189] = 9'b111111111;
assign micromatrizz[78][190] = 9'b111111111;
assign micromatrizz[78][191] = 9'b111111111;
assign micromatrizz[78][192] = 9'b111111111;
assign micromatrizz[78][193] = 9'b111111111;
assign micromatrizz[78][194] = 9'b111111111;
assign micromatrizz[78][195] = 9'b111111111;
assign micromatrizz[78][196] = 9'b111111111;
assign micromatrizz[78][197] = 9'b111111111;
assign micromatrizz[78][198] = 9'b111111111;
assign micromatrizz[78][199] = 9'b111111111;
assign micromatrizz[78][200] = 9'b111111111;
assign micromatrizz[78][201] = 9'b111111111;
assign micromatrizz[78][202] = 9'b111111111;
assign micromatrizz[78][203] = 9'b111111111;
assign micromatrizz[78][204] = 9'b111111111;
assign micromatrizz[78][205] = 9'b111111111;
assign micromatrizz[78][206] = 9'b111111111;
assign micromatrizz[78][207] = 9'b111111111;
assign micromatrizz[78][208] = 9'b111111111;
assign micromatrizz[78][209] = 9'b111111111;
assign micromatrizz[78][210] = 9'b111111111;
assign micromatrizz[78][211] = 9'b111111111;
assign micromatrizz[78][212] = 9'b111111111;
assign micromatrizz[78][213] = 9'b111111111;
assign micromatrizz[78][214] = 9'b111111111;
assign micromatrizz[78][215] = 9'b111111111;
assign micromatrizz[78][216] = 9'b111111111;
assign micromatrizz[78][217] = 9'b111111111;
assign micromatrizz[78][218] = 9'b111111111;
assign micromatrizz[78][219] = 9'b111111111;
assign micromatrizz[78][220] = 9'b111111111;
assign micromatrizz[78][221] = 9'b111111111;
assign micromatrizz[78][222] = 9'b111111111;
assign micromatrizz[78][223] = 9'b111111111;
assign micromatrizz[78][224] = 9'b111111111;
assign micromatrizz[78][225] = 9'b111111111;
assign micromatrizz[78][226] = 9'b111111111;
assign micromatrizz[78][227] = 9'b111111111;
assign micromatrizz[78][228] = 9'b111111111;
assign micromatrizz[78][229] = 9'b111111111;
assign micromatrizz[78][230] = 9'b111111111;
assign micromatrizz[78][231] = 9'b111111111;
assign micromatrizz[78][232] = 9'b111111111;
assign micromatrizz[78][233] = 9'b111111111;
assign micromatrizz[78][234] = 9'b111111111;
assign micromatrizz[78][235] = 9'b111111111;
assign micromatrizz[78][236] = 9'b111111111;
assign micromatrizz[78][237] = 9'b111111111;
assign micromatrizz[78][238] = 9'b111111111;
assign micromatrizz[78][239] = 9'b111111111;
assign micromatrizz[78][240] = 9'b111111111;
assign micromatrizz[78][241] = 9'b111111111;
assign micromatrizz[78][242] = 9'b111111111;
assign micromatrizz[78][243] = 9'b111111111;
assign micromatrizz[78][244] = 9'b111111111;
assign micromatrizz[78][245] = 9'b111111111;
assign micromatrizz[78][246] = 9'b111111111;
assign micromatrizz[78][247] = 9'b111111111;
assign micromatrizz[78][248] = 9'b111111111;
assign micromatrizz[78][249] = 9'b111111111;
assign micromatrizz[78][250] = 9'b111111111;
assign micromatrizz[78][251] = 9'b111111111;
assign micromatrizz[78][252] = 9'b111111111;
assign micromatrizz[78][253] = 9'b111111111;
assign micromatrizz[78][254] = 9'b111111111;
assign micromatrizz[78][255] = 9'b111111111;
assign micromatrizz[78][256] = 9'b111111111;
assign micromatrizz[78][257] = 9'b111111111;
assign micromatrizz[78][258] = 9'b111111111;
assign micromatrizz[78][259] = 9'b111111111;
assign micromatrizz[78][260] = 9'b111111111;
assign micromatrizz[78][261] = 9'b111111111;
assign micromatrizz[78][262] = 9'b111111111;
assign micromatrizz[78][263] = 9'b111111111;
assign micromatrizz[78][264] = 9'b111111111;
assign micromatrizz[78][265] = 9'b111111111;
assign micromatrizz[78][266] = 9'b111111111;
assign micromatrizz[78][267] = 9'b111111111;
assign micromatrizz[78][268] = 9'b111111111;
assign micromatrizz[78][269] = 9'b111111111;
assign micromatrizz[78][270] = 9'b111111111;
assign micromatrizz[78][271] = 9'b111111111;
assign micromatrizz[78][272] = 9'b111111111;
assign micromatrizz[78][273] = 9'b111111111;
assign micromatrizz[78][274] = 9'b111111111;
assign micromatrizz[78][275] = 9'b111111111;
assign micromatrizz[78][276] = 9'b111111111;
assign micromatrizz[78][277] = 9'b111111111;
assign micromatrizz[78][278] = 9'b111111111;
assign micromatrizz[78][279] = 9'b111111111;
assign micromatrizz[78][280] = 9'b111111111;
assign micromatrizz[78][281] = 9'b111111111;
assign micromatrizz[78][282] = 9'b111111111;
assign micromatrizz[78][283] = 9'b111111111;
assign micromatrizz[78][284] = 9'b111111111;
assign micromatrizz[78][285] = 9'b111111111;
assign micromatrizz[78][286] = 9'b111111111;
assign micromatrizz[78][287] = 9'b111111111;
assign micromatrizz[78][288] = 9'b111111111;
assign micromatrizz[78][289] = 9'b111111111;
assign micromatrizz[78][290] = 9'b111111111;
assign micromatrizz[78][291] = 9'b111111111;
assign micromatrizz[78][292] = 9'b111111111;
assign micromatrizz[78][293] = 9'b111111111;
assign micromatrizz[78][294] = 9'b111111111;
assign micromatrizz[78][295] = 9'b111111111;
assign micromatrizz[78][296] = 9'b111111111;
assign micromatrizz[78][297] = 9'b111111111;
assign micromatrizz[78][298] = 9'b111111111;
assign micromatrizz[78][299] = 9'b111111111;
assign micromatrizz[78][300] = 9'b111111111;
assign micromatrizz[78][301] = 9'b111111111;
assign micromatrizz[78][302] = 9'b111111111;
assign micromatrizz[78][303] = 9'b111111111;
assign micromatrizz[78][304] = 9'b111111111;
assign micromatrizz[78][305] = 9'b111111111;
assign micromatrizz[78][306] = 9'b111111111;
assign micromatrizz[78][307] = 9'b111111111;
assign micromatrizz[78][308] = 9'b111111111;
assign micromatrizz[78][309] = 9'b111111111;
assign micromatrizz[78][310] = 9'b111111111;
assign micromatrizz[78][311] = 9'b111111111;
assign micromatrizz[78][312] = 9'b111111111;
assign micromatrizz[78][313] = 9'b111111111;
assign micromatrizz[78][314] = 9'b111111111;
assign micromatrizz[78][315] = 9'b111111111;
assign micromatrizz[78][316] = 9'b111111111;
assign micromatrizz[78][317] = 9'b111111111;
assign micromatrizz[78][318] = 9'b111111111;
assign micromatrizz[78][319] = 9'b111111111;
assign micromatrizz[78][320] = 9'b111111111;
assign micromatrizz[78][321] = 9'b111111111;
assign micromatrizz[78][322] = 9'b111111111;
assign micromatrizz[78][323] = 9'b111111111;
assign micromatrizz[78][324] = 9'b111111111;
assign micromatrizz[78][325] = 9'b111111111;
assign micromatrizz[78][326] = 9'b111111111;
assign micromatrizz[78][327] = 9'b111111111;
assign micromatrizz[78][328] = 9'b111111111;
assign micromatrizz[78][329] = 9'b111111111;
assign micromatrizz[78][330] = 9'b111111111;
assign micromatrizz[78][331] = 9'b111111111;
assign micromatrizz[78][332] = 9'b111111111;
assign micromatrizz[78][333] = 9'b111111111;
assign micromatrizz[78][334] = 9'b111111111;
assign micromatrizz[78][335] = 9'b111111111;
assign micromatrizz[78][336] = 9'b111111111;
assign micromatrizz[78][337] = 9'b111111111;
assign micromatrizz[78][338] = 9'b111111111;
assign micromatrizz[78][339] = 9'b111111111;
assign micromatrizz[78][340] = 9'b111111111;
assign micromatrizz[78][341] = 9'b111111111;
assign micromatrizz[78][342] = 9'b111111111;
assign micromatrizz[78][343] = 9'b111111111;
assign micromatrizz[78][344] = 9'b111111111;
assign micromatrizz[78][345] = 9'b111111111;
assign micromatrizz[78][346] = 9'b111111111;
assign micromatrizz[78][347] = 9'b111111111;
assign micromatrizz[78][348] = 9'b111111111;
assign micromatrizz[78][349] = 9'b111111111;
assign micromatrizz[78][350] = 9'b111111111;
assign micromatrizz[78][351] = 9'b111111111;
assign micromatrizz[78][352] = 9'b111111111;
assign micromatrizz[78][353] = 9'b111111111;
assign micromatrizz[78][354] = 9'b111111111;
assign micromatrizz[78][355] = 9'b111111111;
assign micromatrizz[78][356] = 9'b111111111;
assign micromatrizz[78][357] = 9'b111111111;
assign micromatrizz[78][358] = 9'b111111111;
assign micromatrizz[78][359] = 9'b111111111;
assign micromatrizz[78][360] = 9'b111111111;
assign micromatrizz[78][361] = 9'b111111111;
assign micromatrizz[78][362] = 9'b111111111;
assign micromatrizz[78][363] = 9'b111111111;
assign micromatrizz[78][364] = 9'b111111111;
assign micromatrizz[78][365] = 9'b111111111;
assign micromatrizz[78][366] = 9'b111111111;
assign micromatrizz[78][367] = 9'b111111111;
assign micromatrizz[78][368] = 9'b111111111;
assign micromatrizz[78][369] = 9'b111111111;
assign micromatrizz[78][370] = 9'b111111111;
assign micromatrizz[78][371] = 9'b111111111;
assign micromatrizz[78][372] = 9'b111111111;
assign micromatrizz[78][373] = 9'b111111111;
assign micromatrizz[78][374] = 9'b111111111;
assign micromatrizz[78][375] = 9'b111111111;
assign micromatrizz[78][376] = 9'b111111111;
assign micromatrizz[78][377] = 9'b111111111;
assign micromatrizz[78][378] = 9'b111111111;
assign micromatrizz[78][379] = 9'b111111111;
assign micromatrizz[78][380] = 9'b111111111;
assign micromatrizz[78][381] = 9'b111111111;
assign micromatrizz[78][382] = 9'b111111111;
assign micromatrizz[78][383] = 9'b111111111;
assign micromatrizz[78][384] = 9'b111111111;
assign micromatrizz[78][385] = 9'b111111111;
assign micromatrizz[78][386] = 9'b111111111;
assign micromatrizz[78][387] = 9'b111111111;
assign micromatrizz[78][388] = 9'b111111111;
assign micromatrizz[78][389] = 9'b111111111;
assign micromatrizz[78][390] = 9'b111111111;
assign micromatrizz[78][391] = 9'b111111111;
assign micromatrizz[78][392] = 9'b111111111;
assign micromatrizz[78][393] = 9'b111111111;
assign micromatrizz[78][394] = 9'b111111111;
assign micromatrizz[78][395] = 9'b111111111;
assign micromatrizz[78][396] = 9'b111111111;
assign micromatrizz[78][397] = 9'b111111111;
assign micromatrizz[78][398] = 9'b111111111;
assign micromatrizz[78][399] = 9'b111111111;
assign micromatrizz[78][400] = 9'b111111111;
assign micromatrizz[78][401] = 9'b111111111;
assign micromatrizz[78][402] = 9'b111111111;
assign micromatrizz[78][403] = 9'b111111111;
assign micromatrizz[78][404] = 9'b111111111;
assign micromatrizz[78][405] = 9'b111111111;
assign micromatrizz[78][406] = 9'b111111111;
assign micromatrizz[78][407] = 9'b111111111;
assign micromatrizz[78][408] = 9'b111111111;
assign micromatrizz[78][409] = 9'b111111111;
assign micromatrizz[78][410] = 9'b111111111;
assign micromatrizz[78][411] = 9'b111111111;
assign micromatrizz[78][412] = 9'b111111111;
assign micromatrizz[78][413] = 9'b111111111;
assign micromatrizz[78][414] = 9'b111111111;
assign micromatrizz[78][415] = 9'b111111111;
assign micromatrizz[78][416] = 9'b111111111;
assign micromatrizz[78][417] = 9'b111111111;
assign micromatrizz[78][418] = 9'b111111111;
assign micromatrizz[78][419] = 9'b111111111;
assign micromatrizz[78][420] = 9'b111111111;
assign micromatrizz[78][421] = 9'b111111111;
assign micromatrizz[78][422] = 9'b111111111;
assign micromatrizz[78][423] = 9'b111111111;
assign micromatrizz[78][424] = 9'b111111111;
assign micromatrizz[78][425] = 9'b111111111;
assign micromatrizz[78][426] = 9'b111111111;
assign micromatrizz[78][427] = 9'b111111111;
assign micromatrizz[78][428] = 9'b111111111;
assign micromatrizz[78][429] = 9'b111111111;
assign micromatrizz[78][430] = 9'b111111111;
assign micromatrizz[78][431] = 9'b111111111;
assign micromatrizz[78][432] = 9'b111111111;
assign micromatrizz[78][433] = 9'b111111111;
assign micromatrizz[78][434] = 9'b111111111;
assign micromatrizz[78][435] = 9'b111111111;
assign micromatrizz[78][436] = 9'b111111111;
assign micromatrizz[78][437] = 9'b111111111;
assign micromatrizz[78][438] = 9'b111111111;
assign micromatrizz[78][439] = 9'b111111111;
assign micromatrizz[78][440] = 9'b111111111;
assign micromatrizz[78][441] = 9'b111111111;
assign micromatrizz[78][442] = 9'b111111111;
assign micromatrizz[78][443] = 9'b111111111;
assign micromatrizz[78][444] = 9'b111111111;
assign micromatrizz[78][445] = 9'b111111111;
assign micromatrizz[78][446] = 9'b111111111;
assign micromatrizz[78][447] = 9'b111111111;
assign micromatrizz[78][448] = 9'b111111111;
assign micromatrizz[78][449] = 9'b111111111;
assign micromatrizz[78][450] = 9'b111111111;
assign micromatrizz[78][451] = 9'b111111111;
assign micromatrizz[78][452] = 9'b111111111;
assign micromatrizz[78][453] = 9'b111111111;
assign micromatrizz[78][454] = 9'b111111111;
assign micromatrizz[78][455] = 9'b111111111;
assign micromatrizz[78][456] = 9'b111111111;
assign micromatrizz[78][457] = 9'b111111111;
assign micromatrizz[78][458] = 9'b111111111;
assign micromatrizz[78][459] = 9'b111111111;
assign micromatrizz[78][460] = 9'b111111111;
assign micromatrizz[78][461] = 9'b111111111;
assign micromatrizz[78][462] = 9'b111111111;
assign micromatrizz[78][463] = 9'b111111111;
assign micromatrizz[78][464] = 9'b111111111;
assign micromatrizz[78][465] = 9'b111111111;
assign micromatrizz[78][466] = 9'b111111111;
assign micromatrizz[78][467] = 9'b111111111;
assign micromatrizz[78][468] = 9'b111111111;
assign micromatrizz[78][469] = 9'b111111111;
assign micromatrizz[78][470] = 9'b111111111;
assign micromatrizz[78][471] = 9'b111111111;
assign micromatrizz[78][472] = 9'b111111111;
assign micromatrizz[78][473] = 9'b111111111;
assign micromatrizz[78][474] = 9'b111111111;
assign micromatrizz[78][475] = 9'b111111111;
assign micromatrizz[78][476] = 9'b111111111;
assign micromatrizz[78][477] = 9'b111111111;
assign micromatrizz[78][478] = 9'b111111111;
assign micromatrizz[78][479] = 9'b111111111;
assign micromatrizz[78][480] = 9'b111111111;
assign micromatrizz[78][481] = 9'b111111111;
assign micromatrizz[78][482] = 9'b111111111;
assign micromatrizz[78][483] = 9'b111111111;
assign micromatrizz[78][484] = 9'b111111111;
assign micromatrizz[78][485] = 9'b111111111;
assign micromatrizz[78][486] = 9'b111111111;
assign micromatrizz[78][487] = 9'b111111111;
assign micromatrizz[78][488] = 9'b111111111;
assign micromatrizz[78][489] = 9'b111111111;
assign micromatrizz[78][490] = 9'b111111111;
assign micromatrizz[78][491] = 9'b111111111;
assign micromatrizz[78][492] = 9'b111111111;
assign micromatrizz[78][493] = 9'b111111111;
assign micromatrizz[78][494] = 9'b111111111;
assign micromatrizz[78][495] = 9'b111111111;
assign micromatrizz[78][496] = 9'b111111111;
assign micromatrizz[78][497] = 9'b111111111;
assign micromatrizz[78][498] = 9'b111111111;
assign micromatrizz[78][499] = 9'b111111111;
assign micromatrizz[78][500] = 9'b111111111;
assign micromatrizz[78][501] = 9'b111111111;
assign micromatrizz[78][502] = 9'b111111111;
assign micromatrizz[78][503] = 9'b111111111;
assign micromatrizz[78][504] = 9'b111111111;
assign micromatrizz[78][505] = 9'b111111111;
assign micromatrizz[78][506] = 9'b111111111;
assign micromatrizz[78][507] = 9'b111111111;
assign micromatrizz[78][508] = 9'b111111111;
assign micromatrizz[78][509] = 9'b111111111;
assign micromatrizz[78][510] = 9'b111111111;
assign micromatrizz[78][511] = 9'b111111111;
assign micromatrizz[78][512] = 9'b111111111;
assign micromatrizz[78][513] = 9'b111111111;
assign micromatrizz[78][514] = 9'b111111111;
assign micromatrizz[78][515] = 9'b111111111;
assign micromatrizz[78][516] = 9'b111111111;
assign micromatrizz[78][517] = 9'b111111111;
assign micromatrizz[78][518] = 9'b111111111;
assign micromatrizz[78][519] = 9'b111111111;
assign micromatrizz[78][520] = 9'b111111111;
assign micromatrizz[78][521] = 9'b111111111;
assign micromatrizz[78][522] = 9'b111111111;
assign micromatrizz[78][523] = 9'b111111111;
assign micromatrizz[78][524] = 9'b111111111;
assign micromatrizz[78][525] = 9'b111111111;
assign micromatrizz[78][526] = 9'b111111111;
assign micromatrizz[78][527] = 9'b111111111;
assign micromatrizz[78][528] = 9'b111111111;
assign micromatrizz[78][529] = 9'b111111111;
assign micromatrizz[78][530] = 9'b111111111;
assign micromatrizz[78][531] = 9'b111111111;
assign micromatrizz[78][532] = 9'b111111111;
assign micromatrizz[78][533] = 9'b111111111;
assign micromatrizz[78][534] = 9'b111111111;
assign micromatrizz[78][535] = 9'b111111111;
assign micromatrizz[78][536] = 9'b111111111;
assign micromatrizz[78][537] = 9'b111111111;
assign micromatrizz[78][538] = 9'b111111111;
assign micromatrizz[78][539] = 9'b111111111;
assign micromatrizz[78][540] = 9'b111111111;
assign micromatrizz[78][541] = 9'b111111111;
assign micromatrizz[78][542] = 9'b111111111;
assign micromatrizz[78][543] = 9'b111111111;
assign micromatrizz[78][544] = 9'b111111111;
assign micromatrizz[78][545] = 9'b111111111;
assign micromatrizz[78][546] = 9'b111111111;
assign micromatrizz[78][547] = 9'b111111111;
assign micromatrizz[78][548] = 9'b111111111;
assign micromatrizz[78][549] = 9'b111111111;
assign micromatrizz[78][550] = 9'b111111111;
assign micromatrizz[78][551] = 9'b111111111;
assign micromatrizz[78][552] = 9'b111111111;
assign micromatrizz[78][553] = 9'b111111111;
assign micromatrizz[78][554] = 9'b111111111;
assign micromatrizz[78][555] = 9'b111111111;
assign micromatrizz[78][556] = 9'b111111111;
assign micromatrizz[78][557] = 9'b111111111;
assign micromatrizz[78][558] = 9'b111111111;
assign micromatrizz[78][559] = 9'b111111111;
assign micromatrizz[78][560] = 9'b111111111;
assign micromatrizz[78][561] = 9'b111111111;
assign micromatrizz[78][562] = 9'b111111111;
assign micromatrizz[78][563] = 9'b111111111;
assign micromatrizz[78][564] = 9'b111111111;
assign micromatrizz[78][565] = 9'b111111111;
assign micromatrizz[78][566] = 9'b111111111;
assign micromatrizz[78][567] = 9'b111111111;
assign micromatrizz[78][568] = 9'b111111111;
assign micromatrizz[78][569] = 9'b111111111;
assign micromatrizz[78][570] = 9'b111111111;
assign micromatrizz[78][571] = 9'b111111111;
assign micromatrizz[78][572] = 9'b111111111;
assign micromatrizz[78][573] = 9'b111111111;
assign micromatrizz[78][574] = 9'b111111111;
assign micromatrizz[78][575] = 9'b111111111;
assign micromatrizz[78][576] = 9'b111111111;
assign micromatrizz[78][577] = 9'b111111111;
assign micromatrizz[78][578] = 9'b111111111;
assign micromatrizz[78][579] = 9'b111111111;
assign micromatrizz[78][580] = 9'b111111111;
assign micromatrizz[78][581] = 9'b111111111;
assign micromatrizz[78][582] = 9'b111111111;
assign micromatrizz[78][583] = 9'b111111111;
assign micromatrizz[78][584] = 9'b111111111;
assign micromatrizz[78][585] = 9'b111111111;
assign micromatrizz[78][586] = 9'b111111111;
assign micromatrizz[78][587] = 9'b111111111;
assign micromatrizz[78][588] = 9'b111111111;
assign micromatrizz[78][589] = 9'b111111111;
assign micromatrizz[78][590] = 9'b111111111;
assign micromatrizz[78][591] = 9'b111111111;
assign micromatrizz[78][592] = 9'b111111111;
assign micromatrizz[78][593] = 9'b111111111;
assign micromatrizz[78][594] = 9'b111111111;
assign micromatrizz[78][595] = 9'b111111111;
assign micromatrizz[78][596] = 9'b111111111;
assign micromatrizz[78][597] = 9'b111111111;
assign micromatrizz[78][598] = 9'b111111111;
assign micromatrizz[78][599] = 9'b111111111;
assign micromatrizz[78][600] = 9'b111111111;
assign micromatrizz[78][601] = 9'b111111111;
assign micromatrizz[78][602] = 9'b111111111;
assign micromatrizz[78][603] = 9'b111111111;
assign micromatrizz[78][604] = 9'b111111111;
assign micromatrizz[78][605] = 9'b111111111;
assign micromatrizz[78][606] = 9'b111111111;
assign micromatrizz[78][607] = 9'b111111111;
assign micromatrizz[78][608] = 9'b111111111;
assign micromatrizz[78][609] = 9'b111111111;
assign micromatrizz[78][610] = 9'b111111111;
assign micromatrizz[78][611] = 9'b111111111;
assign micromatrizz[78][612] = 9'b111111111;
assign micromatrizz[78][613] = 9'b111111111;
assign micromatrizz[78][614] = 9'b111111111;
assign micromatrizz[78][615] = 9'b111111111;
assign micromatrizz[78][616] = 9'b111111111;
assign micromatrizz[78][617] = 9'b111111111;
assign micromatrizz[78][618] = 9'b111111111;
assign micromatrizz[78][619] = 9'b111111111;
assign micromatrizz[78][620] = 9'b111111111;
assign micromatrizz[78][621] = 9'b111111111;
assign micromatrizz[78][622] = 9'b111111111;
assign micromatrizz[78][623] = 9'b111111111;
assign micromatrizz[78][624] = 9'b111111111;
assign micromatrizz[78][625] = 9'b111111111;
assign micromatrizz[78][626] = 9'b111111111;
assign micromatrizz[78][627] = 9'b111111111;
assign micromatrizz[78][628] = 9'b111111111;
assign micromatrizz[78][629] = 9'b111111111;
assign micromatrizz[78][630] = 9'b111111111;
assign micromatrizz[78][631] = 9'b111111111;
assign micromatrizz[78][632] = 9'b111111111;
assign micromatrizz[78][633] = 9'b111111111;
assign micromatrizz[78][634] = 9'b111111111;
assign micromatrizz[78][635] = 9'b111111111;
assign micromatrizz[78][636] = 9'b111111111;
assign micromatrizz[78][637] = 9'b111111111;
assign micromatrizz[78][638] = 9'b111111111;
assign micromatrizz[78][639] = 9'b111111111;
assign micromatrizz[79][0] = 9'b111111111;
assign micromatrizz[79][1] = 9'b111111111;
assign micromatrizz[79][2] = 9'b111111111;
assign micromatrizz[79][3] = 9'b111111111;
assign micromatrizz[79][4] = 9'b111111111;
assign micromatrizz[79][5] = 9'b111111111;
assign micromatrizz[79][6] = 9'b111111111;
assign micromatrizz[79][7] = 9'b111111111;
assign micromatrizz[79][8] = 9'b111111111;
assign micromatrizz[79][9] = 9'b111111111;
assign micromatrizz[79][10] = 9'b111111111;
assign micromatrizz[79][11] = 9'b111111111;
assign micromatrizz[79][12] = 9'b111111111;
assign micromatrizz[79][13] = 9'b111111111;
assign micromatrizz[79][14] = 9'b111111111;
assign micromatrizz[79][15] = 9'b111111111;
assign micromatrizz[79][16] = 9'b111111111;
assign micromatrizz[79][17] = 9'b111111111;
assign micromatrizz[79][18] = 9'b111111111;
assign micromatrizz[79][19] = 9'b111111111;
assign micromatrizz[79][20] = 9'b111111111;
assign micromatrizz[79][21] = 9'b111111111;
assign micromatrizz[79][22] = 9'b111111111;
assign micromatrizz[79][23] = 9'b111111111;
assign micromatrizz[79][24] = 9'b111111111;
assign micromatrizz[79][25] = 9'b111111111;
assign micromatrizz[79][26] = 9'b111111111;
assign micromatrizz[79][27] = 9'b111111111;
assign micromatrizz[79][28] = 9'b111111111;
assign micromatrizz[79][29] = 9'b111111111;
assign micromatrizz[79][30] = 9'b111111111;
assign micromatrizz[79][31] = 9'b111111111;
assign micromatrizz[79][32] = 9'b111111111;
assign micromatrizz[79][33] = 9'b111111111;
assign micromatrizz[79][34] = 9'b111111111;
assign micromatrizz[79][35] = 9'b111111111;
assign micromatrizz[79][36] = 9'b111111111;
assign micromatrizz[79][37] = 9'b111111111;
assign micromatrizz[79][38] = 9'b111111111;
assign micromatrizz[79][39] = 9'b111111111;
assign micromatrizz[79][40] = 9'b111111111;
assign micromatrizz[79][41] = 9'b111111111;
assign micromatrizz[79][42] = 9'b111111111;
assign micromatrizz[79][43] = 9'b111111111;
assign micromatrizz[79][44] = 9'b111111111;
assign micromatrizz[79][45] = 9'b111111111;
assign micromatrizz[79][46] = 9'b111111111;
assign micromatrizz[79][47] = 9'b111111111;
assign micromatrizz[79][48] = 9'b111111111;
assign micromatrizz[79][49] = 9'b111111111;
assign micromatrizz[79][50] = 9'b111111111;
assign micromatrizz[79][51] = 9'b111111111;
assign micromatrizz[79][52] = 9'b111111111;
assign micromatrizz[79][53] = 9'b111111111;
assign micromatrizz[79][54] = 9'b111111111;
assign micromatrizz[79][55] = 9'b111111111;
assign micromatrizz[79][56] = 9'b111111111;
assign micromatrizz[79][57] = 9'b111111111;
assign micromatrizz[79][58] = 9'b111111111;
assign micromatrizz[79][59] = 9'b111111111;
assign micromatrizz[79][60] = 9'b111111111;
assign micromatrizz[79][61] = 9'b111111111;
assign micromatrizz[79][62] = 9'b111111111;
assign micromatrizz[79][63] = 9'b111111111;
assign micromatrizz[79][64] = 9'b111111111;
assign micromatrizz[79][65] = 9'b111111111;
assign micromatrizz[79][66] = 9'b111111111;
assign micromatrizz[79][67] = 9'b111111111;
assign micromatrizz[79][68] = 9'b111111111;
assign micromatrizz[79][69] = 9'b111111111;
assign micromatrizz[79][70] = 9'b111111111;
assign micromatrizz[79][71] = 9'b111111111;
assign micromatrizz[79][72] = 9'b111111111;
assign micromatrizz[79][73] = 9'b111111111;
assign micromatrizz[79][74] = 9'b111111111;
assign micromatrizz[79][75] = 9'b111111111;
assign micromatrizz[79][76] = 9'b111111111;
assign micromatrizz[79][77] = 9'b111111111;
assign micromatrizz[79][78] = 9'b111111111;
assign micromatrizz[79][79] = 9'b111111111;
assign micromatrizz[79][80] = 9'b111111111;
assign micromatrizz[79][81] = 9'b111111111;
assign micromatrizz[79][82] = 9'b111111111;
assign micromatrizz[79][83] = 9'b111111111;
assign micromatrizz[79][84] = 9'b111111111;
assign micromatrizz[79][85] = 9'b111111111;
assign micromatrizz[79][86] = 9'b111111111;
assign micromatrizz[79][87] = 9'b111111111;
assign micromatrizz[79][88] = 9'b111111111;
assign micromatrizz[79][89] = 9'b111111111;
assign micromatrizz[79][90] = 9'b111111111;
assign micromatrizz[79][91] = 9'b111111111;
assign micromatrizz[79][92] = 9'b111111111;
assign micromatrizz[79][93] = 9'b111111111;
assign micromatrizz[79][94] = 9'b111111111;
assign micromatrizz[79][95] = 9'b111111111;
assign micromatrizz[79][96] = 9'b111111111;
assign micromatrizz[79][97] = 9'b111111111;
assign micromatrizz[79][98] = 9'b111111111;
assign micromatrizz[79][99] = 9'b111111111;
assign micromatrizz[79][100] = 9'b111111111;
assign micromatrizz[79][101] = 9'b111111111;
assign micromatrizz[79][102] = 9'b111111111;
assign micromatrizz[79][103] = 9'b111111111;
assign micromatrizz[79][104] = 9'b111111111;
assign micromatrizz[79][105] = 9'b111111111;
assign micromatrizz[79][106] = 9'b111111111;
assign micromatrizz[79][107] = 9'b111111111;
assign micromatrizz[79][108] = 9'b111111111;
assign micromatrizz[79][109] = 9'b111111111;
assign micromatrizz[79][110] = 9'b111111111;
assign micromatrizz[79][111] = 9'b111111111;
assign micromatrizz[79][112] = 9'b111111111;
assign micromatrizz[79][113] = 9'b111111111;
assign micromatrizz[79][114] = 9'b111111111;
assign micromatrizz[79][115] = 9'b111111111;
assign micromatrizz[79][116] = 9'b111111111;
assign micromatrizz[79][117] = 9'b111111111;
assign micromatrizz[79][118] = 9'b111111111;
assign micromatrizz[79][119] = 9'b111111111;
assign micromatrizz[79][120] = 9'b111111111;
assign micromatrizz[79][121] = 9'b111111111;
assign micromatrizz[79][122] = 9'b111111111;
assign micromatrizz[79][123] = 9'b111111111;
assign micromatrizz[79][124] = 9'b111111111;
assign micromatrizz[79][125] = 9'b111111111;
assign micromatrizz[79][126] = 9'b111111111;
assign micromatrizz[79][127] = 9'b111111111;
assign micromatrizz[79][128] = 9'b111111111;
assign micromatrizz[79][129] = 9'b111111111;
assign micromatrizz[79][130] = 9'b111111111;
assign micromatrizz[79][131] = 9'b111111111;
assign micromatrizz[79][132] = 9'b111111111;
assign micromatrizz[79][133] = 9'b111111111;
assign micromatrizz[79][134] = 9'b111111111;
assign micromatrizz[79][135] = 9'b111111111;
assign micromatrizz[79][136] = 9'b111111111;
assign micromatrizz[79][137] = 9'b111111111;
assign micromatrizz[79][138] = 9'b111111111;
assign micromatrizz[79][139] = 9'b111111111;
assign micromatrizz[79][140] = 9'b111111111;
assign micromatrizz[79][141] = 9'b111111111;
assign micromatrizz[79][142] = 9'b111111111;
assign micromatrizz[79][143] = 9'b111111111;
assign micromatrizz[79][144] = 9'b111111111;
assign micromatrizz[79][145] = 9'b111111111;
assign micromatrizz[79][146] = 9'b111111111;
assign micromatrizz[79][147] = 9'b111111111;
assign micromatrizz[79][148] = 9'b111111111;
assign micromatrizz[79][149] = 9'b111111111;
assign micromatrizz[79][150] = 9'b111111111;
assign micromatrizz[79][151] = 9'b111111111;
assign micromatrizz[79][152] = 9'b111111111;
assign micromatrizz[79][153] = 9'b111111111;
assign micromatrizz[79][154] = 9'b111111111;
assign micromatrizz[79][155] = 9'b111111111;
assign micromatrizz[79][156] = 9'b111111111;
assign micromatrizz[79][157] = 9'b111111111;
assign micromatrizz[79][158] = 9'b111111111;
assign micromatrizz[79][159] = 9'b111111111;
assign micromatrizz[79][160] = 9'b111111111;
assign micromatrizz[79][161] = 9'b111111111;
assign micromatrizz[79][162] = 9'b111111111;
assign micromatrizz[79][163] = 9'b111111111;
assign micromatrizz[79][164] = 9'b111111111;
assign micromatrizz[79][165] = 9'b111111111;
assign micromatrizz[79][166] = 9'b111111111;
assign micromatrizz[79][167] = 9'b111111111;
assign micromatrizz[79][168] = 9'b111111111;
assign micromatrizz[79][169] = 9'b111111111;
assign micromatrizz[79][170] = 9'b111111111;
assign micromatrizz[79][171] = 9'b111111111;
assign micromatrizz[79][172] = 9'b111111111;
assign micromatrizz[79][173] = 9'b111111111;
assign micromatrizz[79][174] = 9'b111111111;
assign micromatrizz[79][175] = 9'b111111111;
assign micromatrizz[79][176] = 9'b111111111;
assign micromatrizz[79][177] = 9'b111111111;
assign micromatrizz[79][178] = 9'b111111111;
assign micromatrizz[79][179] = 9'b111111111;
assign micromatrizz[79][180] = 9'b111111111;
assign micromatrizz[79][181] = 9'b111111111;
assign micromatrizz[79][182] = 9'b111111111;
assign micromatrizz[79][183] = 9'b111111111;
assign micromatrizz[79][184] = 9'b111111111;
assign micromatrizz[79][185] = 9'b111111111;
assign micromatrizz[79][186] = 9'b111111111;
assign micromatrizz[79][187] = 9'b111111111;
assign micromatrizz[79][188] = 9'b111111111;
assign micromatrizz[79][189] = 9'b111111111;
assign micromatrizz[79][190] = 9'b111111111;
assign micromatrizz[79][191] = 9'b111111111;
assign micromatrizz[79][192] = 9'b111111111;
assign micromatrizz[79][193] = 9'b111111111;
assign micromatrizz[79][194] = 9'b111111111;
assign micromatrizz[79][195] = 9'b111111111;
assign micromatrizz[79][196] = 9'b111111111;
assign micromatrizz[79][197] = 9'b111111111;
assign micromatrizz[79][198] = 9'b111111111;
assign micromatrizz[79][199] = 9'b111111111;
assign micromatrizz[79][200] = 9'b111111111;
assign micromatrizz[79][201] = 9'b111111111;
assign micromatrizz[79][202] = 9'b111111111;
assign micromatrizz[79][203] = 9'b111111111;
assign micromatrizz[79][204] = 9'b111111111;
assign micromatrizz[79][205] = 9'b111111111;
assign micromatrizz[79][206] = 9'b111111111;
assign micromatrizz[79][207] = 9'b111111111;
assign micromatrizz[79][208] = 9'b111111111;
assign micromatrizz[79][209] = 9'b111111111;
assign micromatrizz[79][210] = 9'b111111111;
assign micromatrizz[79][211] = 9'b111111111;
assign micromatrizz[79][212] = 9'b111111111;
assign micromatrizz[79][213] = 9'b111111111;
assign micromatrizz[79][214] = 9'b111111111;
assign micromatrizz[79][215] = 9'b111111111;
assign micromatrizz[79][216] = 9'b111111111;
assign micromatrizz[79][217] = 9'b111111111;
assign micromatrizz[79][218] = 9'b111111111;
assign micromatrizz[79][219] = 9'b111111111;
assign micromatrizz[79][220] = 9'b111111111;
assign micromatrizz[79][221] = 9'b111111111;
assign micromatrizz[79][222] = 9'b111111111;
assign micromatrizz[79][223] = 9'b111111111;
assign micromatrizz[79][224] = 9'b111111111;
assign micromatrizz[79][225] = 9'b111111111;
assign micromatrizz[79][226] = 9'b111111111;
assign micromatrizz[79][227] = 9'b111111111;
assign micromatrizz[79][228] = 9'b111111111;
assign micromatrizz[79][229] = 9'b111111111;
assign micromatrizz[79][230] = 9'b111111111;
assign micromatrizz[79][231] = 9'b111111111;
assign micromatrizz[79][232] = 9'b111111111;
assign micromatrizz[79][233] = 9'b111111111;
assign micromatrizz[79][234] = 9'b111111111;
assign micromatrizz[79][235] = 9'b111111111;
assign micromatrizz[79][236] = 9'b111111111;
assign micromatrizz[79][237] = 9'b111111111;
assign micromatrizz[79][238] = 9'b111111111;
assign micromatrizz[79][239] = 9'b111111111;
assign micromatrizz[79][240] = 9'b111111111;
assign micromatrizz[79][241] = 9'b111111111;
assign micromatrizz[79][242] = 9'b111111111;
assign micromatrizz[79][243] = 9'b111111111;
assign micromatrizz[79][244] = 9'b111111111;
assign micromatrizz[79][245] = 9'b111111111;
assign micromatrizz[79][246] = 9'b111111111;
assign micromatrizz[79][247] = 9'b111111111;
assign micromatrizz[79][248] = 9'b111111111;
assign micromatrizz[79][249] = 9'b111111111;
assign micromatrizz[79][250] = 9'b111111111;
assign micromatrizz[79][251] = 9'b111111111;
assign micromatrizz[79][252] = 9'b111111111;
assign micromatrizz[79][253] = 9'b111111111;
assign micromatrizz[79][254] = 9'b111111111;
assign micromatrizz[79][255] = 9'b111111111;
assign micromatrizz[79][256] = 9'b111111111;
assign micromatrizz[79][257] = 9'b111111111;
assign micromatrizz[79][258] = 9'b111111111;
assign micromatrizz[79][259] = 9'b111111111;
assign micromatrizz[79][260] = 9'b111111111;
assign micromatrizz[79][261] = 9'b111111111;
assign micromatrizz[79][262] = 9'b111111111;
assign micromatrizz[79][263] = 9'b111111111;
assign micromatrizz[79][264] = 9'b111111111;
assign micromatrizz[79][265] = 9'b111111111;
assign micromatrizz[79][266] = 9'b111111111;
assign micromatrizz[79][267] = 9'b111111111;
assign micromatrizz[79][268] = 9'b111111111;
assign micromatrizz[79][269] = 9'b111111111;
assign micromatrizz[79][270] = 9'b111111111;
assign micromatrizz[79][271] = 9'b111111111;
assign micromatrizz[79][272] = 9'b111111111;
assign micromatrizz[79][273] = 9'b111111111;
assign micromatrizz[79][274] = 9'b111111111;
assign micromatrizz[79][275] = 9'b111111111;
assign micromatrizz[79][276] = 9'b111111111;
assign micromatrizz[79][277] = 9'b111111111;
assign micromatrizz[79][278] = 9'b111111111;
assign micromatrizz[79][279] = 9'b111111111;
assign micromatrizz[79][280] = 9'b111111111;
assign micromatrizz[79][281] = 9'b111111111;
assign micromatrizz[79][282] = 9'b111111111;
assign micromatrizz[79][283] = 9'b111111111;
assign micromatrizz[79][284] = 9'b111111111;
assign micromatrizz[79][285] = 9'b111111111;
assign micromatrizz[79][286] = 9'b111111111;
assign micromatrizz[79][287] = 9'b111111111;
assign micromatrizz[79][288] = 9'b111111111;
assign micromatrizz[79][289] = 9'b111111111;
assign micromatrizz[79][290] = 9'b111111111;
assign micromatrizz[79][291] = 9'b111111111;
assign micromatrizz[79][292] = 9'b111111111;
assign micromatrizz[79][293] = 9'b111111111;
assign micromatrizz[79][294] = 9'b111111111;
assign micromatrizz[79][295] = 9'b111111111;
assign micromatrizz[79][296] = 9'b111111111;
assign micromatrizz[79][297] = 9'b111111111;
assign micromatrizz[79][298] = 9'b111111111;
assign micromatrizz[79][299] = 9'b111111111;
assign micromatrizz[79][300] = 9'b111111111;
assign micromatrizz[79][301] = 9'b111111111;
assign micromatrizz[79][302] = 9'b111111111;
assign micromatrizz[79][303] = 9'b111111111;
assign micromatrizz[79][304] = 9'b111111111;
assign micromatrizz[79][305] = 9'b111111111;
assign micromatrizz[79][306] = 9'b111111111;
assign micromatrizz[79][307] = 9'b111111111;
assign micromatrizz[79][308] = 9'b111111111;
assign micromatrizz[79][309] = 9'b111111111;
assign micromatrizz[79][310] = 9'b111111111;
assign micromatrizz[79][311] = 9'b111111111;
assign micromatrizz[79][312] = 9'b111111111;
assign micromatrizz[79][313] = 9'b111111111;
assign micromatrizz[79][314] = 9'b111111111;
assign micromatrizz[79][315] = 9'b111111111;
assign micromatrizz[79][316] = 9'b111111111;
assign micromatrizz[79][317] = 9'b111111111;
assign micromatrizz[79][318] = 9'b111111111;
assign micromatrizz[79][319] = 9'b111111111;
assign micromatrizz[79][320] = 9'b111111111;
assign micromatrizz[79][321] = 9'b111111111;
assign micromatrizz[79][322] = 9'b111111111;
assign micromatrizz[79][323] = 9'b111111111;
assign micromatrizz[79][324] = 9'b111111111;
assign micromatrizz[79][325] = 9'b111111111;
assign micromatrizz[79][326] = 9'b111111111;
assign micromatrizz[79][327] = 9'b111111111;
assign micromatrizz[79][328] = 9'b111111111;
assign micromatrizz[79][329] = 9'b111111111;
assign micromatrizz[79][330] = 9'b111111111;
assign micromatrizz[79][331] = 9'b111111111;
assign micromatrizz[79][332] = 9'b111111111;
assign micromatrizz[79][333] = 9'b111111111;
assign micromatrizz[79][334] = 9'b111111111;
assign micromatrizz[79][335] = 9'b111111111;
assign micromatrizz[79][336] = 9'b111111111;
assign micromatrizz[79][337] = 9'b111111111;
assign micromatrizz[79][338] = 9'b111111111;
assign micromatrizz[79][339] = 9'b111111111;
assign micromatrizz[79][340] = 9'b111111111;
assign micromatrizz[79][341] = 9'b111111111;
assign micromatrizz[79][342] = 9'b111111111;
assign micromatrizz[79][343] = 9'b111111111;
assign micromatrizz[79][344] = 9'b111111111;
assign micromatrizz[79][345] = 9'b111111111;
assign micromatrizz[79][346] = 9'b111111111;
assign micromatrizz[79][347] = 9'b111111111;
assign micromatrizz[79][348] = 9'b111111111;
assign micromatrizz[79][349] = 9'b111111111;
assign micromatrizz[79][350] = 9'b111111111;
assign micromatrizz[79][351] = 9'b111111111;
assign micromatrizz[79][352] = 9'b111111111;
assign micromatrizz[79][353] = 9'b111111111;
assign micromatrizz[79][354] = 9'b111111111;
assign micromatrizz[79][355] = 9'b111111111;
assign micromatrizz[79][356] = 9'b111111111;
assign micromatrizz[79][357] = 9'b111111111;
assign micromatrizz[79][358] = 9'b111111111;
assign micromatrizz[79][359] = 9'b111111111;
assign micromatrizz[79][360] = 9'b111111111;
assign micromatrizz[79][361] = 9'b111111111;
assign micromatrizz[79][362] = 9'b111111111;
assign micromatrizz[79][363] = 9'b111111111;
assign micromatrizz[79][364] = 9'b111111111;
assign micromatrizz[79][365] = 9'b111111111;
assign micromatrizz[79][366] = 9'b111111111;
assign micromatrizz[79][367] = 9'b111111111;
assign micromatrizz[79][368] = 9'b111111111;
assign micromatrizz[79][369] = 9'b111111111;
assign micromatrizz[79][370] = 9'b111111111;
assign micromatrizz[79][371] = 9'b111111111;
assign micromatrizz[79][372] = 9'b111111111;
assign micromatrizz[79][373] = 9'b111111111;
assign micromatrizz[79][374] = 9'b111111111;
assign micromatrizz[79][375] = 9'b111111111;
assign micromatrizz[79][376] = 9'b111111111;
assign micromatrizz[79][377] = 9'b111111111;
assign micromatrizz[79][378] = 9'b111111111;
assign micromatrizz[79][379] = 9'b111111111;
assign micromatrizz[79][380] = 9'b111111111;
assign micromatrizz[79][381] = 9'b111111111;
assign micromatrizz[79][382] = 9'b111111111;
assign micromatrizz[79][383] = 9'b111111111;
assign micromatrizz[79][384] = 9'b111111111;
assign micromatrizz[79][385] = 9'b111111111;
assign micromatrizz[79][386] = 9'b111111111;
assign micromatrizz[79][387] = 9'b111111111;
assign micromatrizz[79][388] = 9'b111111111;
assign micromatrizz[79][389] = 9'b111111111;
assign micromatrizz[79][390] = 9'b111111111;
assign micromatrizz[79][391] = 9'b111111111;
assign micromatrizz[79][392] = 9'b111111111;
assign micromatrizz[79][393] = 9'b111111111;
assign micromatrizz[79][394] = 9'b111111111;
assign micromatrizz[79][395] = 9'b111111111;
assign micromatrizz[79][396] = 9'b111111111;
assign micromatrizz[79][397] = 9'b111111111;
assign micromatrizz[79][398] = 9'b111111111;
assign micromatrizz[79][399] = 9'b111111111;
assign micromatrizz[79][400] = 9'b111111111;
assign micromatrizz[79][401] = 9'b111111111;
assign micromatrizz[79][402] = 9'b111111111;
assign micromatrizz[79][403] = 9'b111111111;
assign micromatrizz[79][404] = 9'b111111111;
assign micromatrizz[79][405] = 9'b111111111;
assign micromatrizz[79][406] = 9'b111111111;
assign micromatrizz[79][407] = 9'b111111111;
assign micromatrizz[79][408] = 9'b111111111;
assign micromatrizz[79][409] = 9'b111111111;
assign micromatrizz[79][410] = 9'b111111111;
assign micromatrizz[79][411] = 9'b111111111;
assign micromatrizz[79][412] = 9'b111111111;
assign micromatrizz[79][413] = 9'b111111111;
assign micromatrizz[79][414] = 9'b111111111;
assign micromatrizz[79][415] = 9'b111111111;
assign micromatrizz[79][416] = 9'b111111111;
assign micromatrizz[79][417] = 9'b111111111;
assign micromatrizz[79][418] = 9'b111111111;
assign micromatrizz[79][419] = 9'b111111111;
assign micromatrizz[79][420] = 9'b111111111;
assign micromatrizz[79][421] = 9'b111111111;
assign micromatrizz[79][422] = 9'b111111111;
assign micromatrizz[79][423] = 9'b111111111;
assign micromatrizz[79][424] = 9'b111111111;
assign micromatrizz[79][425] = 9'b111111111;
assign micromatrizz[79][426] = 9'b111111111;
assign micromatrizz[79][427] = 9'b111111111;
assign micromatrizz[79][428] = 9'b111111111;
assign micromatrizz[79][429] = 9'b111111111;
assign micromatrizz[79][430] = 9'b111111111;
assign micromatrizz[79][431] = 9'b111111111;
assign micromatrizz[79][432] = 9'b111111111;
assign micromatrizz[79][433] = 9'b111111111;
assign micromatrizz[79][434] = 9'b111111111;
assign micromatrizz[79][435] = 9'b111111111;
assign micromatrizz[79][436] = 9'b111111111;
assign micromatrizz[79][437] = 9'b111111111;
assign micromatrizz[79][438] = 9'b111111111;
assign micromatrizz[79][439] = 9'b111111111;
assign micromatrizz[79][440] = 9'b111111111;
assign micromatrizz[79][441] = 9'b111111111;
assign micromatrizz[79][442] = 9'b111111111;
assign micromatrizz[79][443] = 9'b111111111;
assign micromatrizz[79][444] = 9'b111111111;
assign micromatrizz[79][445] = 9'b111111111;
assign micromatrizz[79][446] = 9'b111111111;
assign micromatrizz[79][447] = 9'b111111111;
assign micromatrizz[79][448] = 9'b111111111;
assign micromatrizz[79][449] = 9'b111111111;
assign micromatrizz[79][450] = 9'b111111111;
assign micromatrizz[79][451] = 9'b111111111;
assign micromatrizz[79][452] = 9'b111111111;
assign micromatrizz[79][453] = 9'b111111111;
assign micromatrizz[79][454] = 9'b111111111;
assign micromatrizz[79][455] = 9'b111111111;
assign micromatrizz[79][456] = 9'b111111111;
assign micromatrizz[79][457] = 9'b111111111;
assign micromatrizz[79][458] = 9'b111111111;
assign micromatrizz[79][459] = 9'b111111111;
assign micromatrizz[79][460] = 9'b111111111;
assign micromatrizz[79][461] = 9'b111111111;
assign micromatrizz[79][462] = 9'b111111111;
assign micromatrizz[79][463] = 9'b111111111;
assign micromatrizz[79][464] = 9'b111111111;
assign micromatrizz[79][465] = 9'b111111111;
assign micromatrizz[79][466] = 9'b111111111;
assign micromatrizz[79][467] = 9'b111111111;
assign micromatrizz[79][468] = 9'b111111111;
assign micromatrizz[79][469] = 9'b111111111;
assign micromatrizz[79][470] = 9'b111111111;
assign micromatrizz[79][471] = 9'b111111111;
assign micromatrizz[79][472] = 9'b111111111;
assign micromatrizz[79][473] = 9'b111111111;
assign micromatrizz[79][474] = 9'b111111111;
assign micromatrizz[79][475] = 9'b111111111;
assign micromatrizz[79][476] = 9'b111111111;
assign micromatrizz[79][477] = 9'b111111111;
assign micromatrizz[79][478] = 9'b111111111;
assign micromatrizz[79][479] = 9'b111111111;
assign micromatrizz[79][480] = 9'b111111111;
assign micromatrizz[79][481] = 9'b111111111;
assign micromatrizz[79][482] = 9'b111111111;
assign micromatrizz[79][483] = 9'b111111111;
assign micromatrizz[79][484] = 9'b111111111;
assign micromatrizz[79][485] = 9'b111111111;
assign micromatrizz[79][486] = 9'b111111111;
assign micromatrizz[79][487] = 9'b111111111;
assign micromatrizz[79][488] = 9'b111111111;
assign micromatrizz[79][489] = 9'b111111111;
assign micromatrizz[79][490] = 9'b111111111;
assign micromatrizz[79][491] = 9'b111111111;
assign micromatrizz[79][492] = 9'b111111111;
assign micromatrizz[79][493] = 9'b111111111;
assign micromatrizz[79][494] = 9'b111111111;
assign micromatrizz[79][495] = 9'b111111111;
assign micromatrizz[79][496] = 9'b111111111;
assign micromatrizz[79][497] = 9'b111111111;
assign micromatrizz[79][498] = 9'b111111111;
assign micromatrizz[79][499] = 9'b111111111;
assign micromatrizz[79][500] = 9'b111111111;
assign micromatrizz[79][501] = 9'b111111111;
assign micromatrizz[79][502] = 9'b111111111;
assign micromatrizz[79][503] = 9'b111111111;
assign micromatrizz[79][504] = 9'b111111111;
assign micromatrizz[79][505] = 9'b111111111;
assign micromatrizz[79][506] = 9'b111111111;
assign micromatrizz[79][507] = 9'b111111111;
assign micromatrizz[79][508] = 9'b111111111;
assign micromatrizz[79][509] = 9'b111111111;
assign micromatrizz[79][510] = 9'b111111111;
assign micromatrizz[79][511] = 9'b111111111;
assign micromatrizz[79][512] = 9'b111111111;
assign micromatrizz[79][513] = 9'b111111111;
assign micromatrizz[79][514] = 9'b111111111;
assign micromatrizz[79][515] = 9'b111111111;
assign micromatrizz[79][516] = 9'b111111111;
assign micromatrizz[79][517] = 9'b111111111;
assign micromatrizz[79][518] = 9'b111111111;
assign micromatrizz[79][519] = 9'b111111111;
assign micromatrizz[79][520] = 9'b111111111;
assign micromatrizz[79][521] = 9'b111111111;
assign micromatrizz[79][522] = 9'b111111111;
assign micromatrizz[79][523] = 9'b111111111;
assign micromatrizz[79][524] = 9'b111111111;
assign micromatrizz[79][525] = 9'b111111111;
assign micromatrizz[79][526] = 9'b111111111;
assign micromatrizz[79][527] = 9'b111111111;
assign micromatrizz[79][528] = 9'b111111111;
assign micromatrizz[79][529] = 9'b111111111;
assign micromatrizz[79][530] = 9'b111111111;
assign micromatrizz[79][531] = 9'b111111111;
assign micromatrizz[79][532] = 9'b111111111;
assign micromatrizz[79][533] = 9'b111111111;
assign micromatrizz[79][534] = 9'b111111111;
assign micromatrizz[79][535] = 9'b111111111;
assign micromatrizz[79][536] = 9'b111111111;
assign micromatrizz[79][537] = 9'b111111111;
assign micromatrizz[79][538] = 9'b111111111;
assign micromatrizz[79][539] = 9'b111111111;
assign micromatrizz[79][540] = 9'b111111111;
assign micromatrizz[79][541] = 9'b111111111;
assign micromatrizz[79][542] = 9'b111111111;
assign micromatrizz[79][543] = 9'b111111111;
assign micromatrizz[79][544] = 9'b111111111;
assign micromatrizz[79][545] = 9'b111111111;
assign micromatrizz[79][546] = 9'b111111111;
assign micromatrizz[79][547] = 9'b111111111;
assign micromatrizz[79][548] = 9'b111111111;
assign micromatrizz[79][549] = 9'b111111111;
assign micromatrizz[79][550] = 9'b111111111;
assign micromatrizz[79][551] = 9'b111111111;
assign micromatrizz[79][552] = 9'b111111111;
assign micromatrizz[79][553] = 9'b111111111;
assign micromatrizz[79][554] = 9'b111111111;
assign micromatrizz[79][555] = 9'b111111111;
assign micromatrizz[79][556] = 9'b111111111;
assign micromatrizz[79][557] = 9'b111111111;
assign micromatrizz[79][558] = 9'b111111111;
assign micromatrizz[79][559] = 9'b111111111;
assign micromatrizz[79][560] = 9'b111111111;
assign micromatrizz[79][561] = 9'b111111111;
assign micromatrizz[79][562] = 9'b111111111;
assign micromatrizz[79][563] = 9'b111111111;
assign micromatrizz[79][564] = 9'b111111111;
assign micromatrizz[79][565] = 9'b111111111;
assign micromatrizz[79][566] = 9'b111111111;
assign micromatrizz[79][567] = 9'b111111111;
assign micromatrizz[79][568] = 9'b111111111;
assign micromatrizz[79][569] = 9'b111111111;
assign micromatrizz[79][570] = 9'b111111111;
assign micromatrizz[79][571] = 9'b111111111;
assign micromatrizz[79][572] = 9'b111111111;
assign micromatrizz[79][573] = 9'b111111111;
assign micromatrizz[79][574] = 9'b111111111;
assign micromatrizz[79][575] = 9'b111111111;
assign micromatrizz[79][576] = 9'b111111111;
assign micromatrizz[79][577] = 9'b111111111;
assign micromatrizz[79][578] = 9'b111111111;
assign micromatrizz[79][579] = 9'b111111111;
assign micromatrizz[79][580] = 9'b111111111;
assign micromatrizz[79][581] = 9'b111111111;
assign micromatrizz[79][582] = 9'b111111111;
assign micromatrizz[79][583] = 9'b111111111;
assign micromatrizz[79][584] = 9'b111111111;
assign micromatrizz[79][585] = 9'b111111111;
assign micromatrizz[79][586] = 9'b111111111;
assign micromatrizz[79][587] = 9'b111111111;
assign micromatrizz[79][588] = 9'b111111111;
assign micromatrizz[79][589] = 9'b111111111;
assign micromatrizz[79][590] = 9'b111111111;
assign micromatrizz[79][591] = 9'b111111111;
assign micromatrizz[79][592] = 9'b111111111;
assign micromatrizz[79][593] = 9'b111111111;
assign micromatrizz[79][594] = 9'b111111111;
assign micromatrizz[79][595] = 9'b111111111;
assign micromatrizz[79][596] = 9'b111111111;
assign micromatrizz[79][597] = 9'b111111111;
assign micromatrizz[79][598] = 9'b111111111;
assign micromatrizz[79][599] = 9'b111111111;
assign micromatrizz[79][600] = 9'b111111111;
assign micromatrizz[79][601] = 9'b111111111;
assign micromatrizz[79][602] = 9'b111111111;
assign micromatrizz[79][603] = 9'b111111111;
assign micromatrizz[79][604] = 9'b111111111;
assign micromatrizz[79][605] = 9'b111111111;
assign micromatrizz[79][606] = 9'b111111111;
assign micromatrizz[79][607] = 9'b111111111;
assign micromatrizz[79][608] = 9'b111111111;
assign micromatrizz[79][609] = 9'b111111111;
assign micromatrizz[79][610] = 9'b111111111;
assign micromatrizz[79][611] = 9'b111111111;
assign micromatrizz[79][612] = 9'b111111111;
assign micromatrizz[79][613] = 9'b111111111;
assign micromatrizz[79][614] = 9'b111111111;
assign micromatrizz[79][615] = 9'b111111111;
assign micromatrizz[79][616] = 9'b111111111;
assign micromatrizz[79][617] = 9'b111111111;
assign micromatrizz[79][618] = 9'b111111111;
assign micromatrizz[79][619] = 9'b111111111;
assign micromatrizz[79][620] = 9'b111111111;
assign micromatrizz[79][621] = 9'b111111111;
assign micromatrizz[79][622] = 9'b111111111;
assign micromatrizz[79][623] = 9'b111111111;
assign micromatrizz[79][624] = 9'b111111111;
assign micromatrizz[79][625] = 9'b111111111;
assign micromatrizz[79][626] = 9'b111111111;
assign micromatrizz[79][627] = 9'b111111111;
assign micromatrizz[79][628] = 9'b111111111;
assign micromatrizz[79][629] = 9'b111111111;
assign micromatrizz[79][630] = 9'b111111111;
assign micromatrizz[79][631] = 9'b111111111;
assign micromatrizz[79][632] = 9'b111111111;
assign micromatrizz[79][633] = 9'b111111111;
assign micromatrizz[79][634] = 9'b111111111;
assign micromatrizz[79][635] = 9'b111111111;
assign micromatrizz[79][636] = 9'b111111111;
assign micromatrizz[79][637] = 9'b111111111;
assign micromatrizz[79][638] = 9'b111111111;
assign micromatrizz[79][639] = 9'b111111111;
assign micromatrizz[80][0] = 9'b111111111;
assign micromatrizz[80][1] = 9'b111111111;
assign micromatrizz[80][2] = 9'b111111111;
assign micromatrizz[80][3] = 9'b111111111;
assign micromatrizz[80][4] = 9'b111111111;
assign micromatrizz[80][5] = 9'b111111111;
assign micromatrizz[80][6] = 9'b111111111;
assign micromatrizz[80][7] = 9'b111111111;
assign micromatrizz[80][8] = 9'b111111111;
assign micromatrizz[80][9] = 9'b111111111;
assign micromatrizz[80][10] = 9'b111111111;
assign micromatrizz[80][11] = 9'b111111111;
assign micromatrizz[80][12] = 9'b111111111;
assign micromatrizz[80][13] = 9'b111111111;
assign micromatrizz[80][14] = 9'b111111111;
assign micromatrizz[80][15] = 9'b111111111;
assign micromatrizz[80][16] = 9'b111111111;
assign micromatrizz[80][17] = 9'b111111111;
assign micromatrizz[80][18] = 9'b111111111;
assign micromatrizz[80][19] = 9'b111111111;
assign micromatrizz[80][20] = 9'b111111111;
assign micromatrizz[80][21] = 9'b111111111;
assign micromatrizz[80][22] = 9'b111111111;
assign micromatrizz[80][23] = 9'b111111111;
assign micromatrizz[80][24] = 9'b111111111;
assign micromatrizz[80][25] = 9'b111111111;
assign micromatrizz[80][26] = 9'b111111111;
assign micromatrizz[80][27] = 9'b111111111;
assign micromatrizz[80][28] = 9'b111111111;
assign micromatrizz[80][29] = 9'b111111111;
assign micromatrizz[80][30] = 9'b111111111;
assign micromatrizz[80][31] = 9'b111111111;
assign micromatrizz[80][32] = 9'b111111111;
assign micromatrizz[80][33] = 9'b111111111;
assign micromatrizz[80][34] = 9'b111111111;
assign micromatrizz[80][35] = 9'b111111111;
assign micromatrizz[80][36] = 9'b111111111;
assign micromatrizz[80][37] = 9'b111111111;
assign micromatrizz[80][38] = 9'b111111111;
assign micromatrizz[80][39] = 9'b111111111;
assign micromatrizz[80][40] = 9'b111111111;
assign micromatrizz[80][41] = 9'b111111111;
assign micromatrizz[80][42] = 9'b111111111;
assign micromatrizz[80][43] = 9'b111111111;
assign micromatrizz[80][44] = 9'b111111111;
assign micromatrizz[80][45] = 9'b111111111;
assign micromatrizz[80][46] = 9'b111111111;
assign micromatrizz[80][47] = 9'b111111111;
assign micromatrizz[80][48] = 9'b111111111;
assign micromatrizz[80][49] = 9'b111111111;
assign micromatrizz[80][50] = 9'b111111111;
assign micromatrizz[80][51] = 9'b111111111;
assign micromatrizz[80][52] = 9'b111111111;
assign micromatrizz[80][53] = 9'b111111111;
assign micromatrizz[80][54] = 9'b111111111;
assign micromatrizz[80][55] = 9'b111111111;
assign micromatrizz[80][56] = 9'b111111111;
assign micromatrizz[80][57] = 9'b111111111;
assign micromatrizz[80][58] = 9'b111111111;
assign micromatrizz[80][59] = 9'b111111111;
assign micromatrizz[80][60] = 9'b111111111;
assign micromatrizz[80][61] = 9'b111111111;
assign micromatrizz[80][62] = 9'b111111111;
assign micromatrizz[80][63] = 9'b111111111;
assign micromatrizz[80][64] = 9'b111111111;
assign micromatrizz[80][65] = 9'b111111111;
assign micromatrizz[80][66] = 9'b111111111;
assign micromatrizz[80][67] = 9'b111111111;
assign micromatrizz[80][68] = 9'b111111111;
assign micromatrizz[80][69] = 9'b111111111;
assign micromatrizz[80][70] = 9'b111111111;
assign micromatrizz[80][71] = 9'b111111111;
assign micromatrizz[80][72] = 9'b111111111;
assign micromatrizz[80][73] = 9'b111111111;
assign micromatrizz[80][74] = 9'b111111111;
assign micromatrizz[80][75] = 9'b111111111;
assign micromatrizz[80][76] = 9'b111111111;
assign micromatrizz[80][77] = 9'b111111111;
assign micromatrizz[80][78] = 9'b111111111;
assign micromatrizz[80][79] = 9'b111111111;
assign micromatrizz[80][80] = 9'b111111111;
assign micromatrizz[80][81] = 9'b111111111;
assign micromatrizz[80][82] = 9'b111111111;
assign micromatrizz[80][83] = 9'b111111111;
assign micromatrizz[80][84] = 9'b111111111;
assign micromatrizz[80][85] = 9'b111111111;
assign micromatrizz[80][86] = 9'b111111111;
assign micromatrizz[80][87] = 9'b111111111;
assign micromatrizz[80][88] = 9'b111111111;
assign micromatrizz[80][89] = 9'b111111111;
assign micromatrizz[80][90] = 9'b111111111;
assign micromatrizz[80][91] = 9'b111111111;
assign micromatrizz[80][92] = 9'b111111111;
assign micromatrizz[80][93] = 9'b111111111;
assign micromatrizz[80][94] = 9'b111111111;
assign micromatrizz[80][95] = 9'b111111111;
assign micromatrizz[80][96] = 9'b111111111;
assign micromatrizz[80][97] = 9'b111111111;
assign micromatrizz[80][98] = 9'b111111111;
assign micromatrizz[80][99] = 9'b111111111;
assign micromatrizz[80][100] = 9'b111111111;
assign micromatrizz[80][101] = 9'b111111111;
assign micromatrizz[80][102] = 9'b111111111;
assign micromatrizz[80][103] = 9'b111111111;
assign micromatrizz[80][104] = 9'b111111111;
assign micromatrizz[80][105] = 9'b111111111;
assign micromatrizz[80][106] = 9'b111111111;
assign micromatrizz[80][107] = 9'b111111111;
assign micromatrizz[80][108] = 9'b111111111;
assign micromatrizz[80][109] = 9'b111111111;
assign micromatrizz[80][110] = 9'b111111111;
assign micromatrizz[80][111] = 9'b111111111;
assign micromatrizz[80][112] = 9'b111111111;
assign micromatrizz[80][113] = 9'b111111111;
assign micromatrizz[80][114] = 9'b111111111;
assign micromatrizz[80][115] = 9'b111111111;
assign micromatrizz[80][116] = 9'b111111111;
assign micromatrizz[80][117] = 9'b111111111;
assign micromatrizz[80][118] = 9'b111111111;
assign micromatrizz[80][119] = 9'b111111111;
assign micromatrizz[80][120] = 9'b111111111;
assign micromatrizz[80][121] = 9'b111111111;
assign micromatrizz[80][122] = 9'b111111111;
assign micromatrizz[80][123] = 9'b111111111;
assign micromatrizz[80][124] = 9'b111111111;
assign micromatrizz[80][125] = 9'b111111111;
assign micromatrizz[80][126] = 9'b111111111;
assign micromatrizz[80][127] = 9'b111111111;
assign micromatrizz[80][128] = 9'b111111111;
assign micromatrizz[80][129] = 9'b111111111;
assign micromatrizz[80][130] = 9'b111111111;
assign micromatrizz[80][131] = 9'b111111111;
assign micromatrizz[80][132] = 9'b111111111;
assign micromatrizz[80][133] = 9'b111111111;
assign micromatrizz[80][134] = 9'b111111111;
assign micromatrizz[80][135] = 9'b111111111;
assign micromatrizz[80][136] = 9'b111111111;
assign micromatrizz[80][137] = 9'b111111111;
assign micromatrizz[80][138] = 9'b111111111;
assign micromatrizz[80][139] = 9'b111111111;
assign micromatrizz[80][140] = 9'b111111111;
assign micromatrizz[80][141] = 9'b111111111;
assign micromatrizz[80][142] = 9'b111111111;
assign micromatrizz[80][143] = 9'b111111111;
assign micromatrizz[80][144] = 9'b111111111;
assign micromatrizz[80][145] = 9'b111111111;
assign micromatrizz[80][146] = 9'b111111111;
assign micromatrizz[80][147] = 9'b111111111;
assign micromatrizz[80][148] = 9'b111111111;
assign micromatrizz[80][149] = 9'b111111111;
assign micromatrizz[80][150] = 9'b111111111;
assign micromatrizz[80][151] = 9'b111111111;
assign micromatrizz[80][152] = 9'b111111111;
assign micromatrizz[80][153] = 9'b111111111;
assign micromatrizz[80][154] = 9'b111111111;
assign micromatrizz[80][155] = 9'b111111111;
assign micromatrizz[80][156] = 9'b111111111;
assign micromatrizz[80][157] = 9'b111111111;
assign micromatrizz[80][158] = 9'b111111111;
assign micromatrizz[80][159] = 9'b111111111;
assign micromatrizz[80][160] = 9'b111111111;
assign micromatrizz[80][161] = 9'b111111111;
assign micromatrizz[80][162] = 9'b111111111;
assign micromatrizz[80][163] = 9'b111111111;
assign micromatrizz[80][164] = 9'b111111111;
assign micromatrizz[80][165] = 9'b111111111;
assign micromatrizz[80][166] = 9'b111111111;
assign micromatrizz[80][167] = 9'b111111111;
assign micromatrizz[80][168] = 9'b111111111;
assign micromatrizz[80][169] = 9'b111111111;
assign micromatrizz[80][170] = 9'b111111111;
assign micromatrizz[80][171] = 9'b111111111;
assign micromatrizz[80][172] = 9'b111111111;
assign micromatrizz[80][173] = 9'b111111111;
assign micromatrizz[80][174] = 9'b111111111;
assign micromatrizz[80][175] = 9'b111111111;
assign micromatrizz[80][176] = 9'b111111111;
assign micromatrizz[80][177] = 9'b111111111;
assign micromatrizz[80][178] = 9'b111111111;
assign micromatrizz[80][179] = 9'b111111111;
assign micromatrizz[80][180] = 9'b111111111;
assign micromatrizz[80][181] = 9'b111111111;
assign micromatrizz[80][182] = 9'b111111111;
assign micromatrizz[80][183] = 9'b111111111;
assign micromatrizz[80][184] = 9'b111111111;
assign micromatrizz[80][185] = 9'b111111111;
assign micromatrizz[80][186] = 9'b111111111;
assign micromatrizz[80][187] = 9'b111111111;
assign micromatrizz[80][188] = 9'b111111111;
assign micromatrizz[80][189] = 9'b111111111;
assign micromatrizz[80][190] = 9'b111111111;
assign micromatrizz[80][191] = 9'b111111111;
assign micromatrizz[80][192] = 9'b111111111;
assign micromatrizz[80][193] = 9'b111111111;
assign micromatrizz[80][194] = 9'b111111111;
assign micromatrizz[80][195] = 9'b111111111;
assign micromatrizz[80][196] = 9'b111111111;
assign micromatrizz[80][197] = 9'b111111111;
assign micromatrizz[80][198] = 9'b111111111;
assign micromatrizz[80][199] = 9'b111111111;
assign micromatrizz[80][200] = 9'b111111111;
assign micromatrizz[80][201] = 9'b111111111;
assign micromatrizz[80][202] = 9'b111111111;
assign micromatrizz[80][203] = 9'b111111111;
assign micromatrizz[80][204] = 9'b111111111;
assign micromatrizz[80][205] = 9'b111111111;
assign micromatrizz[80][206] = 9'b111111111;
assign micromatrizz[80][207] = 9'b111111111;
assign micromatrizz[80][208] = 9'b111111111;
assign micromatrizz[80][209] = 9'b111111111;
assign micromatrizz[80][210] = 9'b111111111;
assign micromatrizz[80][211] = 9'b111111111;
assign micromatrizz[80][212] = 9'b111111111;
assign micromatrizz[80][213] = 9'b111111111;
assign micromatrizz[80][214] = 9'b111111111;
assign micromatrizz[80][215] = 9'b111111111;
assign micromatrizz[80][216] = 9'b111111111;
assign micromatrizz[80][217] = 9'b111111111;
assign micromatrizz[80][218] = 9'b111111111;
assign micromatrizz[80][219] = 9'b111111111;
assign micromatrizz[80][220] = 9'b111111111;
assign micromatrizz[80][221] = 9'b111111111;
assign micromatrizz[80][222] = 9'b111111111;
assign micromatrizz[80][223] = 9'b111111111;
assign micromatrizz[80][224] = 9'b111111111;
assign micromatrizz[80][225] = 9'b111111111;
assign micromatrizz[80][226] = 9'b111111111;
assign micromatrizz[80][227] = 9'b111111111;
assign micromatrizz[80][228] = 9'b111111111;
assign micromatrizz[80][229] = 9'b111111111;
assign micromatrizz[80][230] = 9'b111111111;
assign micromatrizz[80][231] = 9'b111111111;
assign micromatrizz[80][232] = 9'b111111111;
assign micromatrizz[80][233] = 9'b111111111;
assign micromatrizz[80][234] = 9'b111111111;
assign micromatrizz[80][235] = 9'b111111111;
assign micromatrizz[80][236] = 9'b111111111;
assign micromatrizz[80][237] = 9'b111111111;
assign micromatrizz[80][238] = 9'b111111111;
assign micromatrizz[80][239] = 9'b111111111;
assign micromatrizz[80][240] = 9'b111111111;
assign micromatrizz[80][241] = 9'b111111111;
assign micromatrizz[80][242] = 9'b111111111;
assign micromatrizz[80][243] = 9'b111111111;
assign micromatrizz[80][244] = 9'b111111111;
assign micromatrizz[80][245] = 9'b111111111;
assign micromatrizz[80][246] = 9'b111111111;
assign micromatrizz[80][247] = 9'b111111111;
assign micromatrizz[80][248] = 9'b111111111;
assign micromatrizz[80][249] = 9'b111111111;
assign micromatrizz[80][250] = 9'b111111111;
assign micromatrizz[80][251] = 9'b111111111;
assign micromatrizz[80][252] = 9'b111111111;
assign micromatrizz[80][253] = 9'b111111111;
assign micromatrizz[80][254] = 9'b111111111;
assign micromatrizz[80][255] = 9'b111111111;
assign micromatrizz[80][256] = 9'b111111111;
assign micromatrizz[80][257] = 9'b111111111;
assign micromatrizz[80][258] = 9'b111111111;
assign micromatrizz[80][259] = 9'b111111111;
assign micromatrizz[80][260] = 9'b111111111;
assign micromatrizz[80][261] = 9'b111111111;
assign micromatrizz[80][262] = 9'b111111111;
assign micromatrizz[80][263] = 9'b111111111;
assign micromatrizz[80][264] = 9'b111111111;
assign micromatrizz[80][265] = 9'b111111111;
assign micromatrizz[80][266] = 9'b111111111;
assign micromatrizz[80][267] = 9'b111111111;
assign micromatrizz[80][268] = 9'b111111111;
assign micromatrizz[80][269] = 9'b111111111;
assign micromatrizz[80][270] = 9'b111111111;
assign micromatrizz[80][271] = 9'b111111111;
assign micromatrizz[80][272] = 9'b111111111;
assign micromatrizz[80][273] = 9'b111111111;
assign micromatrizz[80][274] = 9'b111111111;
assign micromatrizz[80][275] = 9'b111111111;
assign micromatrizz[80][276] = 9'b111111111;
assign micromatrizz[80][277] = 9'b111111111;
assign micromatrizz[80][278] = 9'b111111111;
assign micromatrizz[80][279] = 9'b111111111;
assign micromatrizz[80][280] = 9'b111111111;
assign micromatrizz[80][281] = 9'b111111111;
assign micromatrizz[80][282] = 9'b111111111;
assign micromatrizz[80][283] = 9'b111111111;
assign micromatrizz[80][284] = 9'b111111111;
assign micromatrizz[80][285] = 9'b111111111;
assign micromatrizz[80][286] = 9'b111111111;
assign micromatrizz[80][287] = 9'b111111111;
assign micromatrizz[80][288] = 9'b111111111;
assign micromatrizz[80][289] = 9'b111111111;
assign micromatrizz[80][290] = 9'b111111111;
assign micromatrizz[80][291] = 9'b111111111;
assign micromatrizz[80][292] = 9'b111111111;
assign micromatrizz[80][293] = 9'b111111111;
assign micromatrizz[80][294] = 9'b111111111;
assign micromatrizz[80][295] = 9'b111111111;
assign micromatrizz[80][296] = 9'b111111111;
assign micromatrizz[80][297] = 9'b111111111;
assign micromatrizz[80][298] = 9'b111111111;
assign micromatrizz[80][299] = 9'b111111111;
assign micromatrizz[80][300] = 9'b111111111;
assign micromatrizz[80][301] = 9'b111111111;
assign micromatrizz[80][302] = 9'b111111111;
assign micromatrizz[80][303] = 9'b111111111;
assign micromatrizz[80][304] = 9'b111111111;
assign micromatrizz[80][305] = 9'b111111111;
assign micromatrizz[80][306] = 9'b111111111;
assign micromatrizz[80][307] = 9'b111111111;
assign micromatrizz[80][308] = 9'b111111111;
assign micromatrizz[80][309] = 9'b111111111;
assign micromatrizz[80][310] = 9'b111111111;
assign micromatrizz[80][311] = 9'b111111111;
assign micromatrizz[80][312] = 9'b111111111;
assign micromatrizz[80][313] = 9'b111111111;
assign micromatrizz[80][314] = 9'b111111111;
assign micromatrizz[80][315] = 9'b111111111;
assign micromatrizz[80][316] = 9'b111111111;
assign micromatrizz[80][317] = 9'b111111111;
assign micromatrizz[80][318] = 9'b111111111;
assign micromatrizz[80][319] = 9'b111111111;
assign micromatrizz[80][320] = 9'b111111111;
assign micromatrizz[80][321] = 9'b111111111;
assign micromatrizz[80][322] = 9'b111111111;
assign micromatrizz[80][323] = 9'b111111111;
assign micromatrizz[80][324] = 9'b111111111;
assign micromatrizz[80][325] = 9'b111111111;
assign micromatrizz[80][326] = 9'b111111111;
assign micromatrizz[80][327] = 9'b111111111;
assign micromatrizz[80][328] = 9'b111111111;
assign micromatrizz[80][329] = 9'b111111111;
assign micromatrizz[80][330] = 9'b111111111;
assign micromatrizz[80][331] = 9'b111111111;
assign micromatrizz[80][332] = 9'b111111111;
assign micromatrizz[80][333] = 9'b111111111;
assign micromatrizz[80][334] = 9'b111111111;
assign micromatrizz[80][335] = 9'b111111111;
assign micromatrizz[80][336] = 9'b111111111;
assign micromatrizz[80][337] = 9'b111111111;
assign micromatrizz[80][338] = 9'b111111111;
assign micromatrizz[80][339] = 9'b111111111;
assign micromatrizz[80][340] = 9'b111111111;
assign micromatrizz[80][341] = 9'b111111111;
assign micromatrizz[80][342] = 9'b111111111;
assign micromatrizz[80][343] = 9'b111111111;
assign micromatrizz[80][344] = 9'b111111111;
assign micromatrizz[80][345] = 9'b111111111;
assign micromatrizz[80][346] = 9'b111111111;
assign micromatrizz[80][347] = 9'b111111111;
assign micromatrizz[80][348] = 9'b111111111;
assign micromatrizz[80][349] = 9'b111111111;
assign micromatrizz[80][350] = 9'b111111111;
assign micromatrizz[80][351] = 9'b111111111;
assign micromatrizz[80][352] = 9'b111111111;
assign micromatrizz[80][353] = 9'b111111111;
assign micromatrizz[80][354] = 9'b111111111;
assign micromatrizz[80][355] = 9'b111111111;
assign micromatrizz[80][356] = 9'b111111111;
assign micromatrizz[80][357] = 9'b111111111;
assign micromatrizz[80][358] = 9'b111111111;
assign micromatrizz[80][359] = 9'b111111111;
assign micromatrizz[80][360] = 9'b111111111;
assign micromatrizz[80][361] = 9'b111111111;
assign micromatrizz[80][362] = 9'b111111111;
assign micromatrizz[80][363] = 9'b111111111;
assign micromatrizz[80][364] = 9'b111111111;
assign micromatrizz[80][365] = 9'b111111111;
assign micromatrizz[80][366] = 9'b111111111;
assign micromatrizz[80][367] = 9'b111111111;
assign micromatrizz[80][368] = 9'b111111111;
assign micromatrizz[80][369] = 9'b111111111;
assign micromatrizz[80][370] = 9'b111111111;
assign micromatrizz[80][371] = 9'b111111111;
assign micromatrizz[80][372] = 9'b111111111;
assign micromatrizz[80][373] = 9'b111111111;
assign micromatrizz[80][374] = 9'b111111111;
assign micromatrizz[80][375] = 9'b111111111;
assign micromatrizz[80][376] = 9'b111111111;
assign micromatrizz[80][377] = 9'b111111111;
assign micromatrizz[80][378] = 9'b111111111;
assign micromatrizz[80][379] = 9'b111111111;
assign micromatrizz[80][380] = 9'b111111111;
assign micromatrizz[80][381] = 9'b111111111;
assign micromatrizz[80][382] = 9'b111111111;
assign micromatrizz[80][383] = 9'b111111111;
assign micromatrizz[80][384] = 9'b111111111;
assign micromatrizz[80][385] = 9'b111111111;
assign micromatrizz[80][386] = 9'b111111111;
assign micromatrizz[80][387] = 9'b111111111;
assign micromatrizz[80][388] = 9'b111111111;
assign micromatrizz[80][389] = 9'b111111111;
assign micromatrizz[80][390] = 9'b111111111;
assign micromatrizz[80][391] = 9'b111111111;
assign micromatrizz[80][392] = 9'b111111111;
assign micromatrizz[80][393] = 9'b111111111;
assign micromatrizz[80][394] = 9'b111111111;
assign micromatrizz[80][395] = 9'b111111111;
assign micromatrizz[80][396] = 9'b111111111;
assign micromatrizz[80][397] = 9'b111111111;
assign micromatrizz[80][398] = 9'b111111111;
assign micromatrizz[80][399] = 9'b111111111;
assign micromatrizz[80][400] = 9'b111111111;
assign micromatrizz[80][401] = 9'b111111111;
assign micromatrizz[80][402] = 9'b111111111;
assign micromatrizz[80][403] = 9'b111111111;
assign micromatrizz[80][404] = 9'b111111111;
assign micromatrizz[80][405] = 9'b111111111;
assign micromatrizz[80][406] = 9'b111111111;
assign micromatrizz[80][407] = 9'b111111111;
assign micromatrizz[80][408] = 9'b111111111;
assign micromatrizz[80][409] = 9'b111111111;
assign micromatrizz[80][410] = 9'b111111111;
assign micromatrizz[80][411] = 9'b111111111;
assign micromatrizz[80][412] = 9'b111111111;
assign micromatrizz[80][413] = 9'b111111111;
assign micromatrizz[80][414] = 9'b111111111;
assign micromatrizz[80][415] = 9'b111111111;
assign micromatrizz[80][416] = 9'b111111111;
assign micromatrizz[80][417] = 9'b111111111;
assign micromatrizz[80][418] = 9'b111111111;
assign micromatrizz[80][419] = 9'b111111111;
assign micromatrizz[80][420] = 9'b111111111;
assign micromatrizz[80][421] = 9'b111111111;
assign micromatrizz[80][422] = 9'b111111111;
assign micromatrizz[80][423] = 9'b111111111;
assign micromatrizz[80][424] = 9'b111111111;
assign micromatrizz[80][425] = 9'b111111111;
assign micromatrizz[80][426] = 9'b111111111;
assign micromatrizz[80][427] = 9'b111111111;
assign micromatrizz[80][428] = 9'b111111111;
assign micromatrizz[80][429] = 9'b111111111;
assign micromatrizz[80][430] = 9'b111111111;
assign micromatrizz[80][431] = 9'b111111111;
assign micromatrizz[80][432] = 9'b111111111;
assign micromatrizz[80][433] = 9'b111111111;
assign micromatrizz[80][434] = 9'b111111111;
assign micromatrizz[80][435] = 9'b111111111;
assign micromatrizz[80][436] = 9'b111111111;
assign micromatrizz[80][437] = 9'b111111111;
assign micromatrizz[80][438] = 9'b111111111;
assign micromatrizz[80][439] = 9'b111111111;
assign micromatrizz[80][440] = 9'b111111111;
assign micromatrizz[80][441] = 9'b111111111;
assign micromatrizz[80][442] = 9'b111111111;
assign micromatrizz[80][443] = 9'b111111111;
assign micromatrizz[80][444] = 9'b111111111;
assign micromatrizz[80][445] = 9'b111111111;
assign micromatrizz[80][446] = 9'b111111111;
assign micromatrizz[80][447] = 9'b111111111;
assign micromatrizz[80][448] = 9'b111111111;
assign micromatrizz[80][449] = 9'b111111111;
assign micromatrizz[80][450] = 9'b111111111;
assign micromatrizz[80][451] = 9'b111111111;
assign micromatrizz[80][452] = 9'b111111111;
assign micromatrizz[80][453] = 9'b111111111;
assign micromatrizz[80][454] = 9'b111111111;
assign micromatrizz[80][455] = 9'b111111111;
assign micromatrizz[80][456] = 9'b111111111;
assign micromatrizz[80][457] = 9'b111111111;
assign micromatrizz[80][458] = 9'b111111111;
assign micromatrizz[80][459] = 9'b111111111;
assign micromatrizz[80][460] = 9'b111111111;
assign micromatrizz[80][461] = 9'b111111111;
assign micromatrizz[80][462] = 9'b111111111;
assign micromatrizz[80][463] = 9'b111111111;
assign micromatrizz[80][464] = 9'b111111111;
assign micromatrizz[80][465] = 9'b111111111;
assign micromatrizz[80][466] = 9'b111111111;
assign micromatrizz[80][467] = 9'b111111111;
assign micromatrizz[80][468] = 9'b111111111;
assign micromatrizz[80][469] = 9'b111111111;
assign micromatrizz[80][470] = 9'b111111111;
assign micromatrizz[80][471] = 9'b111111111;
assign micromatrizz[80][472] = 9'b111111111;
assign micromatrizz[80][473] = 9'b111111111;
assign micromatrizz[80][474] = 9'b111111111;
assign micromatrizz[80][475] = 9'b111111111;
assign micromatrizz[80][476] = 9'b111111111;
assign micromatrizz[80][477] = 9'b111111111;
assign micromatrizz[80][478] = 9'b111111111;
assign micromatrizz[80][479] = 9'b111111111;
assign micromatrizz[80][480] = 9'b111111111;
assign micromatrizz[80][481] = 9'b111111111;
assign micromatrizz[80][482] = 9'b111111111;
assign micromatrizz[80][483] = 9'b111111111;
assign micromatrizz[80][484] = 9'b111111111;
assign micromatrizz[80][485] = 9'b111111111;
assign micromatrizz[80][486] = 9'b111111111;
assign micromatrizz[80][487] = 9'b111111111;
assign micromatrizz[80][488] = 9'b111111111;
assign micromatrizz[80][489] = 9'b111111111;
assign micromatrizz[80][490] = 9'b111111111;
assign micromatrizz[80][491] = 9'b111111111;
assign micromatrizz[80][492] = 9'b111111111;
assign micromatrizz[80][493] = 9'b111111111;
assign micromatrizz[80][494] = 9'b111111111;
assign micromatrizz[80][495] = 9'b111111111;
assign micromatrizz[80][496] = 9'b111111111;
assign micromatrizz[80][497] = 9'b111111111;
assign micromatrizz[80][498] = 9'b111111111;
assign micromatrizz[80][499] = 9'b111111111;
assign micromatrizz[80][500] = 9'b111111111;
assign micromatrizz[80][501] = 9'b111111111;
assign micromatrizz[80][502] = 9'b111111111;
assign micromatrizz[80][503] = 9'b111111111;
assign micromatrizz[80][504] = 9'b111111111;
assign micromatrizz[80][505] = 9'b111111111;
assign micromatrizz[80][506] = 9'b111111111;
assign micromatrizz[80][507] = 9'b111111111;
assign micromatrizz[80][508] = 9'b111111111;
assign micromatrizz[80][509] = 9'b111111111;
assign micromatrizz[80][510] = 9'b111111111;
assign micromatrizz[80][511] = 9'b111111111;
assign micromatrizz[80][512] = 9'b111111111;
assign micromatrizz[80][513] = 9'b111111111;
assign micromatrizz[80][514] = 9'b111111111;
assign micromatrizz[80][515] = 9'b111111111;
assign micromatrizz[80][516] = 9'b111111111;
assign micromatrizz[80][517] = 9'b111111111;
assign micromatrizz[80][518] = 9'b111111111;
assign micromatrizz[80][519] = 9'b111111111;
assign micromatrizz[80][520] = 9'b111111111;
assign micromatrizz[80][521] = 9'b111111111;
assign micromatrizz[80][522] = 9'b111111111;
assign micromatrizz[80][523] = 9'b111111111;
assign micromatrizz[80][524] = 9'b111111111;
assign micromatrizz[80][525] = 9'b111111111;
assign micromatrizz[80][526] = 9'b111111111;
assign micromatrizz[80][527] = 9'b111111111;
assign micromatrizz[80][528] = 9'b111111111;
assign micromatrizz[80][529] = 9'b111111111;
assign micromatrizz[80][530] = 9'b111111111;
assign micromatrizz[80][531] = 9'b111111111;
assign micromatrizz[80][532] = 9'b111111111;
assign micromatrizz[80][533] = 9'b111111111;
assign micromatrizz[80][534] = 9'b111111111;
assign micromatrizz[80][535] = 9'b111111111;
assign micromatrizz[80][536] = 9'b111111111;
assign micromatrizz[80][537] = 9'b111111111;
assign micromatrizz[80][538] = 9'b111111111;
assign micromatrizz[80][539] = 9'b111111111;
assign micromatrizz[80][540] = 9'b111111111;
assign micromatrizz[80][541] = 9'b111111111;
assign micromatrizz[80][542] = 9'b111111111;
assign micromatrizz[80][543] = 9'b111111111;
assign micromatrizz[80][544] = 9'b111111111;
assign micromatrizz[80][545] = 9'b111111111;
assign micromatrizz[80][546] = 9'b111111111;
assign micromatrizz[80][547] = 9'b111111111;
assign micromatrizz[80][548] = 9'b111111111;
assign micromatrizz[80][549] = 9'b111111111;
assign micromatrizz[80][550] = 9'b111111111;
assign micromatrizz[80][551] = 9'b111111111;
assign micromatrizz[80][552] = 9'b111111111;
assign micromatrizz[80][553] = 9'b111111111;
assign micromatrizz[80][554] = 9'b111111111;
assign micromatrizz[80][555] = 9'b111111111;
assign micromatrizz[80][556] = 9'b111111111;
assign micromatrizz[80][557] = 9'b111111111;
assign micromatrizz[80][558] = 9'b111111111;
assign micromatrizz[80][559] = 9'b111111111;
assign micromatrizz[80][560] = 9'b111111111;
assign micromatrizz[80][561] = 9'b111111111;
assign micromatrizz[80][562] = 9'b111111111;
assign micromatrizz[80][563] = 9'b111111111;
assign micromatrizz[80][564] = 9'b111111111;
assign micromatrizz[80][565] = 9'b111111111;
assign micromatrizz[80][566] = 9'b111111111;
assign micromatrizz[80][567] = 9'b111111111;
assign micromatrizz[80][568] = 9'b111111111;
assign micromatrizz[80][569] = 9'b111111111;
assign micromatrizz[80][570] = 9'b111111111;
assign micromatrizz[80][571] = 9'b111111111;
assign micromatrizz[80][572] = 9'b111111111;
assign micromatrizz[80][573] = 9'b111111111;
assign micromatrizz[80][574] = 9'b111111111;
assign micromatrizz[80][575] = 9'b111111111;
assign micromatrizz[80][576] = 9'b111111111;
assign micromatrizz[80][577] = 9'b111111111;
assign micromatrizz[80][578] = 9'b111111111;
assign micromatrizz[80][579] = 9'b111111111;
assign micromatrizz[80][580] = 9'b111111111;
assign micromatrizz[80][581] = 9'b111111111;
assign micromatrizz[80][582] = 9'b111111111;
assign micromatrizz[80][583] = 9'b111111111;
assign micromatrizz[80][584] = 9'b111111111;
assign micromatrizz[80][585] = 9'b111111111;
assign micromatrizz[80][586] = 9'b111111111;
assign micromatrizz[80][587] = 9'b111111111;
assign micromatrizz[80][588] = 9'b111111111;
assign micromatrizz[80][589] = 9'b111111111;
assign micromatrizz[80][590] = 9'b111111111;
assign micromatrizz[80][591] = 9'b111111111;
assign micromatrizz[80][592] = 9'b111111111;
assign micromatrizz[80][593] = 9'b111111111;
assign micromatrizz[80][594] = 9'b111111111;
assign micromatrizz[80][595] = 9'b111111111;
assign micromatrizz[80][596] = 9'b111111111;
assign micromatrizz[80][597] = 9'b111111111;
assign micromatrizz[80][598] = 9'b111111111;
assign micromatrizz[80][599] = 9'b111111111;
assign micromatrizz[80][600] = 9'b111111111;
assign micromatrizz[80][601] = 9'b111111111;
assign micromatrizz[80][602] = 9'b111111111;
assign micromatrizz[80][603] = 9'b111111111;
assign micromatrizz[80][604] = 9'b111111111;
assign micromatrizz[80][605] = 9'b111111111;
assign micromatrizz[80][606] = 9'b111111111;
assign micromatrizz[80][607] = 9'b111111111;
assign micromatrizz[80][608] = 9'b111111111;
assign micromatrizz[80][609] = 9'b111111111;
assign micromatrizz[80][610] = 9'b111111111;
assign micromatrizz[80][611] = 9'b111111111;
assign micromatrizz[80][612] = 9'b111111111;
assign micromatrizz[80][613] = 9'b111111111;
assign micromatrizz[80][614] = 9'b111111111;
assign micromatrizz[80][615] = 9'b111111111;
assign micromatrizz[80][616] = 9'b111111111;
assign micromatrizz[80][617] = 9'b111111111;
assign micromatrizz[80][618] = 9'b111111111;
assign micromatrizz[80][619] = 9'b111111111;
assign micromatrizz[80][620] = 9'b111111111;
assign micromatrizz[80][621] = 9'b111111111;
assign micromatrizz[80][622] = 9'b111111111;
assign micromatrizz[80][623] = 9'b111111111;
assign micromatrizz[80][624] = 9'b111111111;
assign micromatrizz[80][625] = 9'b111111111;
assign micromatrizz[80][626] = 9'b111111111;
assign micromatrizz[80][627] = 9'b111111111;
assign micromatrizz[80][628] = 9'b111111111;
assign micromatrizz[80][629] = 9'b111111111;
assign micromatrizz[80][630] = 9'b111111111;
assign micromatrizz[80][631] = 9'b111111111;
assign micromatrizz[80][632] = 9'b111111111;
assign micromatrizz[80][633] = 9'b111111111;
assign micromatrizz[80][634] = 9'b111111111;
assign micromatrizz[80][635] = 9'b111111111;
assign micromatrizz[80][636] = 9'b111111111;
assign micromatrizz[80][637] = 9'b111111111;
assign micromatrizz[80][638] = 9'b111111111;
assign micromatrizz[80][639] = 9'b111111111;
assign micromatrizz[81][0] = 9'b111111111;
assign micromatrizz[81][1] = 9'b111111111;
assign micromatrizz[81][2] = 9'b111111111;
assign micromatrizz[81][3] = 9'b111111111;
assign micromatrizz[81][4] = 9'b111111111;
assign micromatrizz[81][5] = 9'b111111111;
assign micromatrizz[81][6] = 9'b111111111;
assign micromatrizz[81][7] = 9'b111111111;
assign micromatrizz[81][8] = 9'b111111111;
assign micromatrizz[81][9] = 9'b111111111;
assign micromatrizz[81][10] = 9'b111111111;
assign micromatrizz[81][11] = 9'b111111111;
assign micromatrizz[81][12] = 9'b111111111;
assign micromatrizz[81][13] = 9'b111111111;
assign micromatrizz[81][14] = 9'b111111111;
assign micromatrizz[81][15] = 9'b111111111;
assign micromatrizz[81][16] = 9'b111111111;
assign micromatrizz[81][17] = 9'b111111111;
assign micromatrizz[81][18] = 9'b111111111;
assign micromatrizz[81][19] = 9'b111111111;
assign micromatrizz[81][20] = 9'b111111111;
assign micromatrizz[81][21] = 9'b111111111;
assign micromatrizz[81][22] = 9'b111111111;
assign micromatrizz[81][23] = 9'b111111111;
assign micromatrizz[81][24] = 9'b111111111;
assign micromatrizz[81][25] = 9'b111111111;
assign micromatrizz[81][26] = 9'b111111111;
assign micromatrizz[81][27] = 9'b111111111;
assign micromatrizz[81][28] = 9'b111111111;
assign micromatrizz[81][29] = 9'b111111111;
assign micromatrizz[81][30] = 9'b111111111;
assign micromatrizz[81][31] = 9'b111111111;
assign micromatrizz[81][32] = 9'b111111111;
assign micromatrizz[81][33] = 9'b111111111;
assign micromatrizz[81][34] = 9'b111111111;
assign micromatrizz[81][35] = 9'b111111111;
assign micromatrizz[81][36] = 9'b111111111;
assign micromatrizz[81][37] = 9'b111111111;
assign micromatrizz[81][38] = 9'b111111111;
assign micromatrizz[81][39] = 9'b111111111;
assign micromatrizz[81][40] = 9'b111111111;
assign micromatrizz[81][41] = 9'b111111111;
assign micromatrizz[81][42] = 9'b111111111;
assign micromatrizz[81][43] = 9'b111111111;
assign micromatrizz[81][44] = 9'b111111111;
assign micromatrizz[81][45] = 9'b111111111;
assign micromatrizz[81][46] = 9'b111111111;
assign micromatrizz[81][47] = 9'b111111111;
assign micromatrizz[81][48] = 9'b111111111;
assign micromatrizz[81][49] = 9'b111111111;
assign micromatrizz[81][50] = 9'b111111111;
assign micromatrizz[81][51] = 9'b111111111;
assign micromatrizz[81][52] = 9'b111111111;
assign micromatrizz[81][53] = 9'b111111111;
assign micromatrizz[81][54] = 9'b111111111;
assign micromatrizz[81][55] = 9'b111111111;
assign micromatrizz[81][56] = 9'b111111111;
assign micromatrizz[81][57] = 9'b111111111;
assign micromatrizz[81][58] = 9'b111111111;
assign micromatrizz[81][59] = 9'b111111111;
assign micromatrizz[81][60] = 9'b111111111;
assign micromatrizz[81][61] = 9'b111111111;
assign micromatrizz[81][62] = 9'b111111111;
assign micromatrizz[81][63] = 9'b111111111;
assign micromatrizz[81][64] = 9'b111111111;
assign micromatrizz[81][65] = 9'b111111111;
assign micromatrizz[81][66] = 9'b111111111;
assign micromatrizz[81][67] = 9'b111111111;
assign micromatrizz[81][68] = 9'b111111111;
assign micromatrizz[81][69] = 9'b111111111;
assign micromatrizz[81][70] = 9'b111111111;
assign micromatrizz[81][71] = 9'b111111111;
assign micromatrizz[81][72] = 9'b111111111;
assign micromatrizz[81][73] = 9'b111111111;
assign micromatrizz[81][74] = 9'b111111111;
assign micromatrizz[81][75] = 9'b111111111;
assign micromatrizz[81][76] = 9'b111111111;
assign micromatrizz[81][77] = 9'b111111111;
assign micromatrizz[81][78] = 9'b111111111;
assign micromatrizz[81][79] = 9'b111111111;
assign micromatrizz[81][80] = 9'b111111111;
assign micromatrizz[81][81] = 9'b111111111;
assign micromatrizz[81][82] = 9'b111111111;
assign micromatrizz[81][83] = 9'b111111111;
assign micromatrizz[81][84] = 9'b111111111;
assign micromatrizz[81][85] = 9'b111111111;
assign micromatrizz[81][86] = 9'b111111111;
assign micromatrizz[81][87] = 9'b111111111;
assign micromatrizz[81][88] = 9'b111111111;
assign micromatrizz[81][89] = 9'b111111111;
assign micromatrizz[81][90] = 9'b111111111;
assign micromatrizz[81][91] = 9'b111111111;
assign micromatrizz[81][92] = 9'b111111111;
assign micromatrizz[81][93] = 9'b111111111;
assign micromatrizz[81][94] = 9'b111111111;
assign micromatrizz[81][95] = 9'b111111111;
assign micromatrizz[81][96] = 9'b111111111;
assign micromatrizz[81][97] = 9'b111111111;
assign micromatrizz[81][98] = 9'b111111111;
assign micromatrizz[81][99] = 9'b111111111;
assign micromatrizz[81][100] = 9'b111111111;
assign micromatrizz[81][101] = 9'b111111111;
assign micromatrizz[81][102] = 9'b111111111;
assign micromatrizz[81][103] = 9'b111111111;
assign micromatrizz[81][104] = 9'b111111111;
assign micromatrizz[81][105] = 9'b111111111;
assign micromatrizz[81][106] = 9'b111111111;
assign micromatrizz[81][107] = 9'b111111111;
assign micromatrizz[81][108] = 9'b111111111;
assign micromatrizz[81][109] = 9'b111111111;
assign micromatrizz[81][110] = 9'b111111111;
assign micromatrizz[81][111] = 9'b111111111;
assign micromatrizz[81][112] = 9'b111111111;
assign micromatrizz[81][113] = 9'b111111111;
assign micromatrizz[81][114] = 9'b111111111;
assign micromatrizz[81][115] = 9'b111111111;
assign micromatrizz[81][116] = 9'b111111111;
assign micromatrizz[81][117] = 9'b111111111;
assign micromatrizz[81][118] = 9'b111111111;
assign micromatrizz[81][119] = 9'b111111111;
assign micromatrizz[81][120] = 9'b111111111;
assign micromatrizz[81][121] = 9'b111111111;
assign micromatrizz[81][122] = 9'b111111111;
assign micromatrizz[81][123] = 9'b111111111;
assign micromatrizz[81][124] = 9'b111111111;
assign micromatrizz[81][125] = 9'b111111111;
assign micromatrizz[81][126] = 9'b111111111;
assign micromatrizz[81][127] = 9'b111111111;
assign micromatrizz[81][128] = 9'b111111111;
assign micromatrizz[81][129] = 9'b111111111;
assign micromatrizz[81][130] = 9'b111111111;
assign micromatrizz[81][131] = 9'b111111111;
assign micromatrizz[81][132] = 9'b111111111;
assign micromatrizz[81][133] = 9'b111111111;
assign micromatrizz[81][134] = 9'b111111111;
assign micromatrizz[81][135] = 9'b111111111;
assign micromatrizz[81][136] = 9'b111111111;
assign micromatrizz[81][137] = 9'b111111111;
assign micromatrizz[81][138] = 9'b111111111;
assign micromatrizz[81][139] = 9'b111111111;
assign micromatrizz[81][140] = 9'b111111111;
assign micromatrizz[81][141] = 9'b111111111;
assign micromatrizz[81][142] = 9'b111111111;
assign micromatrizz[81][143] = 9'b111111111;
assign micromatrizz[81][144] = 9'b111111111;
assign micromatrizz[81][145] = 9'b111111111;
assign micromatrizz[81][146] = 9'b111111111;
assign micromatrizz[81][147] = 9'b111111111;
assign micromatrizz[81][148] = 9'b111111111;
assign micromatrizz[81][149] = 9'b111111111;
assign micromatrizz[81][150] = 9'b111111111;
assign micromatrizz[81][151] = 9'b111111111;
assign micromatrizz[81][152] = 9'b111111111;
assign micromatrizz[81][153] = 9'b111111111;
assign micromatrizz[81][154] = 9'b111111111;
assign micromatrizz[81][155] = 9'b111111111;
assign micromatrizz[81][156] = 9'b111111111;
assign micromatrizz[81][157] = 9'b111111111;
assign micromatrizz[81][158] = 9'b111111111;
assign micromatrizz[81][159] = 9'b111111111;
assign micromatrizz[81][160] = 9'b111111111;
assign micromatrizz[81][161] = 9'b111111111;
assign micromatrizz[81][162] = 9'b111111111;
assign micromatrizz[81][163] = 9'b111111111;
assign micromatrizz[81][164] = 9'b111111111;
assign micromatrizz[81][165] = 9'b111111111;
assign micromatrizz[81][166] = 9'b111111111;
assign micromatrizz[81][167] = 9'b111111111;
assign micromatrizz[81][168] = 9'b111111111;
assign micromatrizz[81][169] = 9'b111111111;
assign micromatrizz[81][170] = 9'b111111111;
assign micromatrizz[81][171] = 9'b111111111;
assign micromatrizz[81][172] = 9'b111111111;
assign micromatrizz[81][173] = 9'b111111111;
assign micromatrizz[81][174] = 9'b111111111;
assign micromatrizz[81][175] = 9'b111111111;
assign micromatrizz[81][176] = 9'b111111111;
assign micromatrizz[81][177] = 9'b111111111;
assign micromatrizz[81][178] = 9'b111111111;
assign micromatrizz[81][179] = 9'b111111111;
assign micromatrizz[81][180] = 9'b111111111;
assign micromatrizz[81][181] = 9'b111111111;
assign micromatrizz[81][182] = 9'b111111111;
assign micromatrizz[81][183] = 9'b111111111;
assign micromatrizz[81][184] = 9'b111111111;
assign micromatrizz[81][185] = 9'b111111111;
assign micromatrizz[81][186] = 9'b111111111;
assign micromatrizz[81][187] = 9'b111111111;
assign micromatrizz[81][188] = 9'b111111111;
assign micromatrizz[81][189] = 9'b111111111;
assign micromatrizz[81][190] = 9'b111111111;
assign micromatrizz[81][191] = 9'b111111111;
assign micromatrizz[81][192] = 9'b111111111;
assign micromatrizz[81][193] = 9'b111111111;
assign micromatrizz[81][194] = 9'b111111111;
assign micromatrizz[81][195] = 9'b111111111;
assign micromatrizz[81][196] = 9'b111111111;
assign micromatrizz[81][197] = 9'b111111111;
assign micromatrizz[81][198] = 9'b111111111;
assign micromatrizz[81][199] = 9'b111111111;
assign micromatrizz[81][200] = 9'b111111111;
assign micromatrizz[81][201] = 9'b111111111;
assign micromatrizz[81][202] = 9'b111111111;
assign micromatrizz[81][203] = 9'b111111111;
assign micromatrizz[81][204] = 9'b111111111;
assign micromatrizz[81][205] = 9'b111111111;
assign micromatrizz[81][206] = 9'b111111111;
assign micromatrizz[81][207] = 9'b111111111;
assign micromatrizz[81][208] = 9'b111111111;
assign micromatrizz[81][209] = 9'b111111111;
assign micromatrizz[81][210] = 9'b111111111;
assign micromatrizz[81][211] = 9'b111111111;
assign micromatrizz[81][212] = 9'b111111111;
assign micromatrizz[81][213] = 9'b111111111;
assign micromatrizz[81][214] = 9'b111111111;
assign micromatrizz[81][215] = 9'b111111111;
assign micromatrizz[81][216] = 9'b111111111;
assign micromatrizz[81][217] = 9'b111111111;
assign micromatrizz[81][218] = 9'b111111111;
assign micromatrizz[81][219] = 9'b111111111;
assign micromatrizz[81][220] = 9'b111111111;
assign micromatrizz[81][221] = 9'b111111111;
assign micromatrizz[81][222] = 9'b111111111;
assign micromatrizz[81][223] = 9'b111111111;
assign micromatrizz[81][224] = 9'b111111111;
assign micromatrizz[81][225] = 9'b111111111;
assign micromatrizz[81][226] = 9'b111111111;
assign micromatrizz[81][227] = 9'b111111111;
assign micromatrizz[81][228] = 9'b111111111;
assign micromatrizz[81][229] = 9'b111111111;
assign micromatrizz[81][230] = 9'b111111111;
assign micromatrizz[81][231] = 9'b111111111;
assign micromatrizz[81][232] = 9'b111111111;
assign micromatrizz[81][233] = 9'b111111111;
assign micromatrizz[81][234] = 9'b111111111;
assign micromatrizz[81][235] = 9'b111111111;
assign micromatrizz[81][236] = 9'b111111111;
assign micromatrizz[81][237] = 9'b111111111;
assign micromatrizz[81][238] = 9'b111111111;
assign micromatrizz[81][239] = 9'b111111111;
assign micromatrizz[81][240] = 9'b111111111;
assign micromatrizz[81][241] = 9'b111111111;
assign micromatrizz[81][242] = 9'b111111111;
assign micromatrizz[81][243] = 9'b111111111;
assign micromatrizz[81][244] = 9'b111111111;
assign micromatrizz[81][245] = 9'b111111111;
assign micromatrizz[81][246] = 9'b111111111;
assign micromatrizz[81][247] = 9'b111111111;
assign micromatrizz[81][248] = 9'b111111111;
assign micromatrizz[81][249] = 9'b111111111;
assign micromatrizz[81][250] = 9'b111111111;
assign micromatrizz[81][251] = 9'b111111111;
assign micromatrizz[81][252] = 9'b111111111;
assign micromatrizz[81][253] = 9'b111111111;
assign micromatrizz[81][254] = 9'b111111111;
assign micromatrizz[81][255] = 9'b111111111;
assign micromatrizz[81][256] = 9'b111111111;
assign micromatrizz[81][257] = 9'b111111111;
assign micromatrizz[81][258] = 9'b111111111;
assign micromatrizz[81][259] = 9'b111111111;
assign micromatrizz[81][260] = 9'b111111111;
assign micromatrizz[81][261] = 9'b111111111;
assign micromatrizz[81][262] = 9'b111111111;
assign micromatrizz[81][263] = 9'b111111111;
assign micromatrizz[81][264] = 9'b111111111;
assign micromatrizz[81][265] = 9'b111111111;
assign micromatrizz[81][266] = 9'b111111111;
assign micromatrizz[81][267] = 9'b111111111;
assign micromatrizz[81][268] = 9'b111111111;
assign micromatrizz[81][269] = 9'b111111111;
assign micromatrizz[81][270] = 9'b111111111;
assign micromatrizz[81][271] = 9'b111111111;
assign micromatrizz[81][272] = 9'b111111111;
assign micromatrizz[81][273] = 9'b111111111;
assign micromatrizz[81][274] = 9'b111111111;
assign micromatrizz[81][275] = 9'b111111111;
assign micromatrizz[81][276] = 9'b111111111;
assign micromatrizz[81][277] = 9'b111111111;
assign micromatrizz[81][278] = 9'b111111111;
assign micromatrizz[81][279] = 9'b111111111;
assign micromatrizz[81][280] = 9'b111111111;
assign micromatrizz[81][281] = 9'b111111111;
assign micromatrizz[81][282] = 9'b111111111;
assign micromatrizz[81][283] = 9'b111111111;
assign micromatrizz[81][284] = 9'b111111111;
assign micromatrizz[81][285] = 9'b111111111;
assign micromatrizz[81][286] = 9'b111111111;
assign micromatrizz[81][287] = 9'b111111111;
assign micromatrizz[81][288] = 9'b111111111;
assign micromatrizz[81][289] = 9'b111111111;
assign micromatrizz[81][290] = 9'b111111111;
assign micromatrizz[81][291] = 9'b111111111;
assign micromatrizz[81][292] = 9'b111111111;
assign micromatrizz[81][293] = 9'b111111111;
assign micromatrizz[81][294] = 9'b111111111;
assign micromatrizz[81][295] = 9'b111111111;
assign micromatrizz[81][296] = 9'b111111111;
assign micromatrizz[81][297] = 9'b111111111;
assign micromatrizz[81][298] = 9'b111111111;
assign micromatrizz[81][299] = 9'b111111111;
assign micromatrizz[81][300] = 9'b111111111;
assign micromatrizz[81][301] = 9'b111111111;
assign micromatrizz[81][302] = 9'b111111111;
assign micromatrizz[81][303] = 9'b111111111;
assign micromatrizz[81][304] = 9'b111111111;
assign micromatrizz[81][305] = 9'b111111111;
assign micromatrizz[81][306] = 9'b111111111;
assign micromatrizz[81][307] = 9'b111111111;
assign micromatrizz[81][308] = 9'b111111111;
assign micromatrizz[81][309] = 9'b111111111;
assign micromatrizz[81][310] = 9'b111111111;
assign micromatrizz[81][311] = 9'b111111111;
assign micromatrizz[81][312] = 9'b111111111;
assign micromatrizz[81][313] = 9'b111111111;
assign micromatrizz[81][314] = 9'b111111111;
assign micromatrizz[81][315] = 9'b111111111;
assign micromatrizz[81][316] = 9'b111111111;
assign micromatrizz[81][317] = 9'b111111111;
assign micromatrizz[81][318] = 9'b111111111;
assign micromatrizz[81][319] = 9'b111111111;
assign micromatrizz[81][320] = 9'b111111111;
assign micromatrizz[81][321] = 9'b111111111;
assign micromatrizz[81][322] = 9'b111111111;
assign micromatrizz[81][323] = 9'b111111111;
assign micromatrizz[81][324] = 9'b111111111;
assign micromatrizz[81][325] = 9'b111111111;
assign micromatrizz[81][326] = 9'b111111111;
assign micromatrizz[81][327] = 9'b111111111;
assign micromatrizz[81][328] = 9'b111111111;
assign micromatrizz[81][329] = 9'b111111111;
assign micromatrizz[81][330] = 9'b111111111;
assign micromatrizz[81][331] = 9'b111111111;
assign micromatrizz[81][332] = 9'b111111111;
assign micromatrizz[81][333] = 9'b111111111;
assign micromatrizz[81][334] = 9'b111111111;
assign micromatrizz[81][335] = 9'b111111111;
assign micromatrizz[81][336] = 9'b111111111;
assign micromatrizz[81][337] = 9'b111111111;
assign micromatrizz[81][338] = 9'b111111111;
assign micromatrizz[81][339] = 9'b111111111;
assign micromatrizz[81][340] = 9'b111111111;
assign micromatrizz[81][341] = 9'b111111111;
assign micromatrizz[81][342] = 9'b111111111;
assign micromatrizz[81][343] = 9'b111111111;
assign micromatrizz[81][344] = 9'b111111111;
assign micromatrizz[81][345] = 9'b111111111;
assign micromatrizz[81][346] = 9'b111111111;
assign micromatrizz[81][347] = 9'b111111111;
assign micromatrizz[81][348] = 9'b111111111;
assign micromatrizz[81][349] = 9'b111111111;
assign micromatrizz[81][350] = 9'b111111111;
assign micromatrizz[81][351] = 9'b111111111;
assign micromatrizz[81][352] = 9'b111111111;
assign micromatrizz[81][353] = 9'b111111111;
assign micromatrizz[81][354] = 9'b111111111;
assign micromatrizz[81][355] = 9'b111111111;
assign micromatrizz[81][356] = 9'b111111111;
assign micromatrizz[81][357] = 9'b111111111;
assign micromatrizz[81][358] = 9'b111111111;
assign micromatrizz[81][359] = 9'b111111111;
assign micromatrizz[81][360] = 9'b111111111;
assign micromatrizz[81][361] = 9'b111111111;
assign micromatrizz[81][362] = 9'b111111111;
assign micromatrizz[81][363] = 9'b111111111;
assign micromatrizz[81][364] = 9'b111111111;
assign micromatrizz[81][365] = 9'b111111111;
assign micromatrizz[81][366] = 9'b111111111;
assign micromatrizz[81][367] = 9'b111111111;
assign micromatrizz[81][368] = 9'b111111111;
assign micromatrizz[81][369] = 9'b111111111;
assign micromatrizz[81][370] = 9'b111111111;
assign micromatrizz[81][371] = 9'b111111111;
assign micromatrizz[81][372] = 9'b111111111;
assign micromatrizz[81][373] = 9'b111111111;
assign micromatrizz[81][374] = 9'b111111111;
assign micromatrizz[81][375] = 9'b111111111;
assign micromatrizz[81][376] = 9'b111111111;
assign micromatrizz[81][377] = 9'b111111111;
assign micromatrizz[81][378] = 9'b111111111;
assign micromatrizz[81][379] = 9'b111111111;
assign micromatrizz[81][380] = 9'b111111111;
assign micromatrizz[81][381] = 9'b111111111;
assign micromatrizz[81][382] = 9'b111111111;
assign micromatrizz[81][383] = 9'b111111111;
assign micromatrizz[81][384] = 9'b111111111;
assign micromatrizz[81][385] = 9'b111111111;
assign micromatrizz[81][386] = 9'b111111111;
assign micromatrizz[81][387] = 9'b111111111;
assign micromatrizz[81][388] = 9'b111111111;
assign micromatrizz[81][389] = 9'b111111111;
assign micromatrizz[81][390] = 9'b111111111;
assign micromatrizz[81][391] = 9'b111111111;
assign micromatrizz[81][392] = 9'b111111111;
assign micromatrizz[81][393] = 9'b111111111;
assign micromatrizz[81][394] = 9'b111111111;
assign micromatrizz[81][395] = 9'b111111111;
assign micromatrizz[81][396] = 9'b111111111;
assign micromatrizz[81][397] = 9'b111111111;
assign micromatrizz[81][398] = 9'b111111111;
assign micromatrizz[81][399] = 9'b111111111;
assign micromatrizz[81][400] = 9'b111111111;
assign micromatrizz[81][401] = 9'b111111111;
assign micromatrizz[81][402] = 9'b111111111;
assign micromatrizz[81][403] = 9'b111111111;
assign micromatrizz[81][404] = 9'b111111111;
assign micromatrizz[81][405] = 9'b111111111;
assign micromatrizz[81][406] = 9'b111111111;
assign micromatrizz[81][407] = 9'b111111111;
assign micromatrizz[81][408] = 9'b111111111;
assign micromatrizz[81][409] = 9'b111111111;
assign micromatrizz[81][410] = 9'b111111111;
assign micromatrizz[81][411] = 9'b111111111;
assign micromatrizz[81][412] = 9'b111111111;
assign micromatrizz[81][413] = 9'b111111111;
assign micromatrizz[81][414] = 9'b111111111;
assign micromatrizz[81][415] = 9'b111111111;
assign micromatrizz[81][416] = 9'b111111111;
assign micromatrizz[81][417] = 9'b111111111;
assign micromatrizz[81][418] = 9'b111111111;
assign micromatrizz[81][419] = 9'b111111111;
assign micromatrizz[81][420] = 9'b111111111;
assign micromatrizz[81][421] = 9'b111111111;
assign micromatrizz[81][422] = 9'b111111111;
assign micromatrizz[81][423] = 9'b111111111;
assign micromatrizz[81][424] = 9'b111111111;
assign micromatrizz[81][425] = 9'b111111111;
assign micromatrizz[81][426] = 9'b111111111;
assign micromatrizz[81][427] = 9'b111111111;
assign micromatrizz[81][428] = 9'b111111111;
assign micromatrizz[81][429] = 9'b111111111;
assign micromatrizz[81][430] = 9'b111111111;
assign micromatrizz[81][431] = 9'b111111111;
assign micromatrizz[81][432] = 9'b111111111;
assign micromatrizz[81][433] = 9'b111111111;
assign micromatrizz[81][434] = 9'b111111111;
assign micromatrizz[81][435] = 9'b111111111;
assign micromatrizz[81][436] = 9'b111111111;
assign micromatrizz[81][437] = 9'b111111111;
assign micromatrizz[81][438] = 9'b111111111;
assign micromatrizz[81][439] = 9'b111111111;
assign micromatrizz[81][440] = 9'b111111111;
assign micromatrizz[81][441] = 9'b111111111;
assign micromatrizz[81][442] = 9'b111111111;
assign micromatrizz[81][443] = 9'b111111111;
assign micromatrizz[81][444] = 9'b111111111;
assign micromatrizz[81][445] = 9'b111111111;
assign micromatrizz[81][446] = 9'b111111111;
assign micromatrizz[81][447] = 9'b111111111;
assign micromatrizz[81][448] = 9'b111111111;
assign micromatrizz[81][449] = 9'b111111111;
assign micromatrizz[81][450] = 9'b111111111;
assign micromatrizz[81][451] = 9'b111111111;
assign micromatrizz[81][452] = 9'b111111111;
assign micromatrizz[81][453] = 9'b111111111;
assign micromatrizz[81][454] = 9'b111111111;
assign micromatrizz[81][455] = 9'b111111111;
assign micromatrizz[81][456] = 9'b111111111;
assign micromatrizz[81][457] = 9'b111111111;
assign micromatrizz[81][458] = 9'b111111111;
assign micromatrizz[81][459] = 9'b111111111;
assign micromatrizz[81][460] = 9'b111111111;
assign micromatrizz[81][461] = 9'b111111111;
assign micromatrizz[81][462] = 9'b111111111;
assign micromatrizz[81][463] = 9'b111111111;
assign micromatrizz[81][464] = 9'b111111111;
assign micromatrizz[81][465] = 9'b111111111;
assign micromatrizz[81][466] = 9'b111111111;
assign micromatrizz[81][467] = 9'b111111111;
assign micromatrizz[81][468] = 9'b111111111;
assign micromatrizz[81][469] = 9'b111111111;
assign micromatrizz[81][470] = 9'b111111111;
assign micromatrizz[81][471] = 9'b111111111;
assign micromatrizz[81][472] = 9'b111111111;
assign micromatrizz[81][473] = 9'b111111111;
assign micromatrizz[81][474] = 9'b111111111;
assign micromatrizz[81][475] = 9'b111111111;
assign micromatrizz[81][476] = 9'b111111111;
assign micromatrizz[81][477] = 9'b111111111;
assign micromatrizz[81][478] = 9'b111111111;
assign micromatrizz[81][479] = 9'b111111111;
assign micromatrizz[81][480] = 9'b111111111;
assign micromatrizz[81][481] = 9'b111111111;
assign micromatrizz[81][482] = 9'b111111111;
assign micromatrizz[81][483] = 9'b111111111;
assign micromatrizz[81][484] = 9'b111111111;
assign micromatrizz[81][485] = 9'b111111111;
assign micromatrizz[81][486] = 9'b111111111;
assign micromatrizz[81][487] = 9'b111111111;
assign micromatrizz[81][488] = 9'b111111111;
assign micromatrizz[81][489] = 9'b111111111;
assign micromatrizz[81][490] = 9'b111111111;
assign micromatrizz[81][491] = 9'b111111111;
assign micromatrizz[81][492] = 9'b111111111;
assign micromatrizz[81][493] = 9'b111111111;
assign micromatrizz[81][494] = 9'b111111111;
assign micromatrizz[81][495] = 9'b111111111;
assign micromatrizz[81][496] = 9'b111111111;
assign micromatrizz[81][497] = 9'b111111111;
assign micromatrizz[81][498] = 9'b111111111;
assign micromatrizz[81][499] = 9'b111111111;
assign micromatrizz[81][500] = 9'b111111111;
assign micromatrizz[81][501] = 9'b111111111;
assign micromatrizz[81][502] = 9'b111111111;
assign micromatrizz[81][503] = 9'b111111111;
assign micromatrizz[81][504] = 9'b111111111;
assign micromatrizz[81][505] = 9'b111111111;
assign micromatrizz[81][506] = 9'b111111111;
assign micromatrizz[81][507] = 9'b111111111;
assign micromatrizz[81][508] = 9'b111111111;
assign micromatrizz[81][509] = 9'b111111111;
assign micromatrizz[81][510] = 9'b111111111;
assign micromatrizz[81][511] = 9'b111111111;
assign micromatrizz[81][512] = 9'b111111111;
assign micromatrizz[81][513] = 9'b111111111;
assign micromatrizz[81][514] = 9'b111111111;
assign micromatrizz[81][515] = 9'b111111111;
assign micromatrizz[81][516] = 9'b111111111;
assign micromatrizz[81][517] = 9'b111111111;
assign micromatrizz[81][518] = 9'b111111111;
assign micromatrizz[81][519] = 9'b111111111;
assign micromatrizz[81][520] = 9'b111111111;
assign micromatrizz[81][521] = 9'b111111111;
assign micromatrizz[81][522] = 9'b111111111;
assign micromatrizz[81][523] = 9'b111111111;
assign micromatrizz[81][524] = 9'b111111111;
assign micromatrizz[81][525] = 9'b111111111;
assign micromatrizz[81][526] = 9'b111111111;
assign micromatrizz[81][527] = 9'b111111111;
assign micromatrizz[81][528] = 9'b111111111;
assign micromatrizz[81][529] = 9'b111111111;
assign micromatrizz[81][530] = 9'b111111111;
assign micromatrizz[81][531] = 9'b111111111;
assign micromatrizz[81][532] = 9'b111111111;
assign micromatrizz[81][533] = 9'b111111111;
assign micromatrizz[81][534] = 9'b111111111;
assign micromatrizz[81][535] = 9'b111111111;
assign micromatrizz[81][536] = 9'b111111111;
assign micromatrizz[81][537] = 9'b111111111;
assign micromatrizz[81][538] = 9'b111111111;
assign micromatrizz[81][539] = 9'b111111111;
assign micromatrizz[81][540] = 9'b111111111;
assign micromatrizz[81][541] = 9'b111111111;
assign micromatrizz[81][542] = 9'b111111111;
assign micromatrizz[81][543] = 9'b111111111;
assign micromatrizz[81][544] = 9'b111111111;
assign micromatrizz[81][545] = 9'b111111111;
assign micromatrizz[81][546] = 9'b111111111;
assign micromatrizz[81][547] = 9'b111111111;
assign micromatrizz[81][548] = 9'b111111111;
assign micromatrizz[81][549] = 9'b111111111;
assign micromatrizz[81][550] = 9'b111111111;
assign micromatrizz[81][551] = 9'b111111111;
assign micromatrizz[81][552] = 9'b111111111;
assign micromatrizz[81][553] = 9'b111111111;
assign micromatrizz[81][554] = 9'b111111111;
assign micromatrizz[81][555] = 9'b111111111;
assign micromatrizz[81][556] = 9'b111111111;
assign micromatrizz[81][557] = 9'b111111111;
assign micromatrizz[81][558] = 9'b111111111;
assign micromatrizz[81][559] = 9'b111111111;
assign micromatrizz[81][560] = 9'b111111111;
assign micromatrizz[81][561] = 9'b111111111;
assign micromatrizz[81][562] = 9'b111111111;
assign micromatrizz[81][563] = 9'b111111111;
assign micromatrizz[81][564] = 9'b111111111;
assign micromatrizz[81][565] = 9'b111111111;
assign micromatrizz[81][566] = 9'b111111111;
assign micromatrizz[81][567] = 9'b111111111;
assign micromatrizz[81][568] = 9'b111111111;
assign micromatrizz[81][569] = 9'b111111111;
assign micromatrizz[81][570] = 9'b111111111;
assign micromatrizz[81][571] = 9'b111111111;
assign micromatrizz[81][572] = 9'b111111111;
assign micromatrizz[81][573] = 9'b111111111;
assign micromatrizz[81][574] = 9'b111111111;
assign micromatrizz[81][575] = 9'b111111111;
assign micromatrizz[81][576] = 9'b111111111;
assign micromatrizz[81][577] = 9'b111111111;
assign micromatrizz[81][578] = 9'b111111111;
assign micromatrizz[81][579] = 9'b111111111;
assign micromatrizz[81][580] = 9'b111111111;
assign micromatrizz[81][581] = 9'b111111111;
assign micromatrizz[81][582] = 9'b111111111;
assign micromatrizz[81][583] = 9'b111111111;
assign micromatrizz[81][584] = 9'b111111111;
assign micromatrizz[81][585] = 9'b111111111;
assign micromatrizz[81][586] = 9'b111111111;
assign micromatrizz[81][587] = 9'b111111111;
assign micromatrizz[81][588] = 9'b111111111;
assign micromatrizz[81][589] = 9'b111111111;
assign micromatrizz[81][590] = 9'b111111111;
assign micromatrizz[81][591] = 9'b111111111;
assign micromatrizz[81][592] = 9'b111111111;
assign micromatrizz[81][593] = 9'b111111111;
assign micromatrizz[81][594] = 9'b111111111;
assign micromatrizz[81][595] = 9'b111111111;
assign micromatrizz[81][596] = 9'b111111111;
assign micromatrizz[81][597] = 9'b111111111;
assign micromatrizz[81][598] = 9'b111111111;
assign micromatrizz[81][599] = 9'b111111111;
assign micromatrizz[81][600] = 9'b111111111;
assign micromatrizz[81][601] = 9'b111111111;
assign micromatrizz[81][602] = 9'b111111111;
assign micromatrizz[81][603] = 9'b111111111;
assign micromatrizz[81][604] = 9'b111111111;
assign micromatrizz[81][605] = 9'b111111111;
assign micromatrizz[81][606] = 9'b111111111;
assign micromatrizz[81][607] = 9'b111111111;
assign micromatrizz[81][608] = 9'b111111111;
assign micromatrizz[81][609] = 9'b111111111;
assign micromatrizz[81][610] = 9'b111111111;
assign micromatrizz[81][611] = 9'b111111111;
assign micromatrizz[81][612] = 9'b111111111;
assign micromatrizz[81][613] = 9'b111111111;
assign micromatrizz[81][614] = 9'b111111111;
assign micromatrizz[81][615] = 9'b111111111;
assign micromatrizz[81][616] = 9'b111111111;
assign micromatrizz[81][617] = 9'b111111111;
assign micromatrizz[81][618] = 9'b111111111;
assign micromatrizz[81][619] = 9'b111111111;
assign micromatrizz[81][620] = 9'b111111111;
assign micromatrizz[81][621] = 9'b111111111;
assign micromatrizz[81][622] = 9'b111111111;
assign micromatrizz[81][623] = 9'b111111111;
assign micromatrizz[81][624] = 9'b111111111;
assign micromatrizz[81][625] = 9'b111111111;
assign micromatrizz[81][626] = 9'b111111111;
assign micromatrizz[81][627] = 9'b111111111;
assign micromatrizz[81][628] = 9'b111111111;
assign micromatrizz[81][629] = 9'b111111111;
assign micromatrizz[81][630] = 9'b111111111;
assign micromatrizz[81][631] = 9'b111111111;
assign micromatrizz[81][632] = 9'b111111111;
assign micromatrizz[81][633] = 9'b111111111;
assign micromatrizz[81][634] = 9'b111111111;
assign micromatrizz[81][635] = 9'b111111111;
assign micromatrizz[81][636] = 9'b111111111;
assign micromatrizz[81][637] = 9'b111111111;
assign micromatrizz[81][638] = 9'b111111111;
assign micromatrizz[81][639] = 9'b111111111;
assign micromatrizz[82][0] = 9'b111111111;
assign micromatrizz[82][1] = 9'b111111111;
assign micromatrizz[82][2] = 9'b111111111;
assign micromatrizz[82][3] = 9'b111111111;
assign micromatrizz[82][4] = 9'b111111111;
assign micromatrizz[82][5] = 9'b111111111;
assign micromatrizz[82][6] = 9'b111111111;
assign micromatrizz[82][7] = 9'b111111111;
assign micromatrizz[82][8] = 9'b111111111;
assign micromatrizz[82][9] = 9'b111111111;
assign micromatrizz[82][10] = 9'b111111111;
assign micromatrizz[82][11] = 9'b111111111;
assign micromatrizz[82][12] = 9'b111111111;
assign micromatrizz[82][13] = 9'b111111111;
assign micromatrizz[82][14] = 9'b111111111;
assign micromatrizz[82][15] = 9'b111111111;
assign micromatrizz[82][16] = 9'b111111111;
assign micromatrizz[82][17] = 9'b111111111;
assign micromatrizz[82][18] = 9'b111111111;
assign micromatrizz[82][19] = 9'b111111111;
assign micromatrizz[82][20] = 9'b111111111;
assign micromatrizz[82][21] = 9'b111111111;
assign micromatrizz[82][22] = 9'b111111111;
assign micromatrizz[82][23] = 9'b111111111;
assign micromatrizz[82][24] = 9'b111111111;
assign micromatrizz[82][25] = 9'b111111111;
assign micromatrizz[82][26] = 9'b111111111;
assign micromatrizz[82][27] = 9'b111111111;
assign micromatrizz[82][28] = 9'b111111111;
assign micromatrizz[82][29] = 9'b111111111;
assign micromatrizz[82][30] = 9'b111111111;
assign micromatrizz[82][31] = 9'b111111111;
assign micromatrizz[82][32] = 9'b111111111;
assign micromatrizz[82][33] = 9'b111111111;
assign micromatrizz[82][34] = 9'b111111111;
assign micromatrizz[82][35] = 9'b111111111;
assign micromatrizz[82][36] = 9'b111111111;
assign micromatrizz[82][37] = 9'b111111111;
assign micromatrizz[82][38] = 9'b111111111;
assign micromatrizz[82][39] = 9'b111111111;
assign micromatrizz[82][40] = 9'b111111111;
assign micromatrizz[82][41] = 9'b111111111;
assign micromatrizz[82][42] = 9'b111111111;
assign micromatrizz[82][43] = 9'b111111111;
assign micromatrizz[82][44] = 9'b111111111;
assign micromatrizz[82][45] = 9'b111111111;
assign micromatrizz[82][46] = 9'b111111111;
assign micromatrizz[82][47] = 9'b111111111;
assign micromatrizz[82][48] = 9'b111111111;
assign micromatrizz[82][49] = 9'b111111111;
assign micromatrizz[82][50] = 9'b111111111;
assign micromatrizz[82][51] = 9'b111111111;
assign micromatrizz[82][52] = 9'b111111111;
assign micromatrizz[82][53] = 9'b111111111;
assign micromatrizz[82][54] = 9'b111111111;
assign micromatrizz[82][55] = 9'b111111111;
assign micromatrizz[82][56] = 9'b111111111;
assign micromatrizz[82][57] = 9'b111111111;
assign micromatrizz[82][58] = 9'b111111111;
assign micromatrizz[82][59] = 9'b111111111;
assign micromatrizz[82][60] = 9'b111111111;
assign micromatrizz[82][61] = 9'b111111111;
assign micromatrizz[82][62] = 9'b111111111;
assign micromatrizz[82][63] = 9'b111111111;
assign micromatrizz[82][64] = 9'b111111111;
assign micromatrizz[82][65] = 9'b111111111;
assign micromatrizz[82][66] = 9'b111111111;
assign micromatrizz[82][67] = 9'b111111111;
assign micromatrizz[82][68] = 9'b111111111;
assign micromatrizz[82][69] = 9'b111111111;
assign micromatrizz[82][70] = 9'b111111111;
assign micromatrizz[82][71] = 9'b111111111;
assign micromatrizz[82][72] = 9'b111111111;
assign micromatrizz[82][73] = 9'b111111111;
assign micromatrizz[82][74] = 9'b111111111;
assign micromatrizz[82][75] = 9'b111111111;
assign micromatrizz[82][76] = 9'b111111111;
assign micromatrizz[82][77] = 9'b111111111;
assign micromatrizz[82][78] = 9'b111111111;
assign micromatrizz[82][79] = 9'b111111111;
assign micromatrizz[82][80] = 9'b111111111;
assign micromatrizz[82][81] = 9'b111111111;
assign micromatrizz[82][82] = 9'b111111111;
assign micromatrizz[82][83] = 9'b111111111;
assign micromatrizz[82][84] = 9'b111111111;
assign micromatrizz[82][85] = 9'b111111111;
assign micromatrizz[82][86] = 9'b111111111;
assign micromatrizz[82][87] = 9'b111111111;
assign micromatrizz[82][88] = 9'b111111111;
assign micromatrizz[82][89] = 9'b111111111;
assign micromatrizz[82][90] = 9'b111111111;
assign micromatrizz[82][91] = 9'b111111111;
assign micromatrizz[82][92] = 9'b111111111;
assign micromatrizz[82][93] = 9'b111111111;
assign micromatrizz[82][94] = 9'b111111111;
assign micromatrizz[82][95] = 9'b111111111;
assign micromatrizz[82][96] = 9'b111111111;
assign micromatrizz[82][97] = 9'b111111111;
assign micromatrizz[82][98] = 9'b111111111;
assign micromatrizz[82][99] = 9'b111111111;
assign micromatrizz[82][100] = 9'b111111111;
assign micromatrizz[82][101] = 9'b111111111;
assign micromatrizz[82][102] = 9'b111111111;
assign micromatrizz[82][103] = 9'b111111111;
assign micromatrizz[82][104] = 9'b111111111;
assign micromatrizz[82][105] = 9'b111111111;
assign micromatrizz[82][106] = 9'b111111111;
assign micromatrizz[82][107] = 9'b111111111;
assign micromatrizz[82][108] = 9'b111111111;
assign micromatrizz[82][109] = 9'b111111111;
assign micromatrizz[82][110] = 9'b111111111;
assign micromatrizz[82][111] = 9'b111111111;
assign micromatrizz[82][112] = 9'b111111111;
assign micromatrizz[82][113] = 9'b111111111;
assign micromatrizz[82][114] = 9'b111111111;
assign micromatrizz[82][115] = 9'b111111111;
assign micromatrizz[82][116] = 9'b111111111;
assign micromatrizz[82][117] = 9'b111111111;
assign micromatrizz[82][118] = 9'b111111111;
assign micromatrizz[82][119] = 9'b111111111;
assign micromatrizz[82][120] = 9'b111111111;
assign micromatrizz[82][121] = 9'b111111111;
assign micromatrizz[82][122] = 9'b111111111;
assign micromatrizz[82][123] = 9'b111111111;
assign micromatrizz[82][124] = 9'b111111111;
assign micromatrizz[82][125] = 9'b111111111;
assign micromatrizz[82][126] = 9'b111111111;
assign micromatrizz[82][127] = 9'b111111111;
assign micromatrizz[82][128] = 9'b111111111;
assign micromatrizz[82][129] = 9'b111111111;
assign micromatrizz[82][130] = 9'b111111111;
assign micromatrizz[82][131] = 9'b111111111;
assign micromatrizz[82][132] = 9'b111111111;
assign micromatrizz[82][133] = 9'b111111111;
assign micromatrizz[82][134] = 9'b111111111;
assign micromatrizz[82][135] = 9'b111111111;
assign micromatrizz[82][136] = 9'b111111111;
assign micromatrizz[82][137] = 9'b111111111;
assign micromatrizz[82][138] = 9'b111111111;
assign micromatrizz[82][139] = 9'b111111111;
assign micromatrizz[82][140] = 9'b111111111;
assign micromatrizz[82][141] = 9'b111111111;
assign micromatrizz[82][142] = 9'b111111111;
assign micromatrizz[82][143] = 9'b111111111;
assign micromatrizz[82][144] = 9'b111111111;
assign micromatrizz[82][145] = 9'b111111111;
assign micromatrizz[82][146] = 9'b111111111;
assign micromatrizz[82][147] = 9'b111111111;
assign micromatrizz[82][148] = 9'b111111111;
assign micromatrizz[82][149] = 9'b111111111;
assign micromatrizz[82][150] = 9'b111111111;
assign micromatrizz[82][151] = 9'b111111111;
assign micromatrizz[82][152] = 9'b111111111;
assign micromatrizz[82][153] = 9'b111111111;
assign micromatrizz[82][154] = 9'b111111111;
assign micromatrizz[82][155] = 9'b111111111;
assign micromatrizz[82][156] = 9'b111111111;
assign micromatrizz[82][157] = 9'b111111111;
assign micromatrizz[82][158] = 9'b111111111;
assign micromatrizz[82][159] = 9'b111111111;
assign micromatrizz[82][160] = 9'b111111111;
assign micromatrizz[82][161] = 9'b111111111;
assign micromatrizz[82][162] = 9'b111111111;
assign micromatrizz[82][163] = 9'b111111111;
assign micromatrizz[82][164] = 9'b111111111;
assign micromatrizz[82][165] = 9'b111111111;
assign micromatrizz[82][166] = 9'b111111111;
assign micromatrizz[82][167] = 9'b111111111;
assign micromatrizz[82][168] = 9'b111111111;
assign micromatrizz[82][169] = 9'b111111111;
assign micromatrizz[82][170] = 9'b111111111;
assign micromatrizz[82][171] = 9'b111111111;
assign micromatrizz[82][172] = 9'b111111111;
assign micromatrizz[82][173] = 9'b111111111;
assign micromatrizz[82][174] = 9'b111111111;
assign micromatrizz[82][175] = 9'b111111111;
assign micromatrizz[82][176] = 9'b111111111;
assign micromatrizz[82][177] = 9'b111111111;
assign micromatrizz[82][178] = 9'b111111111;
assign micromatrizz[82][179] = 9'b111111111;
assign micromatrizz[82][180] = 9'b111111111;
assign micromatrizz[82][181] = 9'b111111111;
assign micromatrizz[82][182] = 9'b111111111;
assign micromatrizz[82][183] = 9'b111111111;
assign micromatrizz[82][184] = 9'b111111111;
assign micromatrizz[82][185] = 9'b111111111;
assign micromatrizz[82][186] = 9'b111111111;
assign micromatrizz[82][187] = 9'b111111111;
assign micromatrizz[82][188] = 9'b111111111;
assign micromatrizz[82][189] = 9'b111111111;
assign micromatrizz[82][190] = 9'b111111111;
assign micromatrizz[82][191] = 9'b111111111;
assign micromatrizz[82][192] = 9'b111111111;
assign micromatrizz[82][193] = 9'b111111111;
assign micromatrizz[82][194] = 9'b111111111;
assign micromatrizz[82][195] = 9'b111111111;
assign micromatrizz[82][196] = 9'b111111111;
assign micromatrizz[82][197] = 9'b111111111;
assign micromatrizz[82][198] = 9'b111111111;
assign micromatrizz[82][199] = 9'b111111111;
assign micromatrizz[82][200] = 9'b111111111;
assign micromatrizz[82][201] = 9'b111111111;
assign micromatrizz[82][202] = 9'b111111111;
assign micromatrizz[82][203] = 9'b111111111;
assign micromatrizz[82][204] = 9'b111111111;
assign micromatrizz[82][205] = 9'b111111111;
assign micromatrizz[82][206] = 9'b111111111;
assign micromatrizz[82][207] = 9'b111111111;
assign micromatrizz[82][208] = 9'b111111111;
assign micromatrizz[82][209] = 9'b111111111;
assign micromatrizz[82][210] = 9'b111111111;
assign micromatrizz[82][211] = 9'b111111111;
assign micromatrizz[82][212] = 9'b111111111;
assign micromatrizz[82][213] = 9'b111111111;
assign micromatrizz[82][214] = 9'b111111111;
assign micromatrizz[82][215] = 9'b111111111;
assign micromatrizz[82][216] = 9'b111111111;
assign micromatrizz[82][217] = 9'b111111111;
assign micromatrizz[82][218] = 9'b111111111;
assign micromatrizz[82][219] = 9'b111111111;
assign micromatrizz[82][220] = 9'b111111111;
assign micromatrizz[82][221] = 9'b111111111;
assign micromatrizz[82][222] = 9'b111111111;
assign micromatrizz[82][223] = 9'b111111111;
assign micromatrizz[82][224] = 9'b111111111;
assign micromatrizz[82][225] = 9'b111111111;
assign micromatrizz[82][226] = 9'b111111111;
assign micromatrizz[82][227] = 9'b111111111;
assign micromatrizz[82][228] = 9'b111111111;
assign micromatrizz[82][229] = 9'b111111111;
assign micromatrizz[82][230] = 9'b111111111;
assign micromatrizz[82][231] = 9'b111111111;
assign micromatrizz[82][232] = 9'b111111111;
assign micromatrizz[82][233] = 9'b111111111;
assign micromatrizz[82][234] = 9'b111111111;
assign micromatrizz[82][235] = 9'b111111111;
assign micromatrizz[82][236] = 9'b111111111;
assign micromatrizz[82][237] = 9'b111111111;
assign micromatrizz[82][238] = 9'b111111111;
assign micromatrizz[82][239] = 9'b111111111;
assign micromatrizz[82][240] = 9'b111111111;
assign micromatrizz[82][241] = 9'b111111111;
assign micromatrizz[82][242] = 9'b111111111;
assign micromatrizz[82][243] = 9'b111111111;
assign micromatrizz[82][244] = 9'b111111111;
assign micromatrizz[82][245] = 9'b111111111;
assign micromatrizz[82][246] = 9'b111111111;
assign micromatrizz[82][247] = 9'b111111111;
assign micromatrizz[82][248] = 9'b111111111;
assign micromatrizz[82][249] = 9'b111111111;
assign micromatrizz[82][250] = 9'b111111111;
assign micromatrizz[82][251] = 9'b111111111;
assign micromatrizz[82][252] = 9'b111111111;
assign micromatrizz[82][253] = 9'b111111111;
assign micromatrizz[82][254] = 9'b111111111;
assign micromatrizz[82][255] = 9'b111111111;
assign micromatrizz[82][256] = 9'b111111111;
assign micromatrizz[82][257] = 9'b111111111;
assign micromatrizz[82][258] = 9'b111111111;
assign micromatrizz[82][259] = 9'b111111111;
assign micromatrizz[82][260] = 9'b111111111;
assign micromatrizz[82][261] = 9'b111111111;
assign micromatrizz[82][262] = 9'b111111111;
assign micromatrizz[82][263] = 9'b111111111;
assign micromatrizz[82][264] = 9'b111111111;
assign micromatrizz[82][265] = 9'b111111111;
assign micromatrizz[82][266] = 9'b111111111;
assign micromatrizz[82][267] = 9'b111111111;
assign micromatrizz[82][268] = 9'b111111111;
assign micromatrizz[82][269] = 9'b111111111;
assign micromatrizz[82][270] = 9'b111111111;
assign micromatrizz[82][271] = 9'b111111111;
assign micromatrizz[82][272] = 9'b111111111;
assign micromatrizz[82][273] = 9'b111111111;
assign micromatrizz[82][274] = 9'b111111111;
assign micromatrizz[82][275] = 9'b111111111;
assign micromatrizz[82][276] = 9'b111111111;
assign micromatrizz[82][277] = 9'b111111111;
assign micromatrizz[82][278] = 9'b111111111;
assign micromatrizz[82][279] = 9'b111111111;
assign micromatrizz[82][280] = 9'b111111111;
assign micromatrizz[82][281] = 9'b111111111;
assign micromatrizz[82][282] = 9'b111111111;
assign micromatrizz[82][283] = 9'b111111111;
assign micromatrizz[82][284] = 9'b111111111;
assign micromatrizz[82][285] = 9'b111111111;
assign micromatrizz[82][286] = 9'b111111111;
assign micromatrizz[82][287] = 9'b111111111;
assign micromatrizz[82][288] = 9'b111111111;
assign micromatrizz[82][289] = 9'b111111111;
assign micromatrizz[82][290] = 9'b111111111;
assign micromatrizz[82][291] = 9'b111111111;
assign micromatrizz[82][292] = 9'b111111111;
assign micromatrizz[82][293] = 9'b111111111;
assign micromatrizz[82][294] = 9'b111111111;
assign micromatrizz[82][295] = 9'b111111111;
assign micromatrizz[82][296] = 9'b111111111;
assign micromatrizz[82][297] = 9'b111111111;
assign micromatrizz[82][298] = 9'b111111111;
assign micromatrizz[82][299] = 9'b111111111;
assign micromatrizz[82][300] = 9'b111111111;
assign micromatrizz[82][301] = 9'b111111111;
assign micromatrizz[82][302] = 9'b111111111;
assign micromatrizz[82][303] = 9'b111111111;
assign micromatrizz[82][304] = 9'b111111111;
assign micromatrizz[82][305] = 9'b111111111;
assign micromatrizz[82][306] = 9'b111111111;
assign micromatrizz[82][307] = 9'b111111111;
assign micromatrizz[82][308] = 9'b111111111;
assign micromatrizz[82][309] = 9'b111111111;
assign micromatrizz[82][310] = 9'b111111111;
assign micromatrizz[82][311] = 9'b111111111;
assign micromatrizz[82][312] = 9'b111111111;
assign micromatrizz[82][313] = 9'b111111111;
assign micromatrizz[82][314] = 9'b111111111;
assign micromatrizz[82][315] = 9'b111111111;
assign micromatrizz[82][316] = 9'b111111111;
assign micromatrizz[82][317] = 9'b111111111;
assign micromatrizz[82][318] = 9'b111111111;
assign micromatrizz[82][319] = 9'b111111111;
assign micromatrizz[82][320] = 9'b111111111;
assign micromatrizz[82][321] = 9'b111111111;
assign micromatrizz[82][322] = 9'b111111111;
assign micromatrizz[82][323] = 9'b111111111;
assign micromatrizz[82][324] = 9'b111111111;
assign micromatrizz[82][325] = 9'b111111111;
assign micromatrizz[82][326] = 9'b111111111;
assign micromatrizz[82][327] = 9'b111111111;
assign micromatrizz[82][328] = 9'b111111111;
assign micromatrizz[82][329] = 9'b111111111;
assign micromatrizz[82][330] = 9'b111111111;
assign micromatrizz[82][331] = 9'b111111111;
assign micromatrizz[82][332] = 9'b111111111;
assign micromatrizz[82][333] = 9'b111111111;
assign micromatrizz[82][334] = 9'b111111111;
assign micromatrizz[82][335] = 9'b111111111;
assign micromatrizz[82][336] = 9'b111111111;
assign micromatrizz[82][337] = 9'b111111111;
assign micromatrizz[82][338] = 9'b111111111;
assign micromatrizz[82][339] = 9'b111111111;
assign micromatrizz[82][340] = 9'b111111111;
assign micromatrizz[82][341] = 9'b111111111;
assign micromatrizz[82][342] = 9'b111111111;
assign micromatrizz[82][343] = 9'b111111111;
assign micromatrizz[82][344] = 9'b111111111;
assign micromatrizz[82][345] = 9'b111111111;
assign micromatrizz[82][346] = 9'b111111111;
assign micromatrizz[82][347] = 9'b111111111;
assign micromatrizz[82][348] = 9'b111111111;
assign micromatrizz[82][349] = 9'b111111111;
assign micromatrizz[82][350] = 9'b111111111;
assign micromatrizz[82][351] = 9'b111111111;
assign micromatrizz[82][352] = 9'b111111111;
assign micromatrizz[82][353] = 9'b111111111;
assign micromatrizz[82][354] = 9'b111111111;
assign micromatrizz[82][355] = 9'b111111111;
assign micromatrizz[82][356] = 9'b111111111;
assign micromatrizz[82][357] = 9'b111111111;
assign micromatrizz[82][358] = 9'b111111111;
assign micromatrizz[82][359] = 9'b111111111;
assign micromatrizz[82][360] = 9'b111111111;
assign micromatrizz[82][361] = 9'b111111111;
assign micromatrizz[82][362] = 9'b111111111;
assign micromatrizz[82][363] = 9'b111111111;
assign micromatrizz[82][364] = 9'b111111111;
assign micromatrizz[82][365] = 9'b111111111;
assign micromatrizz[82][366] = 9'b111111111;
assign micromatrizz[82][367] = 9'b111111111;
assign micromatrizz[82][368] = 9'b111111111;
assign micromatrizz[82][369] = 9'b111111111;
assign micromatrizz[82][370] = 9'b111111111;
assign micromatrizz[82][371] = 9'b111111111;
assign micromatrizz[82][372] = 9'b111111111;
assign micromatrizz[82][373] = 9'b111111111;
assign micromatrizz[82][374] = 9'b111111111;
assign micromatrizz[82][375] = 9'b111111111;
assign micromatrizz[82][376] = 9'b111111111;
assign micromatrizz[82][377] = 9'b111111111;
assign micromatrizz[82][378] = 9'b111111111;
assign micromatrizz[82][379] = 9'b111111111;
assign micromatrizz[82][380] = 9'b111111111;
assign micromatrizz[82][381] = 9'b111111111;
assign micromatrizz[82][382] = 9'b111111111;
assign micromatrizz[82][383] = 9'b111111111;
assign micromatrizz[82][384] = 9'b111111111;
assign micromatrizz[82][385] = 9'b111111111;
assign micromatrizz[82][386] = 9'b111111111;
assign micromatrizz[82][387] = 9'b111111111;
assign micromatrizz[82][388] = 9'b111111111;
assign micromatrizz[82][389] = 9'b111111111;
assign micromatrizz[82][390] = 9'b111111111;
assign micromatrizz[82][391] = 9'b111111111;
assign micromatrizz[82][392] = 9'b111111111;
assign micromatrizz[82][393] = 9'b111111111;
assign micromatrizz[82][394] = 9'b111111111;
assign micromatrizz[82][395] = 9'b111111111;
assign micromatrizz[82][396] = 9'b111111111;
assign micromatrizz[82][397] = 9'b111111111;
assign micromatrizz[82][398] = 9'b111111111;
assign micromatrizz[82][399] = 9'b111111111;
assign micromatrizz[82][400] = 9'b111111111;
assign micromatrizz[82][401] = 9'b111111111;
assign micromatrizz[82][402] = 9'b111111111;
assign micromatrizz[82][403] = 9'b111111111;
assign micromatrizz[82][404] = 9'b111111111;
assign micromatrizz[82][405] = 9'b111111111;
assign micromatrizz[82][406] = 9'b111111111;
assign micromatrizz[82][407] = 9'b111111111;
assign micromatrizz[82][408] = 9'b111111111;
assign micromatrizz[82][409] = 9'b111111111;
assign micromatrizz[82][410] = 9'b111111111;
assign micromatrizz[82][411] = 9'b111111111;
assign micromatrizz[82][412] = 9'b111111111;
assign micromatrizz[82][413] = 9'b111111111;
assign micromatrizz[82][414] = 9'b111111111;
assign micromatrizz[82][415] = 9'b111111111;
assign micromatrizz[82][416] = 9'b111111111;
assign micromatrizz[82][417] = 9'b111111111;
assign micromatrizz[82][418] = 9'b111111111;
assign micromatrizz[82][419] = 9'b111111111;
assign micromatrizz[82][420] = 9'b111111111;
assign micromatrizz[82][421] = 9'b111111111;
assign micromatrizz[82][422] = 9'b111111111;
assign micromatrizz[82][423] = 9'b111111111;
assign micromatrizz[82][424] = 9'b111111111;
assign micromatrizz[82][425] = 9'b111111111;
assign micromatrizz[82][426] = 9'b111111111;
assign micromatrizz[82][427] = 9'b111111111;
assign micromatrizz[82][428] = 9'b111111111;
assign micromatrizz[82][429] = 9'b111111111;
assign micromatrizz[82][430] = 9'b111111111;
assign micromatrizz[82][431] = 9'b111111111;
assign micromatrizz[82][432] = 9'b111111111;
assign micromatrizz[82][433] = 9'b111111111;
assign micromatrizz[82][434] = 9'b111111111;
assign micromatrizz[82][435] = 9'b111111111;
assign micromatrizz[82][436] = 9'b111111111;
assign micromatrizz[82][437] = 9'b111111111;
assign micromatrizz[82][438] = 9'b111111111;
assign micromatrizz[82][439] = 9'b111111111;
assign micromatrizz[82][440] = 9'b111111111;
assign micromatrizz[82][441] = 9'b111111111;
assign micromatrizz[82][442] = 9'b111111111;
assign micromatrizz[82][443] = 9'b111111111;
assign micromatrizz[82][444] = 9'b111111111;
assign micromatrizz[82][445] = 9'b111111111;
assign micromatrizz[82][446] = 9'b111111111;
assign micromatrizz[82][447] = 9'b111111111;
assign micromatrizz[82][448] = 9'b111111111;
assign micromatrizz[82][449] = 9'b111111111;
assign micromatrizz[82][450] = 9'b111111111;
assign micromatrizz[82][451] = 9'b111111111;
assign micromatrizz[82][452] = 9'b111111111;
assign micromatrizz[82][453] = 9'b111111111;
assign micromatrizz[82][454] = 9'b111111111;
assign micromatrizz[82][455] = 9'b111111111;
assign micromatrizz[82][456] = 9'b111111111;
assign micromatrizz[82][457] = 9'b111111111;
assign micromatrizz[82][458] = 9'b111111111;
assign micromatrizz[82][459] = 9'b111111111;
assign micromatrizz[82][460] = 9'b111111111;
assign micromatrizz[82][461] = 9'b111111111;
assign micromatrizz[82][462] = 9'b111111111;
assign micromatrizz[82][463] = 9'b111111111;
assign micromatrizz[82][464] = 9'b111111111;
assign micromatrizz[82][465] = 9'b111111111;
assign micromatrizz[82][466] = 9'b111111111;
assign micromatrizz[82][467] = 9'b111111111;
assign micromatrizz[82][468] = 9'b111111111;
assign micromatrizz[82][469] = 9'b111111111;
assign micromatrizz[82][470] = 9'b111111111;
assign micromatrizz[82][471] = 9'b111111111;
assign micromatrizz[82][472] = 9'b111111111;
assign micromatrizz[82][473] = 9'b111111111;
assign micromatrizz[82][474] = 9'b111111111;
assign micromatrizz[82][475] = 9'b111111111;
assign micromatrizz[82][476] = 9'b111111111;
assign micromatrizz[82][477] = 9'b111111111;
assign micromatrizz[82][478] = 9'b111111111;
assign micromatrizz[82][479] = 9'b111111111;
assign micromatrizz[82][480] = 9'b111111111;
assign micromatrizz[82][481] = 9'b111111111;
assign micromatrizz[82][482] = 9'b111111111;
assign micromatrizz[82][483] = 9'b111111111;
assign micromatrizz[82][484] = 9'b111111111;
assign micromatrizz[82][485] = 9'b111111111;
assign micromatrizz[82][486] = 9'b111111111;
assign micromatrizz[82][487] = 9'b111111111;
assign micromatrizz[82][488] = 9'b111111111;
assign micromatrizz[82][489] = 9'b111111111;
assign micromatrizz[82][490] = 9'b111111111;
assign micromatrizz[82][491] = 9'b111111111;
assign micromatrizz[82][492] = 9'b111111111;
assign micromatrizz[82][493] = 9'b111111111;
assign micromatrizz[82][494] = 9'b111111111;
assign micromatrizz[82][495] = 9'b111111111;
assign micromatrizz[82][496] = 9'b111111111;
assign micromatrizz[82][497] = 9'b111111111;
assign micromatrizz[82][498] = 9'b111111111;
assign micromatrizz[82][499] = 9'b111111111;
assign micromatrizz[82][500] = 9'b111111111;
assign micromatrizz[82][501] = 9'b111111111;
assign micromatrizz[82][502] = 9'b111111111;
assign micromatrizz[82][503] = 9'b111111111;
assign micromatrizz[82][504] = 9'b111111111;
assign micromatrizz[82][505] = 9'b111111111;
assign micromatrizz[82][506] = 9'b111111111;
assign micromatrizz[82][507] = 9'b111111111;
assign micromatrizz[82][508] = 9'b111111111;
assign micromatrizz[82][509] = 9'b111111111;
assign micromatrizz[82][510] = 9'b111111111;
assign micromatrizz[82][511] = 9'b111111111;
assign micromatrizz[82][512] = 9'b111111111;
assign micromatrizz[82][513] = 9'b111111111;
assign micromatrizz[82][514] = 9'b111111111;
assign micromatrizz[82][515] = 9'b111111111;
assign micromatrizz[82][516] = 9'b111111111;
assign micromatrizz[82][517] = 9'b111111111;
assign micromatrizz[82][518] = 9'b111111111;
assign micromatrizz[82][519] = 9'b111111111;
assign micromatrizz[82][520] = 9'b111111111;
assign micromatrizz[82][521] = 9'b111111111;
assign micromatrizz[82][522] = 9'b111111111;
assign micromatrizz[82][523] = 9'b111111111;
assign micromatrizz[82][524] = 9'b111111111;
assign micromatrizz[82][525] = 9'b111111111;
assign micromatrizz[82][526] = 9'b111111111;
assign micromatrizz[82][527] = 9'b111111111;
assign micromatrizz[82][528] = 9'b111111111;
assign micromatrizz[82][529] = 9'b111111111;
assign micromatrizz[82][530] = 9'b111111111;
assign micromatrizz[82][531] = 9'b111111111;
assign micromatrizz[82][532] = 9'b111111111;
assign micromatrizz[82][533] = 9'b111111111;
assign micromatrizz[82][534] = 9'b111111111;
assign micromatrizz[82][535] = 9'b111111111;
assign micromatrizz[82][536] = 9'b111111111;
assign micromatrizz[82][537] = 9'b111111111;
assign micromatrizz[82][538] = 9'b111111111;
assign micromatrizz[82][539] = 9'b111111111;
assign micromatrizz[82][540] = 9'b111111111;
assign micromatrizz[82][541] = 9'b111111111;
assign micromatrizz[82][542] = 9'b111111111;
assign micromatrizz[82][543] = 9'b111111111;
assign micromatrizz[82][544] = 9'b111111111;
assign micromatrizz[82][545] = 9'b111111111;
assign micromatrizz[82][546] = 9'b111111111;
assign micromatrizz[82][547] = 9'b111111111;
assign micromatrizz[82][548] = 9'b111111111;
assign micromatrizz[82][549] = 9'b111111111;
assign micromatrizz[82][550] = 9'b111111111;
assign micromatrizz[82][551] = 9'b111111111;
assign micromatrizz[82][552] = 9'b111111111;
assign micromatrizz[82][553] = 9'b111111111;
assign micromatrizz[82][554] = 9'b111111111;
assign micromatrizz[82][555] = 9'b111111111;
assign micromatrizz[82][556] = 9'b111111111;
assign micromatrizz[82][557] = 9'b111111111;
assign micromatrizz[82][558] = 9'b111111111;
assign micromatrizz[82][559] = 9'b111111111;
assign micromatrizz[82][560] = 9'b111111111;
assign micromatrizz[82][561] = 9'b111111111;
assign micromatrizz[82][562] = 9'b111111111;
assign micromatrizz[82][563] = 9'b111111111;
assign micromatrizz[82][564] = 9'b111111111;
assign micromatrizz[82][565] = 9'b111111111;
assign micromatrizz[82][566] = 9'b111111111;
assign micromatrizz[82][567] = 9'b111111111;
assign micromatrizz[82][568] = 9'b111111111;
assign micromatrizz[82][569] = 9'b111111111;
assign micromatrizz[82][570] = 9'b111111111;
assign micromatrizz[82][571] = 9'b111111111;
assign micromatrizz[82][572] = 9'b111111111;
assign micromatrizz[82][573] = 9'b111111111;
assign micromatrizz[82][574] = 9'b111111111;
assign micromatrizz[82][575] = 9'b111111111;
assign micromatrizz[82][576] = 9'b111111111;
assign micromatrizz[82][577] = 9'b111111111;
assign micromatrizz[82][578] = 9'b111111111;
assign micromatrizz[82][579] = 9'b111111111;
assign micromatrizz[82][580] = 9'b111111111;
assign micromatrizz[82][581] = 9'b111111111;
assign micromatrizz[82][582] = 9'b111111111;
assign micromatrizz[82][583] = 9'b111111111;
assign micromatrizz[82][584] = 9'b111111111;
assign micromatrizz[82][585] = 9'b111111111;
assign micromatrizz[82][586] = 9'b111111111;
assign micromatrizz[82][587] = 9'b111111111;
assign micromatrizz[82][588] = 9'b111111111;
assign micromatrizz[82][589] = 9'b111111111;
assign micromatrizz[82][590] = 9'b111111111;
assign micromatrizz[82][591] = 9'b111111111;
assign micromatrizz[82][592] = 9'b111111111;
assign micromatrizz[82][593] = 9'b111111111;
assign micromatrizz[82][594] = 9'b111111111;
assign micromatrizz[82][595] = 9'b111111111;
assign micromatrizz[82][596] = 9'b111111111;
assign micromatrizz[82][597] = 9'b111111111;
assign micromatrizz[82][598] = 9'b111111111;
assign micromatrizz[82][599] = 9'b111111111;
assign micromatrizz[82][600] = 9'b111111111;
assign micromatrizz[82][601] = 9'b111111111;
assign micromatrizz[82][602] = 9'b111111111;
assign micromatrizz[82][603] = 9'b111111111;
assign micromatrizz[82][604] = 9'b111111111;
assign micromatrizz[82][605] = 9'b111111111;
assign micromatrizz[82][606] = 9'b111111111;
assign micromatrizz[82][607] = 9'b111111111;
assign micromatrizz[82][608] = 9'b111111111;
assign micromatrizz[82][609] = 9'b111111111;
assign micromatrizz[82][610] = 9'b111111111;
assign micromatrizz[82][611] = 9'b111111111;
assign micromatrizz[82][612] = 9'b111111111;
assign micromatrizz[82][613] = 9'b111111111;
assign micromatrizz[82][614] = 9'b111111111;
assign micromatrizz[82][615] = 9'b111111111;
assign micromatrizz[82][616] = 9'b111111111;
assign micromatrizz[82][617] = 9'b111111111;
assign micromatrizz[82][618] = 9'b111111111;
assign micromatrizz[82][619] = 9'b111111111;
assign micromatrizz[82][620] = 9'b111111111;
assign micromatrizz[82][621] = 9'b111111111;
assign micromatrizz[82][622] = 9'b111111111;
assign micromatrizz[82][623] = 9'b111111111;
assign micromatrizz[82][624] = 9'b111111111;
assign micromatrizz[82][625] = 9'b111111111;
assign micromatrizz[82][626] = 9'b111111111;
assign micromatrizz[82][627] = 9'b111111111;
assign micromatrizz[82][628] = 9'b111111111;
assign micromatrizz[82][629] = 9'b111111111;
assign micromatrizz[82][630] = 9'b111111111;
assign micromatrizz[82][631] = 9'b111111111;
assign micromatrizz[82][632] = 9'b111111111;
assign micromatrizz[82][633] = 9'b111111111;
assign micromatrizz[82][634] = 9'b111111111;
assign micromatrizz[82][635] = 9'b111111111;
assign micromatrizz[82][636] = 9'b111111111;
assign micromatrizz[82][637] = 9'b111111111;
assign micromatrizz[82][638] = 9'b111111111;
assign micromatrizz[82][639] = 9'b111111111;
assign micromatrizz[83][0] = 9'b111111111;
assign micromatrizz[83][1] = 9'b111111111;
assign micromatrizz[83][2] = 9'b111111111;
assign micromatrizz[83][3] = 9'b111111111;
assign micromatrizz[83][4] = 9'b111111111;
assign micromatrizz[83][5] = 9'b111111111;
assign micromatrizz[83][6] = 9'b111111111;
assign micromatrizz[83][7] = 9'b111111111;
assign micromatrizz[83][8] = 9'b111111111;
assign micromatrizz[83][9] = 9'b111111111;
assign micromatrizz[83][10] = 9'b111111111;
assign micromatrizz[83][11] = 9'b111111111;
assign micromatrizz[83][12] = 9'b111111111;
assign micromatrizz[83][13] = 9'b111111111;
assign micromatrizz[83][14] = 9'b111111111;
assign micromatrizz[83][15] = 9'b111111111;
assign micromatrizz[83][16] = 9'b111111111;
assign micromatrizz[83][17] = 9'b111111111;
assign micromatrizz[83][18] = 9'b111111111;
assign micromatrizz[83][19] = 9'b111111111;
assign micromatrizz[83][20] = 9'b111111111;
assign micromatrizz[83][21] = 9'b111111111;
assign micromatrizz[83][22] = 9'b111111111;
assign micromatrizz[83][23] = 9'b111111111;
assign micromatrizz[83][24] = 9'b111111111;
assign micromatrizz[83][25] = 9'b111111111;
assign micromatrizz[83][26] = 9'b111111111;
assign micromatrizz[83][27] = 9'b111111111;
assign micromatrizz[83][28] = 9'b111111111;
assign micromatrizz[83][29] = 9'b111111111;
assign micromatrizz[83][30] = 9'b111111111;
assign micromatrizz[83][31] = 9'b111111111;
assign micromatrizz[83][32] = 9'b111111111;
assign micromatrizz[83][33] = 9'b111111111;
assign micromatrizz[83][34] = 9'b111111111;
assign micromatrizz[83][35] = 9'b111111111;
assign micromatrizz[83][36] = 9'b111111111;
assign micromatrizz[83][37] = 9'b111111111;
assign micromatrizz[83][38] = 9'b111111111;
assign micromatrizz[83][39] = 9'b111111111;
assign micromatrizz[83][40] = 9'b111111111;
assign micromatrizz[83][41] = 9'b111111111;
assign micromatrizz[83][42] = 9'b111111111;
assign micromatrizz[83][43] = 9'b111111111;
assign micromatrizz[83][44] = 9'b111111111;
assign micromatrizz[83][45] = 9'b111111111;
assign micromatrizz[83][46] = 9'b111111111;
assign micromatrizz[83][47] = 9'b111111111;
assign micromatrizz[83][48] = 9'b111111111;
assign micromatrizz[83][49] = 9'b111111111;
assign micromatrizz[83][50] = 9'b111111111;
assign micromatrizz[83][51] = 9'b111111111;
assign micromatrizz[83][52] = 9'b111111111;
assign micromatrizz[83][53] = 9'b111111111;
assign micromatrizz[83][54] = 9'b111111111;
assign micromatrizz[83][55] = 9'b111111111;
assign micromatrizz[83][56] = 9'b111111111;
assign micromatrizz[83][57] = 9'b111111111;
assign micromatrizz[83][58] = 9'b111111111;
assign micromatrizz[83][59] = 9'b111111111;
assign micromatrizz[83][60] = 9'b111111111;
assign micromatrizz[83][61] = 9'b111111111;
assign micromatrizz[83][62] = 9'b111111111;
assign micromatrizz[83][63] = 9'b111111111;
assign micromatrizz[83][64] = 9'b111111111;
assign micromatrizz[83][65] = 9'b111111111;
assign micromatrizz[83][66] = 9'b111111111;
assign micromatrizz[83][67] = 9'b111111111;
assign micromatrizz[83][68] = 9'b111111111;
assign micromatrizz[83][69] = 9'b111111111;
assign micromatrizz[83][70] = 9'b111111111;
assign micromatrizz[83][71] = 9'b111111111;
assign micromatrizz[83][72] = 9'b111111111;
assign micromatrizz[83][73] = 9'b111111111;
assign micromatrizz[83][74] = 9'b111111111;
assign micromatrizz[83][75] = 9'b111111111;
assign micromatrizz[83][76] = 9'b111111111;
assign micromatrizz[83][77] = 9'b111111111;
assign micromatrizz[83][78] = 9'b111111111;
assign micromatrizz[83][79] = 9'b111111111;
assign micromatrizz[83][80] = 9'b111111111;
assign micromatrizz[83][81] = 9'b111111111;
assign micromatrizz[83][82] = 9'b111111111;
assign micromatrizz[83][83] = 9'b111111111;
assign micromatrizz[83][84] = 9'b111111111;
assign micromatrizz[83][85] = 9'b111111111;
assign micromatrizz[83][86] = 9'b111111111;
assign micromatrizz[83][87] = 9'b111111111;
assign micromatrizz[83][88] = 9'b111111111;
assign micromatrizz[83][89] = 9'b111111111;
assign micromatrizz[83][90] = 9'b111111111;
assign micromatrizz[83][91] = 9'b111111111;
assign micromatrizz[83][92] = 9'b111111111;
assign micromatrizz[83][93] = 9'b111111111;
assign micromatrizz[83][94] = 9'b111111111;
assign micromatrizz[83][95] = 9'b111111111;
assign micromatrizz[83][96] = 9'b111111111;
assign micromatrizz[83][97] = 9'b111111111;
assign micromatrizz[83][98] = 9'b111111111;
assign micromatrizz[83][99] = 9'b111111111;
assign micromatrizz[83][100] = 9'b111111111;
assign micromatrizz[83][101] = 9'b111111111;
assign micromatrizz[83][102] = 9'b111111111;
assign micromatrizz[83][103] = 9'b111111111;
assign micromatrizz[83][104] = 9'b111111111;
assign micromatrizz[83][105] = 9'b111111111;
assign micromatrizz[83][106] = 9'b111111111;
assign micromatrizz[83][107] = 9'b111111111;
assign micromatrizz[83][108] = 9'b111111111;
assign micromatrizz[83][109] = 9'b111111111;
assign micromatrizz[83][110] = 9'b111111111;
assign micromatrizz[83][111] = 9'b111111111;
assign micromatrizz[83][112] = 9'b111111111;
assign micromatrizz[83][113] = 9'b111111111;
assign micromatrizz[83][114] = 9'b111111111;
assign micromatrizz[83][115] = 9'b111111111;
assign micromatrizz[83][116] = 9'b111111111;
assign micromatrizz[83][117] = 9'b111111111;
assign micromatrizz[83][118] = 9'b111111111;
assign micromatrizz[83][119] = 9'b111111111;
assign micromatrizz[83][120] = 9'b111111111;
assign micromatrizz[83][121] = 9'b111111111;
assign micromatrizz[83][122] = 9'b111111111;
assign micromatrizz[83][123] = 9'b111111111;
assign micromatrizz[83][124] = 9'b111111111;
assign micromatrizz[83][125] = 9'b111111111;
assign micromatrizz[83][126] = 9'b111111111;
assign micromatrizz[83][127] = 9'b111111111;
assign micromatrizz[83][128] = 9'b111111111;
assign micromatrizz[83][129] = 9'b111111111;
assign micromatrizz[83][130] = 9'b111111111;
assign micromatrizz[83][131] = 9'b111111111;
assign micromatrizz[83][132] = 9'b111111111;
assign micromatrizz[83][133] = 9'b111111111;
assign micromatrizz[83][134] = 9'b111111111;
assign micromatrizz[83][135] = 9'b111111111;
assign micromatrizz[83][136] = 9'b111111111;
assign micromatrizz[83][137] = 9'b111111111;
assign micromatrizz[83][138] = 9'b111111111;
assign micromatrizz[83][139] = 9'b111111111;
assign micromatrizz[83][140] = 9'b111111111;
assign micromatrizz[83][141] = 9'b111111111;
assign micromatrizz[83][142] = 9'b111111111;
assign micromatrizz[83][143] = 9'b111111111;
assign micromatrizz[83][144] = 9'b111111111;
assign micromatrizz[83][145] = 9'b111111111;
assign micromatrizz[83][146] = 9'b111111111;
assign micromatrizz[83][147] = 9'b111111111;
assign micromatrizz[83][148] = 9'b111111111;
assign micromatrizz[83][149] = 9'b111111111;
assign micromatrizz[83][150] = 9'b111111111;
assign micromatrizz[83][151] = 9'b111111111;
assign micromatrizz[83][152] = 9'b111111111;
assign micromatrizz[83][153] = 9'b111111111;
assign micromatrizz[83][154] = 9'b111111111;
assign micromatrizz[83][155] = 9'b111111111;
assign micromatrizz[83][156] = 9'b111111111;
assign micromatrizz[83][157] = 9'b111111111;
assign micromatrizz[83][158] = 9'b111111111;
assign micromatrizz[83][159] = 9'b111111111;
assign micromatrizz[83][160] = 9'b111111111;
assign micromatrizz[83][161] = 9'b111111111;
assign micromatrizz[83][162] = 9'b111111111;
assign micromatrizz[83][163] = 9'b111111111;
assign micromatrizz[83][164] = 9'b111111111;
assign micromatrizz[83][165] = 9'b111111111;
assign micromatrizz[83][166] = 9'b111111111;
assign micromatrizz[83][167] = 9'b111111111;
assign micromatrizz[83][168] = 9'b111111111;
assign micromatrizz[83][169] = 9'b111111111;
assign micromatrizz[83][170] = 9'b111111111;
assign micromatrizz[83][171] = 9'b111111111;
assign micromatrizz[83][172] = 9'b111111111;
assign micromatrizz[83][173] = 9'b111111111;
assign micromatrizz[83][174] = 9'b111111111;
assign micromatrizz[83][175] = 9'b111111111;
assign micromatrizz[83][176] = 9'b111111111;
assign micromatrizz[83][177] = 9'b111111111;
assign micromatrizz[83][178] = 9'b111111111;
assign micromatrizz[83][179] = 9'b111111111;
assign micromatrizz[83][180] = 9'b111111111;
assign micromatrizz[83][181] = 9'b111111111;
assign micromatrizz[83][182] = 9'b111111111;
assign micromatrizz[83][183] = 9'b111111111;
assign micromatrizz[83][184] = 9'b111111111;
assign micromatrizz[83][185] = 9'b111111111;
assign micromatrizz[83][186] = 9'b111111111;
assign micromatrizz[83][187] = 9'b111111111;
assign micromatrizz[83][188] = 9'b111111111;
assign micromatrizz[83][189] = 9'b111111111;
assign micromatrizz[83][190] = 9'b111111111;
assign micromatrizz[83][191] = 9'b111111111;
assign micromatrizz[83][192] = 9'b111111111;
assign micromatrizz[83][193] = 9'b111111111;
assign micromatrizz[83][194] = 9'b111111111;
assign micromatrizz[83][195] = 9'b111111111;
assign micromatrizz[83][196] = 9'b111111111;
assign micromatrizz[83][197] = 9'b111111111;
assign micromatrizz[83][198] = 9'b111111111;
assign micromatrizz[83][199] = 9'b111111111;
assign micromatrizz[83][200] = 9'b111111111;
assign micromatrizz[83][201] = 9'b111111111;
assign micromatrizz[83][202] = 9'b111111111;
assign micromatrizz[83][203] = 9'b111111111;
assign micromatrizz[83][204] = 9'b111111111;
assign micromatrizz[83][205] = 9'b111111111;
assign micromatrizz[83][206] = 9'b111111111;
assign micromatrizz[83][207] = 9'b111111111;
assign micromatrizz[83][208] = 9'b111111111;
assign micromatrizz[83][209] = 9'b111111111;
assign micromatrizz[83][210] = 9'b111111111;
assign micromatrizz[83][211] = 9'b111111111;
assign micromatrizz[83][212] = 9'b111111111;
assign micromatrizz[83][213] = 9'b111111111;
assign micromatrizz[83][214] = 9'b111111111;
assign micromatrizz[83][215] = 9'b111111111;
assign micromatrizz[83][216] = 9'b111111111;
assign micromatrizz[83][217] = 9'b111111111;
assign micromatrizz[83][218] = 9'b111111111;
assign micromatrizz[83][219] = 9'b111111111;
assign micromatrizz[83][220] = 9'b111111111;
assign micromatrizz[83][221] = 9'b111111111;
assign micromatrizz[83][222] = 9'b111111111;
assign micromatrizz[83][223] = 9'b111111111;
assign micromatrizz[83][224] = 9'b111111111;
assign micromatrizz[83][225] = 9'b111111111;
assign micromatrizz[83][226] = 9'b111111111;
assign micromatrizz[83][227] = 9'b111111111;
assign micromatrizz[83][228] = 9'b111111111;
assign micromatrizz[83][229] = 9'b111111111;
assign micromatrizz[83][230] = 9'b111111111;
assign micromatrizz[83][231] = 9'b111111111;
assign micromatrizz[83][232] = 9'b111111111;
assign micromatrizz[83][233] = 9'b111111111;
assign micromatrizz[83][234] = 9'b111111111;
assign micromatrizz[83][235] = 9'b111111111;
assign micromatrizz[83][236] = 9'b111111111;
assign micromatrizz[83][237] = 9'b111111111;
assign micromatrizz[83][238] = 9'b111111111;
assign micromatrizz[83][239] = 9'b111111111;
assign micromatrizz[83][240] = 9'b111111111;
assign micromatrizz[83][241] = 9'b111111111;
assign micromatrizz[83][242] = 9'b111111111;
assign micromatrizz[83][243] = 9'b111111111;
assign micromatrizz[83][244] = 9'b111111111;
assign micromatrizz[83][245] = 9'b111111111;
assign micromatrizz[83][246] = 9'b111111111;
assign micromatrizz[83][247] = 9'b111111111;
assign micromatrizz[83][248] = 9'b111111111;
assign micromatrizz[83][249] = 9'b111111111;
assign micromatrizz[83][250] = 9'b111111111;
assign micromatrizz[83][251] = 9'b111111111;
assign micromatrizz[83][252] = 9'b111111111;
assign micromatrizz[83][253] = 9'b111111111;
assign micromatrizz[83][254] = 9'b111111111;
assign micromatrizz[83][255] = 9'b111111111;
assign micromatrizz[83][256] = 9'b111111111;
assign micromatrizz[83][257] = 9'b111111111;
assign micromatrizz[83][258] = 9'b111111111;
assign micromatrizz[83][259] = 9'b111111111;
assign micromatrizz[83][260] = 9'b111111111;
assign micromatrizz[83][261] = 9'b111111111;
assign micromatrizz[83][262] = 9'b111111111;
assign micromatrizz[83][263] = 9'b111111111;
assign micromatrizz[83][264] = 9'b111111111;
assign micromatrizz[83][265] = 9'b111111111;
assign micromatrizz[83][266] = 9'b111111111;
assign micromatrizz[83][267] = 9'b111111111;
assign micromatrizz[83][268] = 9'b111111111;
assign micromatrizz[83][269] = 9'b111111111;
assign micromatrizz[83][270] = 9'b111111111;
assign micromatrizz[83][271] = 9'b111111111;
assign micromatrizz[83][272] = 9'b111111111;
assign micromatrizz[83][273] = 9'b111111111;
assign micromatrizz[83][274] = 9'b111111111;
assign micromatrizz[83][275] = 9'b111111111;
assign micromatrizz[83][276] = 9'b111111111;
assign micromatrizz[83][277] = 9'b111111111;
assign micromatrizz[83][278] = 9'b111111111;
assign micromatrizz[83][279] = 9'b111111111;
assign micromatrizz[83][280] = 9'b111111111;
assign micromatrizz[83][281] = 9'b111111111;
assign micromatrizz[83][282] = 9'b111111111;
assign micromatrizz[83][283] = 9'b111111111;
assign micromatrizz[83][284] = 9'b111111111;
assign micromatrizz[83][285] = 9'b111111111;
assign micromatrizz[83][286] = 9'b111111111;
assign micromatrizz[83][287] = 9'b111111111;
assign micromatrizz[83][288] = 9'b111111111;
assign micromatrizz[83][289] = 9'b111111111;
assign micromatrizz[83][290] = 9'b111111111;
assign micromatrizz[83][291] = 9'b111111111;
assign micromatrizz[83][292] = 9'b111111111;
assign micromatrizz[83][293] = 9'b111111111;
assign micromatrizz[83][294] = 9'b111111111;
assign micromatrizz[83][295] = 9'b111111111;
assign micromatrizz[83][296] = 9'b111111111;
assign micromatrizz[83][297] = 9'b111111111;
assign micromatrizz[83][298] = 9'b111111111;
assign micromatrizz[83][299] = 9'b111111111;
assign micromatrizz[83][300] = 9'b111111111;
assign micromatrizz[83][301] = 9'b111111111;
assign micromatrizz[83][302] = 9'b111111111;
assign micromatrizz[83][303] = 9'b111111111;
assign micromatrizz[83][304] = 9'b111111111;
assign micromatrizz[83][305] = 9'b111111111;
assign micromatrizz[83][306] = 9'b111111111;
assign micromatrizz[83][307] = 9'b111111111;
assign micromatrizz[83][308] = 9'b111111111;
assign micromatrizz[83][309] = 9'b111111111;
assign micromatrizz[83][310] = 9'b111111111;
assign micromatrizz[83][311] = 9'b111111111;
assign micromatrizz[83][312] = 9'b111111111;
assign micromatrizz[83][313] = 9'b111111111;
assign micromatrizz[83][314] = 9'b111111111;
assign micromatrizz[83][315] = 9'b111111111;
assign micromatrizz[83][316] = 9'b111111111;
assign micromatrizz[83][317] = 9'b111111111;
assign micromatrizz[83][318] = 9'b111111111;
assign micromatrizz[83][319] = 9'b111111111;
assign micromatrizz[83][320] = 9'b111111111;
assign micromatrizz[83][321] = 9'b111111111;
assign micromatrizz[83][322] = 9'b111111111;
assign micromatrizz[83][323] = 9'b111111111;
assign micromatrizz[83][324] = 9'b111111111;
assign micromatrizz[83][325] = 9'b111111111;
assign micromatrizz[83][326] = 9'b111111111;
assign micromatrizz[83][327] = 9'b111111111;
assign micromatrizz[83][328] = 9'b111111111;
assign micromatrizz[83][329] = 9'b111111111;
assign micromatrizz[83][330] = 9'b111111111;
assign micromatrizz[83][331] = 9'b111111111;
assign micromatrizz[83][332] = 9'b111111111;
assign micromatrizz[83][333] = 9'b111111111;
assign micromatrizz[83][334] = 9'b111111111;
assign micromatrizz[83][335] = 9'b111111111;
assign micromatrizz[83][336] = 9'b111111111;
assign micromatrizz[83][337] = 9'b111111111;
assign micromatrizz[83][338] = 9'b111111111;
assign micromatrizz[83][339] = 9'b111111111;
assign micromatrizz[83][340] = 9'b111111111;
assign micromatrizz[83][341] = 9'b111111111;
assign micromatrizz[83][342] = 9'b111111111;
assign micromatrizz[83][343] = 9'b111111111;
assign micromatrizz[83][344] = 9'b111111111;
assign micromatrizz[83][345] = 9'b111111111;
assign micromatrizz[83][346] = 9'b111111111;
assign micromatrizz[83][347] = 9'b111111111;
assign micromatrizz[83][348] = 9'b111111111;
assign micromatrizz[83][349] = 9'b111111111;
assign micromatrizz[83][350] = 9'b111111111;
assign micromatrizz[83][351] = 9'b111111111;
assign micromatrizz[83][352] = 9'b111111111;
assign micromatrizz[83][353] = 9'b111111111;
assign micromatrizz[83][354] = 9'b111111111;
assign micromatrizz[83][355] = 9'b111111111;
assign micromatrizz[83][356] = 9'b111111111;
assign micromatrizz[83][357] = 9'b111111111;
assign micromatrizz[83][358] = 9'b111111111;
assign micromatrizz[83][359] = 9'b111111111;
assign micromatrizz[83][360] = 9'b111111111;
assign micromatrizz[83][361] = 9'b111111111;
assign micromatrizz[83][362] = 9'b111111111;
assign micromatrizz[83][363] = 9'b111111111;
assign micromatrizz[83][364] = 9'b111111111;
assign micromatrizz[83][365] = 9'b111111111;
assign micromatrizz[83][366] = 9'b111111111;
assign micromatrizz[83][367] = 9'b111111111;
assign micromatrizz[83][368] = 9'b111111111;
assign micromatrizz[83][369] = 9'b111111111;
assign micromatrizz[83][370] = 9'b111111111;
assign micromatrizz[83][371] = 9'b111111111;
assign micromatrizz[83][372] = 9'b111111111;
assign micromatrizz[83][373] = 9'b111111111;
assign micromatrizz[83][374] = 9'b111111111;
assign micromatrizz[83][375] = 9'b111111111;
assign micromatrizz[83][376] = 9'b111111111;
assign micromatrizz[83][377] = 9'b111111111;
assign micromatrizz[83][378] = 9'b111111111;
assign micromatrizz[83][379] = 9'b111111111;
assign micromatrizz[83][380] = 9'b111111111;
assign micromatrizz[83][381] = 9'b111111111;
assign micromatrizz[83][382] = 9'b111111111;
assign micromatrizz[83][383] = 9'b111111111;
assign micromatrizz[83][384] = 9'b111111111;
assign micromatrizz[83][385] = 9'b111111111;
assign micromatrizz[83][386] = 9'b111111111;
assign micromatrizz[83][387] = 9'b111111111;
assign micromatrizz[83][388] = 9'b111111111;
assign micromatrizz[83][389] = 9'b111111111;
assign micromatrizz[83][390] = 9'b111111111;
assign micromatrizz[83][391] = 9'b111111111;
assign micromatrizz[83][392] = 9'b111111111;
assign micromatrizz[83][393] = 9'b111111111;
assign micromatrizz[83][394] = 9'b111111111;
assign micromatrizz[83][395] = 9'b111111111;
assign micromatrizz[83][396] = 9'b111111111;
assign micromatrizz[83][397] = 9'b111111111;
assign micromatrizz[83][398] = 9'b111111111;
assign micromatrizz[83][399] = 9'b111111111;
assign micromatrizz[83][400] = 9'b111111111;
assign micromatrizz[83][401] = 9'b111111111;
assign micromatrizz[83][402] = 9'b111111111;
assign micromatrizz[83][403] = 9'b111111111;
assign micromatrizz[83][404] = 9'b111111111;
assign micromatrizz[83][405] = 9'b111111111;
assign micromatrizz[83][406] = 9'b111111111;
assign micromatrizz[83][407] = 9'b111111111;
assign micromatrizz[83][408] = 9'b111111111;
assign micromatrizz[83][409] = 9'b111111111;
assign micromatrizz[83][410] = 9'b111111111;
assign micromatrizz[83][411] = 9'b111111111;
assign micromatrizz[83][412] = 9'b111111111;
assign micromatrizz[83][413] = 9'b111111111;
assign micromatrizz[83][414] = 9'b111111111;
assign micromatrizz[83][415] = 9'b111111111;
assign micromatrizz[83][416] = 9'b111111111;
assign micromatrizz[83][417] = 9'b111111111;
assign micromatrizz[83][418] = 9'b111111111;
assign micromatrizz[83][419] = 9'b111111111;
assign micromatrizz[83][420] = 9'b111111111;
assign micromatrizz[83][421] = 9'b111111111;
assign micromatrizz[83][422] = 9'b111111111;
assign micromatrizz[83][423] = 9'b111111111;
assign micromatrizz[83][424] = 9'b111111111;
assign micromatrizz[83][425] = 9'b111111111;
assign micromatrizz[83][426] = 9'b111111111;
assign micromatrizz[83][427] = 9'b111111111;
assign micromatrizz[83][428] = 9'b111111111;
assign micromatrizz[83][429] = 9'b111111111;
assign micromatrizz[83][430] = 9'b111111111;
assign micromatrizz[83][431] = 9'b111111111;
assign micromatrizz[83][432] = 9'b111111111;
assign micromatrizz[83][433] = 9'b111111111;
assign micromatrizz[83][434] = 9'b111111111;
assign micromatrizz[83][435] = 9'b111111111;
assign micromatrizz[83][436] = 9'b111111111;
assign micromatrizz[83][437] = 9'b111111111;
assign micromatrizz[83][438] = 9'b111111111;
assign micromatrizz[83][439] = 9'b111111111;
assign micromatrizz[83][440] = 9'b111111111;
assign micromatrizz[83][441] = 9'b111111111;
assign micromatrizz[83][442] = 9'b111111111;
assign micromatrizz[83][443] = 9'b111111111;
assign micromatrizz[83][444] = 9'b111111111;
assign micromatrizz[83][445] = 9'b111111111;
assign micromatrizz[83][446] = 9'b111111111;
assign micromatrizz[83][447] = 9'b111111111;
assign micromatrizz[83][448] = 9'b111111111;
assign micromatrizz[83][449] = 9'b111111111;
assign micromatrizz[83][450] = 9'b111111111;
assign micromatrizz[83][451] = 9'b111111111;
assign micromatrizz[83][452] = 9'b111111111;
assign micromatrizz[83][453] = 9'b111111111;
assign micromatrizz[83][454] = 9'b111111111;
assign micromatrizz[83][455] = 9'b111111111;
assign micromatrizz[83][456] = 9'b111111111;
assign micromatrizz[83][457] = 9'b111111111;
assign micromatrizz[83][458] = 9'b111111111;
assign micromatrizz[83][459] = 9'b111111111;
assign micromatrizz[83][460] = 9'b111111111;
assign micromatrizz[83][461] = 9'b111111111;
assign micromatrizz[83][462] = 9'b111111111;
assign micromatrizz[83][463] = 9'b111111111;
assign micromatrizz[83][464] = 9'b111111111;
assign micromatrizz[83][465] = 9'b111111111;
assign micromatrizz[83][466] = 9'b111111111;
assign micromatrizz[83][467] = 9'b111111111;
assign micromatrizz[83][468] = 9'b111111111;
assign micromatrizz[83][469] = 9'b111111111;
assign micromatrizz[83][470] = 9'b111111111;
assign micromatrizz[83][471] = 9'b111111111;
assign micromatrizz[83][472] = 9'b111111111;
assign micromatrizz[83][473] = 9'b111111111;
assign micromatrizz[83][474] = 9'b111111111;
assign micromatrizz[83][475] = 9'b111111111;
assign micromatrizz[83][476] = 9'b111111111;
assign micromatrizz[83][477] = 9'b111111111;
assign micromatrizz[83][478] = 9'b111111111;
assign micromatrizz[83][479] = 9'b111111111;
assign micromatrizz[83][480] = 9'b111111111;
assign micromatrizz[83][481] = 9'b111111111;
assign micromatrizz[83][482] = 9'b111111111;
assign micromatrizz[83][483] = 9'b111111111;
assign micromatrizz[83][484] = 9'b111111111;
assign micromatrizz[83][485] = 9'b111111111;
assign micromatrizz[83][486] = 9'b111111111;
assign micromatrizz[83][487] = 9'b111111111;
assign micromatrizz[83][488] = 9'b111111111;
assign micromatrizz[83][489] = 9'b111111111;
assign micromatrizz[83][490] = 9'b111111111;
assign micromatrizz[83][491] = 9'b111111111;
assign micromatrizz[83][492] = 9'b111111111;
assign micromatrizz[83][493] = 9'b111111111;
assign micromatrizz[83][494] = 9'b111111111;
assign micromatrizz[83][495] = 9'b111111111;
assign micromatrizz[83][496] = 9'b111111111;
assign micromatrizz[83][497] = 9'b111111111;
assign micromatrizz[83][498] = 9'b111111111;
assign micromatrizz[83][499] = 9'b111111111;
assign micromatrizz[83][500] = 9'b111111111;
assign micromatrizz[83][501] = 9'b111111111;
assign micromatrizz[83][502] = 9'b111111111;
assign micromatrizz[83][503] = 9'b111111111;
assign micromatrizz[83][504] = 9'b111111111;
assign micromatrizz[83][505] = 9'b111111111;
assign micromatrizz[83][506] = 9'b111111111;
assign micromatrizz[83][507] = 9'b111111111;
assign micromatrizz[83][508] = 9'b111111111;
assign micromatrizz[83][509] = 9'b111111111;
assign micromatrizz[83][510] = 9'b111111111;
assign micromatrizz[83][511] = 9'b111111111;
assign micromatrizz[83][512] = 9'b111111111;
assign micromatrizz[83][513] = 9'b111111111;
assign micromatrizz[83][514] = 9'b111111111;
assign micromatrizz[83][515] = 9'b111111111;
assign micromatrizz[83][516] = 9'b111111111;
assign micromatrizz[83][517] = 9'b111111111;
assign micromatrizz[83][518] = 9'b111111111;
assign micromatrizz[83][519] = 9'b111111111;
assign micromatrizz[83][520] = 9'b111111111;
assign micromatrizz[83][521] = 9'b111111111;
assign micromatrizz[83][522] = 9'b111111111;
assign micromatrizz[83][523] = 9'b111111111;
assign micromatrizz[83][524] = 9'b111111111;
assign micromatrizz[83][525] = 9'b111111111;
assign micromatrizz[83][526] = 9'b111111111;
assign micromatrizz[83][527] = 9'b111111111;
assign micromatrizz[83][528] = 9'b111111111;
assign micromatrizz[83][529] = 9'b111111111;
assign micromatrizz[83][530] = 9'b111111111;
assign micromatrizz[83][531] = 9'b111111111;
assign micromatrizz[83][532] = 9'b111111111;
assign micromatrizz[83][533] = 9'b111111111;
assign micromatrizz[83][534] = 9'b111111111;
assign micromatrizz[83][535] = 9'b111111111;
assign micromatrizz[83][536] = 9'b111111111;
assign micromatrizz[83][537] = 9'b111111111;
assign micromatrizz[83][538] = 9'b111111111;
assign micromatrizz[83][539] = 9'b111111111;
assign micromatrizz[83][540] = 9'b111111111;
assign micromatrizz[83][541] = 9'b111111111;
assign micromatrizz[83][542] = 9'b111111111;
assign micromatrizz[83][543] = 9'b111111111;
assign micromatrizz[83][544] = 9'b111111111;
assign micromatrizz[83][545] = 9'b111111111;
assign micromatrizz[83][546] = 9'b111111111;
assign micromatrizz[83][547] = 9'b111111111;
assign micromatrizz[83][548] = 9'b111111111;
assign micromatrizz[83][549] = 9'b111111111;
assign micromatrizz[83][550] = 9'b111111111;
assign micromatrizz[83][551] = 9'b111111111;
assign micromatrizz[83][552] = 9'b111111111;
assign micromatrizz[83][553] = 9'b111111111;
assign micromatrizz[83][554] = 9'b111111111;
assign micromatrizz[83][555] = 9'b111111111;
assign micromatrizz[83][556] = 9'b111111111;
assign micromatrizz[83][557] = 9'b111111111;
assign micromatrizz[83][558] = 9'b111111111;
assign micromatrizz[83][559] = 9'b111111111;
assign micromatrizz[83][560] = 9'b111111111;
assign micromatrizz[83][561] = 9'b111111111;
assign micromatrizz[83][562] = 9'b111111111;
assign micromatrizz[83][563] = 9'b111111111;
assign micromatrizz[83][564] = 9'b111111111;
assign micromatrizz[83][565] = 9'b111111111;
assign micromatrizz[83][566] = 9'b111111111;
assign micromatrizz[83][567] = 9'b111111111;
assign micromatrizz[83][568] = 9'b111111111;
assign micromatrizz[83][569] = 9'b111111111;
assign micromatrizz[83][570] = 9'b111111111;
assign micromatrizz[83][571] = 9'b111111111;
assign micromatrizz[83][572] = 9'b111111111;
assign micromatrizz[83][573] = 9'b111111111;
assign micromatrizz[83][574] = 9'b111111111;
assign micromatrizz[83][575] = 9'b111111111;
assign micromatrizz[83][576] = 9'b111111111;
assign micromatrizz[83][577] = 9'b111111111;
assign micromatrizz[83][578] = 9'b111111111;
assign micromatrizz[83][579] = 9'b111111111;
assign micromatrizz[83][580] = 9'b111111111;
assign micromatrizz[83][581] = 9'b111111111;
assign micromatrizz[83][582] = 9'b111111111;
assign micromatrizz[83][583] = 9'b111111111;
assign micromatrizz[83][584] = 9'b111111111;
assign micromatrizz[83][585] = 9'b111111111;
assign micromatrizz[83][586] = 9'b111111111;
assign micromatrizz[83][587] = 9'b111111111;
assign micromatrizz[83][588] = 9'b111111111;
assign micromatrizz[83][589] = 9'b111111111;
assign micromatrizz[83][590] = 9'b111111111;
assign micromatrizz[83][591] = 9'b111111111;
assign micromatrizz[83][592] = 9'b111111111;
assign micromatrizz[83][593] = 9'b111111111;
assign micromatrizz[83][594] = 9'b111111111;
assign micromatrizz[83][595] = 9'b111111111;
assign micromatrizz[83][596] = 9'b111111111;
assign micromatrizz[83][597] = 9'b111111111;
assign micromatrizz[83][598] = 9'b111111111;
assign micromatrizz[83][599] = 9'b111111111;
assign micromatrizz[83][600] = 9'b111111111;
assign micromatrizz[83][601] = 9'b111111111;
assign micromatrizz[83][602] = 9'b111111111;
assign micromatrizz[83][603] = 9'b111111111;
assign micromatrizz[83][604] = 9'b111111111;
assign micromatrizz[83][605] = 9'b111111111;
assign micromatrizz[83][606] = 9'b111111111;
assign micromatrizz[83][607] = 9'b111111111;
assign micromatrizz[83][608] = 9'b111111111;
assign micromatrizz[83][609] = 9'b111111111;
assign micromatrizz[83][610] = 9'b111111111;
assign micromatrizz[83][611] = 9'b111111111;
assign micromatrizz[83][612] = 9'b111111111;
assign micromatrizz[83][613] = 9'b111111111;
assign micromatrizz[83][614] = 9'b111111111;
assign micromatrizz[83][615] = 9'b111111111;
assign micromatrizz[83][616] = 9'b111111111;
assign micromatrizz[83][617] = 9'b111111111;
assign micromatrizz[83][618] = 9'b111111111;
assign micromatrizz[83][619] = 9'b111111111;
assign micromatrizz[83][620] = 9'b111111111;
assign micromatrizz[83][621] = 9'b111111111;
assign micromatrizz[83][622] = 9'b111111111;
assign micromatrizz[83][623] = 9'b111111111;
assign micromatrizz[83][624] = 9'b111111111;
assign micromatrizz[83][625] = 9'b111111111;
assign micromatrizz[83][626] = 9'b111111111;
assign micromatrizz[83][627] = 9'b111111111;
assign micromatrizz[83][628] = 9'b111111111;
assign micromatrizz[83][629] = 9'b111111111;
assign micromatrizz[83][630] = 9'b111111111;
assign micromatrizz[83][631] = 9'b111111111;
assign micromatrizz[83][632] = 9'b111111111;
assign micromatrizz[83][633] = 9'b111111111;
assign micromatrizz[83][634] = 9'b111111111;
assign micromatrizz[83][635] = 9'b111111111;
assign micromatrizz[83][636] = 9'b111111111;
assign micromatrizz[83][637] = 9'b111111111;
assign micromatrizz[83][638] = 9'b111111111;
assign micromatrizz[83][639] = 9'b111111111;
assign micromatrizz[84][0] = 9'b111111111;
assign micromatrizz[84][1] = 9'b111111111;
assign micromatrizz[84][2] = 9'b111111111;
assign micromatrizz[84][3] = 9'b111111111;
assign micromatrizz[84][4] = 9'b111111111;
assign micromatrizz[84][5] = 9'b111111111;
assign micromatrizz[84][6] = 9'b111111111;
assign micromatrizz[84][7] = 9'b111111111;
assign micromatrizz[84][8] = 9'b111111111;
assign micromatrizz[84][9] = 9'b111111111;
assign micromatrizz[84][10] = 9'b111111111;
assign micromatrizz[84][11] = 9'b111111111;
assign micromatrizz[84][12] = 9'b111111111;
assign micromatrizz[84][13] = 9'b111111111;
assign micromatrizz[84][14] = 9'b111111111;
assign micromatrizz[84][15] = 9'b111111111;
assign micromatrizz[84][16] = 9'b111111111;
assign micromatrizz[84][17] = 9'b111111111;
assign micromatrizz[84][18] = 9'b111111111;
assign micromatrizz[84][19] = 9'b111111111;
assign micromatrizz[84][20] = 9'b111111111;
assign micromatrizz[84][21] = 9'b111111111;
assign micromatrizz[84][22] = 9'b111111111;
assign micromatrizz[84][23] = 9'b111111111;
assign micromatrizz[84][24] = 9'b111111111;
assign micromatrizz[84][25] = 9'b111111111;
assign micromatrizz[84][26] = 9'b111111111;
assign micromatrizz[84][27] = 9'b111111111;
assign micromatrizz[84][28] = 9'b111111111;
assign micromatrizz[84][29] = 9'b111111111;
assign micromatrizz[84][30] = 9'b111111111;
assign micromatrizz[84][31] = 9'b111111111;
assign micromatrizz[84][32] = 9'b111111111;
assign micromatrizz[84][33] = 9'b111111111;
assign micromatrizz[84][34] = 9'b111111111;
assign micromatrizz[84][35] = 9'b111111111;
assign micromatrizz[84][36] = 9'b111111111;
assign micromatrizz[84][37] = 9'b111111111;
assign micromatrizz[84][38] = 9'b111111111;
assign micromatrizz[84][39] = 9'b111111111;
assign micromatrizz[84][40] = 9'b111111111;
assign micromatrizz[84][41] = 9'b111111111;
assign micromatrizz[84][42] = 9'b111111111;
assign micromatrizz[84][43] = 9'b111111111;
assign micromatrizz[84][44] = 9'b111111111;
assign micromatrizz[84][45] = 9'b111111111;
assign micromatrizz[84][46] = 9'b111111111;
assign micromatrizz[84][47] = 9'b111111111;
assign micromatrizz[84][48] = 9'b111111111;
assign micromatrizz[84][49] = 9'b111111111;
assign micromatrizz[84][50] = 9'b111111111;
assign micromatrizz[84][51] = 9'b111111111;
assign micromatrizz[84][52] = 9'b111111111;
assign micromatrizz[84][53] = 9'b111111111;
assign micromatrizz[84][54] = 9'b111111111;
assign micromatrizz[84][55] = 9'b111111111;
assign micromatrizz[84][56] = 9'b111111111;
assign micromatrizz[84][57] = 9'b111111111;
assign micromatrizz[84][58] = 9'b111111111;
assign micromatrizz[84][59] = 9'b111111111;
assign micromatrizz[84][60] = 9'b111111111;
assign micromatrizz[84][61] = 9'b111111111;
assign micromatrizz[84][62] = 9'b111111111;
assign micromatrizz[84][63] = 9'b111111111;
assign micromatrizz[84][64] = 9'b111111111;
assign micromatrizz[84][65] = 9'b111111111;
assign micromatrizz[84][66] = 9'b111111111;
assign micromatrizz[84][67] = 9'b111111111;
assign micromatrizz[84][68] = 9'b111111111;
assign micromatrizz[84][69] = 9'b111111111;
assign micromatrizz[84][70] = 9'b111111111;
assign micromatrizz[84][71] = 9'b111111111;
assign micromatrizz[84][72] = 9'b111111111;
assign micromatrizz[84][73] = 9'b111111111;
assign micromatrizz[84][74] = 9'b111111111;
assign micromatrizz[84][75] = 9'b111111111;
assign micromatrizz[84][76] = 9'b111111111;
assign micromatrizz[84][77] = 9'b111111111;
assign micromatrizz[84][78] = 9'b111111111;
assign micromatrizz[84][79] = 9'b111111111;
assign micromatrizz[84][80] = 9'b111111111;
assign micromatrizz[84][81] = 9'b111111111;
assign micromatrizz[84][82] = 9'b111111111;
assign micromatrizz[84][83] = 9'b111111111;
assign micromatrizz[84][84] = 9'b111111111;
assign micromatrizz[84][85] = 9'b111111111;
assign micromatrizz[84][86] = 9'b111111111;
assign micromatrizz[84][87] = 9'b111111111;
assign micromatrizz[84][88] = 9'b111111111;
assign micromatrizz[84][89] = 9'b111111111;
assign micromatrizz[84][90] = 9'b111111111;
assign micromatrizz[84][91] = 9'b111111111;
assign micromatrizz[84][92] = 9'b111111111;
assign micromatrizz[84][93] = 9'b111111111;
assign micromatrizz[84][94] = 9'b111111111;
assign micromatrizz[84][95] = 9'b111111111;
assign micromatrizz[84][96] = 9'b111111111;
assign micromatrizz[84][97] = 9'b111111111;
assign micromatrizz[84][98] = 9'b111111111;
assign micromatrizz[84][99] = 9'b111111111;
assign micromatrizz[84][100] = 9'b111111111;
assign micromatrizz[84][101] = 9'b111111111;
assign micromatrizz[84][102] = 9'b111111111;
assign micromatrizz[84][103] = 9'b111111111;
assign micromatrizz[84][104] = 9'b111111111;
assign micromatrizz[84][105] = 9'b111111111;
assign micromatrizz[84][106] = 9'b111111111;
assign micromatrizz[84][107] = 9'b111111111;
assign micromatrizz[84][108] = 9'b111111111;
assign micromatrizz[84][109] = 9'b111111111;
assign micromatrizz[84][110] = 9'b111111111;
assign micromatrizz[84][111] = 9'b111111111;
assign micromatrizz[84][112] = 9'b111111111;
assign micromatrizz[84][113] = 9'b111111111;
assign micromatrizz[84][114] = 9'b111111111;
assign micromatrizz[84][115] = 9'b111111111;
assign micromatrizz[84][116] = 9'b111111111;
assign micromatrizz[84][117] = 9'b111111111;
assign micromatrizz[84][118] = 9'b111111111;
assign micromatrizz[84][119] = 9'b111111111;
assign micromatrizz[84][120] = 9'b111111111;
assign micromatrizz[84][121] = 9'b111111111;
assign micromatrizz[84][122] = 9'b111111111;
assign micromatrizz[84][123] = 9'b111111111;
assign micromatrizz[84][124] = 9'b111111111;
assign micromatrizz[84][125] = 9'b111111111;
assign micromatrizz[84][126] = 9'b111111111;
assign micromatrizz[84][127] = 9'b111111111;
assign micromatrizz[84][128] = 9'b111111111;
assign micromatrizz[84][129] = 9'b111111111;
assign micromatrizz[84][130] = 9'b111111111;
assign micromatrizz[84][131] = 9'b111111111;
assign micromatrizz[84][132] = 9'b111111111;
assign micromatrizz[84][133] = 9'b111111111;
assign micromatrizz[84][134] = 9'b111111111;
assign micromatrizz[84][135] = 9'b111111111;
assign micromatrizz[84][136] = 9'b111111111;
assign micromatrizz[84][137] = 9'b111111111;
assign micromatrizz[84][138] = 9'b111111111;
assign micromatrizz[84][139] = 9'b111111111;
assign micromatrizz[84][140] = 9'b111111111;
assign micromatrizz[84][141] = 9'b111111111;
assign micromatrizz[84][142] = 9'b111111111;
assign micromatrizz[84][143] = 9'b111111111;
assign micromatrizz[84][144] = 9'b111111111;
assign micromatrizz[84][145] = 9'b111111111;
assign micromatrizz[84][146] = 9'b111111111;
assign micromatrizz[84][147] = 9'b111111111;
assign micromatrizz[84][148] = 9'b111111111;
assign micromatrizz[84][149] = 9'b111111111;
assign micromatrizz[84][150] = 9'b111111111;
assign micromatrizz[84][151] = 9'b111111111;
assign micromatrizz[84][152] = 9'b111111111;
assign micromatrizz[84][153] = 9'b111111111;
assign micromatrizz[84][154] = 9'b111111111;
assign micromatrizz[84][155] = 9'b111111111;
assign micromatrizz[84][156] = 9'b111111111;
assign micromatrizz[84][157] = 9'b111111111;
assign micromatrizz[84][158] = 9'b111111111;
assign micromatrizz[84][159] = 9'b111111111;
assign micromatrizz[84][160] = 9'b111111111;
assign micromatrizz[84][161] = 9'b111111111;
assign micromatrizz[84][162] = 9'b111111111;
assign micromatrizz[84][163] = 9'b111111111;
assign micromatrizz[84][164] = 9'b111111111;
assign micromatrizz[84][165] = 9'b111111111;
assign micromatrizz[84][166] = 9'b111111111;
assign micromatrizz[84][167] = 9'b111111111;
assign micromatrizz[84][168] = 9'b111111111;
assign micromatrizz[84][169] = 9'b111111111;
assign micromatrizz[84][170] = 9'b111111111;
assign micromatrizz[84][171] = 9'b111111111;
assign micromatrizz[84][172] = 9'b111111111;
assign micromatrizz[84][173] = 9'b111111111;
assign micromatrizz[84][174] = 9'b111111111;
assign micromatrizz[84][175] = 9'b111111111;
assign micromatrizz[84][176] = 9'b111111111;
assign micromatrizz[84][177] = 9'b111111111;
assign micromatrizz[84][178] = 9'b111111111;
assign micromatrizz[84][179] = 9'b111111111;
assign micromatrizz[84][180] = 9'b111111111;
assign micromatrizz[84][181] = 9'b111111111;
assign micromatrizz[84][182] = 9'b111111111;
assign micromatrizz[84][183] = 9'b111111111;
assign micromatrizz[84][184] = 9'b111111111;
assign micromatrizz[84][185] = 9'b111111111;
assign micromatrizz[84][186] = 9'b111111111;
assign micromatrizz[84][187] = 9'b111111111;
assign micromatrizz[84][188] = 9'b111111111;
assign micromatrizz[84][189] = 9'b111111111;
assign micromatrizz[84][190] = 9'b111111111;
assign micromatrizz[84][191] = 9'b111111111;
assign micromatrizz[84][192] = 9'b111111111;
assign micromatrizz[84][193] = 9'b111111111;
assign micromatrizz[84][194] = 9'b111111111;
assign micromatrizz[84][195] = 9'b111111111;
assign micromatrizz[84][196] = 9'b111111111;
assign micromatrizz[84][197] = 9'b111111111;
assign micromatrizz[84][198] = 9'b111111111;
assign micromatrizz[84][199] = 9'b111111111;
assign micromatrizz[84][200] = 9'b111111111;
assign micromatrizz[84][201] = 9'b111111111;
assign micromatrizz[84][202] = 9'b111111111;
assign micromatrizz[84][203] = 9'b111111111;
assign micromatrizz[84][204] = 9'b111111111;
assign micromatrizz[84][205] = 9'b111111111;
assign micromatrizz[84][206] = 9'b111111111;
assign micromatrizz[84][207] = 9'b111111111;
assign micromatrizz[84][208] = 9'b111111111;
assign micromatrizz[84][209] = 9'b111111111;
assign micromatrizz[84][210] = 9'b111111111;
assign micromatrizz[84][211] = 9'b111111111;
assign micromatrizz[84][212] = 9'b111111111;
assign micromatrizz[84][213] = 9'b111111111;
assign micromatrizz[84][214] = 9'b111111111;
assign micromatrizz[84][215] = 9'b111111111;
assign micromatrizz[84][216] = 9'b111111111;
assign micromatrizz[84][217] = 9'b111111111;
assign micromatrizz[84][218] = 9'b111111111;
assign micromatrizz[84][219] = 9'b111111111;
assign micromatrizz[84][220] = 9'b111111111;
assign micromatrizz[84][221] = 9'b111111111;
assign micromatrizz[84][222] = 9'b111111111;
assign micromatrizz[84][223] = 9'b111111111;
assign micromatrizz[84][224] = 9'b111111111;
assign micromatrizz[84][225] = 9'b111111111;
assign micromatrizz[84][226] = 9'b111111111;
assign micromatrizz[84][227] = 9'b111111111;
assign micromatrizz[84][228] = 9'b111111111;
assign micromatrizz[84][229] = 9'b111111111;
assign micromatrizz[84][230] = 9'b111111111;
assign micromatrizz[84][231] = 9'b111111111;
assign micromatrizz[84][232] = 9'b111111111;
assign micromatrizz[84][233] = 9'b111111111;
assign micromatrizz[84][234] = 9'b111111111;
assign micromatrizz[84][235] = 9'b111111111;
assign micromatrizz[84][236] = 9'b111111111;
assign micromatrizz[84][237] = 9'b111111111;
assign micromatrizz[84][238] = 9'b111111111;
assign micromatrizz[84][239] = 9'b111111111;
assign micromatrizz[84][240] = 9'b111111111;
assign micromatrizz[84][241] = 9'b111111111;
assign micromatrizz[84][242] = 9'b111111111;
assign micromatrizz[84][243] = 9'b111111111;
assign micromatrizz[84][244] = 9'b111111111;
assign micromatrizz[84][245] = 9'b111111111;
assign micromatrizz[84][246] = 9'b111111111;
assign micromatrizz[84][247] = 9'b111111111;
assign micromatrizz[84][248] = 9'b111111111;
assign micromatrizz[84][249] = 9'b111111111;
assign micromatrizz[84][250] = 9'b111111111;
assign micromatrizz[84][251] = 9'b111111111;
assign micromatrizz[84][252] = 9'b111111111;
assign micromatrizz[84][253] = 9'b111111111;
assign micromatrizz[84][254] = 9'b111111111;
assign micromatrizz[84][255] = 9'b111111111;
assign micromatrizz[84][256] = 9'b111111111;
assign micromatrizz[84][257] = 9'b111111111;
assign micromatrizz[84][258] = 9'b111111111;
assign micromatrizz[84][259] = 9'b111111111;
assign micromatrizz[84][260] = 9'b111111111;
assign micromatrizz[84][261] = 9'b111111111;
assign micromatrizz[84][262] = 9'b111111111;
assign micromatrizz[84][263] = 9'b111111111;
assign micromatrizz[84][264] = 9'b111111111;
assign micromatrizz[84][265] = 9'b111111111;
assign micromatrizz[84][266] = 9'b111111111;
assign micromatrizz[84][267] = 9'b111111111;
assign micromatrizz[84][268] = 9'b111111111;
assign micromatrizz[84][269] = 9'b111111111;
assign micromatrizz[84][270] = 9'b111111111;
assign micromatrizz[84][271] = 9'b111111111;
assign micromatrizz[84][272] = 9'b111111111;
assign micromatrizz[84][273] = 9'b111111111;
assign micromatrizz[84][274] = 9'b111111111;
assign micromatrizz[84][275] = 9'b111111111;
assign micromatrizz[84][276] = 9'b111111111;
assign micromatrizz[84][277] = 9'b111111111;
assign micromatrizz[84][278] = 9'b111111111;
assign micromatrizz[84][279] = 9'b111111111;
assign micromatrizz[84][280] = 9'b111111111;
assign micromatrizz[84][281] = 9'b111111111;
assign micromatrizz[84][282] = 9'b111111111;
assign micromatrizz[84][283] = 9'b111111111;
assign micromatrizz[84][284] = 9'b111111111;
assign micromatrizz[84][285] = 9'b111111111;
assign micromatrizz[84][286] = 9'b111111111;
assign micromatrizz[84][287] = 9'b111111111;
assign micromatrizz[84][288] = 9'b111111111;
assign micromatrizz[84][289] = 9'b111111111;
assign micromatrizz[84][290] = 9'b111111111;
assign micromatrizz[84][291] = 9'b111111111;
assign micromatrizz[84][292] = 9'b111111111;
assign micromatrizz[84][293] = 9'b111111111;
assign micromatrizz[84][294] = 9'b111111111;
assign micromatrizz[84][295] = 9'b111111111;
assign micromatrizz[84][296] = 9'b111111111;
assign micromatrizz[84][297] = 9'b111111111;
assign micromatrizz[84][298] = 9'b111111111;
assign micromatrizz[84][299] = 9'b111111111;
assign micromatrizz[84][300] = 9'b111111111;
assign micromatrizz[84][301] = 9'b111111111;
assign micromatrizz[84][302] = 9'b111111111;
assign micromatrizz[84][303] = 9'b111111111;
assign micromatrizz[84][304] = 9'b111111111;
assign micromatrizz[84][305] = 9'b111111111;
assign micromatrizz[84][306] = 9'b111111111;
assign micromatrizz[84][307] = 9'b111111111;
assign micromatrizz[84][308] = 9'b111111111;
assign micromatrizz[84][309] = 9'b111111111;
assign micromatrizz[84][310] = 9'b111111111;
assign micromatrizz[84][311] = 9'b111111111;
assign micromatrizz[84][312] = 9'b111111111;
assign micromatrizz[84][313] = 9'b111111111;
assign micromatrizz[84][314] = 9'b111111111;
assign micromatrizz[84][315] = 9'b111111111;
assign micromatrizz[84][316] = 9'b111111111;
assign micromatrizz[84][317] = 9'b111111111;
assign micromatrizz[84][318] = 9'b111111111;
assign micromatrizz[84][319] = 9'b111111111;
assign micromatrizz[84][320] = 9'b111111111;
assign micromatrizz[84][321] = 9'b111111111;
assign micromatrizz[84][322] = 9'b111111111;
assign micromatrizz[84][323] = 9'b111111111;
assign micromatrizz[84][324] = 9'b111111111;
assign micromatrizz[84][325] = 9'b111111111;
assign micromatrizz[84][326] = 9'b111111111;
assign micromatrizz[84][327] = 9'b111111111;
assign micromatrizz[84][328] = 9'b111111111;
assign micromatrizz[84][329] = 9'b111111111;
assign micromatrizz[84][330] = 9'b111111111;
assign micromatrizz[84][331] = 9'b111111111;
assign micromatrizz[84][332] = 9'b111111111;
assign micromatrizz[84][333] = 9'b111111111;
assign micromatrizz[84][334] = 9'b111111111;
assign micromatrizz[84][335] = 9'b111111111;
assign micromatrizz[84][336] = 9'b111111111;
assign micromatrizz[84][337] = 9'b111111111;
assign micromatrizz[84][338] = 9'b111111111;
assign micromatrizz[84][339] = 9'b111111111;
assign micromatrizz[84][340] = 9'b111111111;
assign micromatrizz[84][341] = 9'b111111111;
assign micromatrizz[84][342] = 9'b111111111;
assign micromatrizz[84][343] = 9'b111111111;
assign micromatrizz[84][344] = 9'b111111111;
assign micromatrizz[84][345] = 9'b111111111;
assign micromatrizz[84][346] = 9'b111111111;
assign micromatrizz[84][347] = 9'b111111111;
assign micromatrizz[84][348] = 9'b111111111;
assign micromatrizz[84][349] = 9'b111111111;
assign micromatrizz[84][350] = 9'b111111111;
assign micromatrizz[84][351] = 9'b111111111;
assign micromatrizz[84][352] = 9'b111111111;
assign micromatrizz[84][353] = 9'b111111111;
assign micromatrizz[84][354] = 9'b111111111;
assign micromatrizz[84][355] = 9'b111111111;
assign micromatrizz[84][356] = 9'b111111111;
assign micromatrizz[84][357] = 9'b111111111;
assign micromatrizz[84][358] = 9'b111111111;
assign micromatrizz[84][359] = 9'b111111111;
assign micromatrizz[84][360] = 9'b111111111;
assign micromatrizz[84][361] = 9'b111111111;
assign micromatrizz[84][362] = 9'b111111111;
assign micromatrizz[84][363] = 9'b111111111;
assign micromatrizz[84][364] = 9'b111111111;
assign micromatrizz[84][365] = 9'b111111111;
assign micromatrizz[84][366] = 9'b111111111;
assign micromatrizz[84][367] = 9'b111111111;
assign micromatrizz[84][368] = 9'b111111111;
assign micromatrizz[84][369] = 9'b111111111;
assign micromatrizz[84][370] = 9'b111111111;
assign micromatrizz[84][371] = 9'b111111111;
assign micromatrizz[84][372] = 9'b111111111;
assign micromatrizz[84][373] = 9'b111111111;
assign micromatrizz[84][374] = 9'b111111111;
assign micromatrizz[84][375] = 9'b111111111;
assign micromatrizz[84][376] = 9'b111111111;
assign micromatrizz[84][377] = 9'b111111111;
assign micromatrizz[84][378] = 9'b111111111;
assign micromatrizz[84][379] = 9'b111111111;
assign micromatrizz[84][380] = 9'b111111111;
assign micromatrizz[84][381] = 9'b111111111;
assign micromatrizz[84][382] = 9'b111111111;
assign micromatrizz[84][383] = 9'b111111111;
assign micromatrizz[84][384] = 9'b111111111;
assign micromatrizz[84][385] = 9'b111111111;
assign micromatrizz[84][386] = 9'b111111111;
assign micromatrizz[84][387] = 9'b111111111;
assign micromatrizz[84][388] = 9'b111111111;
assign micromatrizz[84][389] = 9'b111111111;
assign micromatrizz[84][390] = 9'b111111111;
assign micromatrizz[84][391] = 9'b111111111;
assign micromatrizz[84][392] = 9'b111111111;
assign micromatrizz[84][393] = 9'b111111111;
assign micromatrizz[84][394] = 9'b111111111;
assign micromatrizz[84][395] = 9'b111111111;
assign micromatrizz[84][396] = 9'b111111111;
assign micromatrizz[84][397] = 9'b111111111;
assign micromatrizz[84][398] = 9'b111111111;
assign micromatrizz[84][399] = 9'b111111111;
assign micromatrizz[84][400] = 9'b111111111;
assign micromatrizz[84][401] = 9'b111111111;
assign micromatrizz[84][402] = 9'b111111111;
assign micromatrizz[84][403] = 9'b111111111;
assign micromatrizz[84][404] = 9'b111111111;
assign micromatrizz[84][405] = 9'b111111111;
assign micromatrizz[84][406] = 9'b111111111;
assign micromatrizz[84][407] = 9'b111111111;
assign micromatrizz[84][408] = 9'b111111111;
assign micromatrizz[84][409] = 9'b111111111;
assign micromatrizz[84][410] = 9'b111111111;
assign micromatrizz[84][411] = 9'b111111111;
assign micromatrizz[84][412] = 9'b111111111;
assign micromatrizz[84][413] = 9'b111111111;
assign micromatrizz[84][414] = 9'b111111111;
assign micromatrizz[84][415] = 9'b111111111;
assign micromatrizz[84][416] = 9'b111111111;
assign micromatrizz[84][417] = 9'b111111111;
assign micromatrizz[84][418] = 9'b111111111;
assign micromatrizz[84][419] = 9'b111111111;
assign micromatrizz[84][420] = 9'b111111111;
assign micromatrizz[84][421] = 9'b111111111;
assign micromatrizz[84][422] = 9'b111111111;
assign micromatrizz[84][423] = 9'b111111111;
assign micromatrizz[84][424] = 9'b111111111;
assign micromatrizz[84][425] = 9'b111111111;
assign micromatrizz[84][426] = 9'b111111111;
assign micromatrizz[84][427] = 9'b111111111;
assign micromatrizz[84][428] = 9'b111111111;
assign micromatrizz[84][429] = 9'b111111111;
assign micromatrizz[84][430] = 9'b111111111;
assign micromatrizz[84][431] = 9'b111111111;
assign micromatrizz[84][432] = 9'b111111111;
assign micromatrizz[84][433] = 9'b111111111;
assign micromatrizz[84][434] = 9'b111111111;
assign micromatrizz[84][435] = 9'b111111111;
assign micromatrizz[84][436] = 9'b111111111;
assign micromatrizz[84][437] = 9'b111111111;
assign micromatrizz[84][438] = 9'b111111111;
assign micromatrizz[84][439] = 9'b111111111;
assign micromatrizz[84][440] = 9'b111111111;
assign micromatrizz[84][441] = 9'b111111111;
assign micromatrizz[84][442] = 9'b111111111;
assign micromatrizz[84][443] = 9'b111111111;
assign micromatrizz[84][444] = 9'b111111111;
assign micromatrizz[84][445] = 9'b111111111;
assign micromatrizz[84][446] = 9'b111111111;
assign micromatrizz[84][447] = 9'b111111111;
assign micromatrizz[84][448] = 9'b111111111;
assign micromatrizz[84][449] = 9'b111111111;
assign micromatrizz[84][450] = 9'b111111111;
assign micromatrizz[84][451] = 9'b111111111;
assign micromatrizz[84][452] = 9'b111111111;
assign micromatrizz[84][453] = 9'b111111111;
assign micromatrizz[84][454] = 9'b111111111;
assign micromatrizz[84][455] = 9'b111111111;
assign micromatrizz[84][456] = 9'b111111111;
assign micromatrizz[84][457] = 9'b111111111;
assign micromatrizz[84][458] = 9'b111111111;
assign micromatrizz[84][459] = 9'b111111111;
assign micromatrizz[84][460] = 9'b111111111;
assign micromatrizz[84][461] = 9'b111111111;
assign micromatrizz[84][462] = 9'b111111111;
assign micromatrizz[84][463] = 9'b111111111;
assign micromatrizz[84][464] = 9'b111111111;
assign micromatrizz[84][465] = 9'b111111111;
assign micromatrizz[84][466] = 9'b111111111;
assign micromatrizz[84][467] = 9'b111111111;
assign micromatrizz[84][468] = 9'b111111111;
assign micromatrizz[84][469] = 9'b111111111;
assign micromatrizz[84][470] = 9'b111111111;
assign micromatrizz[84][471] = 9'b111111111;
assign micromatrizz[84][472] = 9'b111111111;
assign micromatrizz[84][473] = 9'b111111111;
assign micromatrizz[84][474] = 9'b111111111;
assign micromatrizz[84][475] = 9'b111111111;
assign micromatrizz[84][476] = 9'b111111111;
assign micromatrizz[84][477] = 9'b111111111;
assign micromatrizz[84][478] = 9'b111111111;
assign micromatrizz[84][479] = 9'b111111111;
assign micromatrizz[84][480] = 9'b111111111;
assign micromatrizz[84][481] = 9'b111111111;
assign micromatrizz[84][482] = 9'b111111111;
assign micromatrizz[84][483] = 9'b111111111;
assign micromatrizz[84][484] = 9'b111111111;
assign micromatrizz[84][485] = 9'b111111111;
assign micromatrizz[84][486] = 9'b111111111;
assign micromatrizz[84][487] = 9'b111111111;
assign micromatrizz[84][488] = 9'b111111111;
assign micromatrizz[84][489] = 9'b111111111;
assign micromatrizz[84][490] = 9'b111111111;
assign micromatrizz[84][491] = 9'b111111111;
assign micromatrizz[84][492] = 9'b111111111;
assign micromatrizz[84][493] = 9'b111111111;
assign micromatrizz[84][494] = 9'b111111111;
assign micromatrizz[84][495] = 9'b111111111;
assign micromatrizz[84][496] = 9'b111111111;
assign micromatrizz[84][497] = 9'b111111111;
assign micromatrizz[84][498] = 9'b111111111;
assign micromatrizz[84][499] = 9'b111111111;
assign micromatrizz[84][500] = 9'b111111111;
assign micromatrizz[84][501] = 9'b111111111;
assign micromatrizz[84][502] = 9'b111111111;
assign micromatrizz[84][503] = 9'b111111111;
assign micromatrizz[84][504] = 9'b111111111;
assign micromatrizz[84][505] = 9'b111111111;
assign micromatrizz[84][506] = 9'b111111111;
assign micromatrizz[84][507] = 9'b111111111;
assign micromatrizz[84][508] = 9'b111111111;
assign micromatrizz[84][509] = 9'b111111111;
assign micromatrizz[84][510] = 9'b111111111;
assign micromatrizz[84][511] = 9'b111111111;
assign micromatrizz[84][512] = 9'b111111111;
assign micromatrizz[84][513] = 9'b111111111;
assign micromatrizz[84][514] = 9'b111111111;
assign micromatrizz[84][515] = 9'b111111111;
assign micromatrizz[84][516] = 9'b111111111;
assign micromatrizz[84][517] = 9'b111111111;
assign micromatrizz[84][518] = 9'b111111111;
assign micromatrizz[84][519] = 9'b111111111;
assign micromatrizz[84][520] = 9'b111111111;
assign micromatrizz[84][521] = 9'b111111111;
assign micromatrizz[84][522] = 9'b111111111;
assign micromatrizz[84][523] = 9'b111111111;
assign micromatrizz[84][524] = 9'b111111111;
assign micromatrizz[84][525] = 9'b111111111;
assign micromatrizz[84][526] = 9'b111111111;
assign micromatrizz[84][527] = 9'b111111111;
assign micromatrizz[84][528] = 9'b111111111;
assign micromatrizz[84][529] = 9'b111111111;
assign micromatrizz[84][530] = 9'b111111111;
assign micromatrizz[84][531] = 9'b111111111;
assign micromatrizz[84][532] = 9'b111111111;
assign micromatrizz[84][533] = 9'b111111111;
assign micromatrizz[84][534] = 9'b111111111;
assign micromatrizz[84][535] = 9'b111111111;
assign micromatrizz[84][536] = 9'b111111111;
assign micromatrizz[84][537] = 9'b111111111;
assign micromatrizz[84][538] = 9'b111111111;
assign micromatrizz[84][539] = 9'b111111111;
assign micromatrizz[84][540] = 9'b111111111;
assign micromatrizz[84][541] = 9'b111111111;
assign micromatrizz[84][542] = 9'b111111111;
assign micromatrizz[84][543] = 9'b111111111;
assign micromatrizz[84][544] = 9'b111111111;
assign micromatrizz[84][545] = 9'b111111111;
assign micromatrizz[84][546] = 9'b111111111;
assign micromatrizz[84][547] = 9'b111111111;
assign micromatrizz[84][548] = 9'b111111111;
assign micromatrizz[84][549] = 9'b111111111;
assign micromatrizz[84][550] = 9'b111111111;
assign micromatrizz[84][551] = 9'b111111111;
assign micromatrizz[84][552] = 9'b111111111;
assign micromatrizz[84][553] = 9'b111111111;
assign micromatrizz[84][554] = 9'b111111111;
assign micromatrizz[84][555] = 9'b111111111;
assign micromatrizz[84][556] = 9'b111111111;
assign micromatrizz[84][557] = 9'b111111111;
assign micromatrizz[84][558] = 9'b111111111;
assign micromatrizz[84][559] = 9'b111111111;
assign micromatrizz[84][560] = 9'b111111111;
assign micromatrizz[84][561] = 9'b111111111;
assign micromatrizz[84][562] = 9'b111111111;
assign micromatrizz[84][563] = 9'b111111111;
assign micromatrizz[84][564] = 9'b111111111;
assign micromatrizz[84][565] = 9'b111111111;
assign micromatrizz[84][566] = 9'b111111111;
assign micromatrizz[84][567] = 9'b111111111;
assign micromatrizz[84][568] = 9'b111111111;
assign micromatrizz[84][569] = 9'b111111111;
assign micromatrizz[84][570] = 9'b111111111;
assign micromatrizz[84][571] = 9'b111111111;
assign micromatrizz[84][572] = 9'b111111111;
assign micromatrizz[84][573] = 9'b111111111;
assign micromatrizz[84][574] = 9'b111111111;
assign micromatrizz[84][575] = 9'b111111111;
assign micromatrizz[84][576] = 9'b111111111;
assign micromatrizz[84][577] = 9'b111111111;
assign micromatrizz[84][578] = 9'b111111111;
assign micromatrizz[84][579] = 9'b111111111;
assign micromatrizz[84][580] = 9'b111111111;
assign micromatrizz[84][581] = 9'b111111111;
assign micromatrizz[84][582] = 9'b111111111;
assign micromatrizz[84][583] = 9'b111111111;
assign micromatrizz[84][584] = 9'b111111111;
assign micromatrizz[84][585] = 9'b111111111;
assign micromatrizz[84][586] = 9'b111111111;
assign micromatrizz[84][587] = 9'b111111111;
assign micromatrizz[84][588] = 9'b111111111;
assign micromatrizz[84][589] = 9'b111111111;
assign micromatrizz[84][590] = 9'b111111111;
assign micromatrizz[84][591] = 9'b111111111;
assign micromatrizz[84][592] = 9'b111111111;
assign micromatrizz[84][593] = 9'b111111111;
assign micromatrizz[84][594] = 9'b111111111;
assign micromatrizz[84][595] = 9'b111111111;
assign micromatrizz[84][596] = 9'b111111111;
assign micromatrizz[84][597] = 9'b111111111;
assign micromatrizz[84][598] = 9'b111111111;
assign micromatrizz[84][599] = 9'b111111111;
assign micromatrizz[84][600] = 9'b111111111;
assign micromatrizz[84][601] = 9'b111111111;
assign micromatrizz[84][602] = 9'b111111111;
assign micromatrizz[84][603] = 9'b111111111;
assign micromatrizz[84][604] = 9'b111111111;
assign micromatrizz[84][605] = 9'b111111111;
assign micromatrizz[84][606] = 9'b111111111;
assign micromatrizz[84][607] = 9'b111111111;
assign micromatrizz[84][608] = 9'b111111111;
assign micromatrizz[84][609] = 9'b111111111;
assign micromatrizz[84][610] = 9'b111111111;
assign micromatrizz[84][611] = 9'b111111111;
assign micromatrizz[84][612] = 9'b111111111;
assign micromatrizz[84][613] = 9'b111111111;
assign micromatrizz[84][614] = 9'b111111111;
assign micromatrizz[84][615] = 9'b111111111;
assign micromatrizz[84][616] = 9'b111111111;
assign micromatrizz[84][617] = 9'b111111111;
assign micromatrizz[84][618] = 9'b111111111;
assign micromatrizz[84][619] = 9'b111111111;
assign micromatrizz[84][620] = 9'b111111111;
assign micromatrizz[84][621] = 9'b111111111;
assign micromatrizz[84][622] = 9'b111111111;
assign micromatrizz[84][623] = 9'b111111111;
assign micromatrizz[84][624] = 9'b111111111;
assign micromatrizz[84][625] = 9'b111111111;
assign micromatrizz[84][626] = 9'b111111111;
assign micromatrizz[84][627] = 9'b111111111;
assign micromatrizz[84][628] = 9'b111111111;
assign micromatrizz[84][629] = 9'b111111111;
assign micromatrizz[84][630] = 9'b111111111;
assign micromatrizz[84][631] = 9'b111111111;
assign micromatrizz[84][632] = 9'b111111111;
assign micromatrizz[84][633] = 9'b111111111;
assign micromatrizz[84][634] = 9'b111111111;
assign micromatrizz[84][635] = 9'b111111111;
assign micromatrizz[84][636] = 9'b111111111;
assign micromatrizz[84][637] = 9'b111111111;
assign micromatrizz[84][638] = 9'b111111111;
assign micromatrizz[84][639] = 9'b111111111;
assign micromatrizz[85][0] = 9'b111111111;
assign micromatrizz[85][1] = 9'b111111111;
assign micromatrizz[85][2] = 9'b111111111;
assign micromatrizz[85][3] = 9'b111111111;
assign micromatrizz[85][4] = 9'b111111111;
assign micromatrizz[85][5] = 9'b111111111;
assign micromatrizz[85][6] = 9'b111111111;
assign micromatrizz[85][7] = 9'b111111111;
assign micromatrizz[85][8] = 9'b111111111;
assign micromatrizz[85][9] = 9'b111111111;
assign micromatrizz[85][10] = 9'b111111111;
assign micromatrizz[85][11] = 9'b111111111;
assign micromatrizz[85][12] = 9'b111111111;
assign micromatrizz[85][13] = 9'b111111111;
assign micromatrizz[85][14] = 9'b111111111;
assign micromatrizz[85][15] = 9'b111111111;
assign micromatrizz[85][16] = 9'b111111111;
assign micromatrizz[85][17] = 9'b111111111;
assign micromatrizz[85][18] = 9'b111111111;
assign micromatrizz[85][19] = 9'b111111111;
assign micromatrizz[85][20] = 9'b111111111;
assign micromatrizz[85][21] = 9'b111111111;
assign micromatrizz[85][22] = 9'b111111111;
assign micromatrizz[85][23] = 9'b111111111;
assign micromatrizz[85][24] = 9'b111111111;
assign micromatrizz[85][25] = 9'b111111111;
assign micromatrizz[85][26] = 9'b111111111;
assign micromatrizz[85][27] = 9'b111111111;
assign micromatrizz[85][28] = 9'b111111111;
assign micromatrizz[85][29] = 9'b111111111;
assign micromatrizz[85][30] = 9'b111111111;
assign micromatrizz[85][31] = 9'b111111111;
assign micromatrizz[85][32] = 9'b111111111;
assign micromatrizz[85][33] = 9'b111111111;
assign micromatrizz[85][34] = 9'b111111111;
assign micromatrizz[85][35] = 9'b111111111;
assign micromatrizz[85][36] = 9'b111111111;
assign micromatrizz[85][37] = 9'b111111111;
assign micromatrizz[85][38] = 9'b111111111;
assign micromatrizz[85][39] = 9'b111111111;
assign micromatrizz[85][40] = 9'b111111111;
assign micromatrizz[85][41] = 9'b111111111;
assign micromatrizz[85][42] = 9'b111111111;
assign micromatrizz[85][43] = 9'b111111111;
assign micromatrizz[85][44] = 9'b111111111;
assign micromatrizz[85][45] = 9'b111111111;
assign micromatrizz[85][46] = 9'b111111111;
assign micromatrizz[85][47] = 9'b111111111;
assign micromatrizz[85][48] = 9'b111111111;
assign micromatrizz[85][49] = 9'b111111111;
assign micromatrizz[85][50] = 9'b111111111;
assign micromatrizz[85][51] = 9'b111111111;
assign micromatrizz[85][52] = 9'b111111111;
assign micromatrizz[85][53] = 9'b111111111;
assign micromatrizz[85][54] = 9'b111111111;
assign micromatrizz[85][55] = 9'b111111111;
assign micromatrizz[85][56] = 9'b111111111;
assign micromatrizz[85][57] = 9'b111111111;
assign micromatrizz[85][58] = 9'b111111111;
assign micromatrizz[85][59] = 9'b111111111;
assign micromatrizz[85][60] = 9'b111111111;
assign micromatrizz[85][61] = 9'b111111111;
assign micromatrizz[85][62] = 9'b111111111;
assign micromatrizz[85][63] = 9'b111111111;
assign micromatrizz[85][64] = 9'b111111111;
assign micromatrizz[85][65] = 9'b111111111;
assign micromatrizz[85][66] = 9'b111111111;
assign micromatrizz[85][67] = 9'b111111111;
assign micromatrizz[85][68] = 9'b111111111;
assign micromatrizz[85][69] = 9'b111111111;
assign micromatrizz[85][70] = 9'b111111111;
assign micromatrizz[85][71] = 9'b111111111;
assign micromatrizz[85][72] = 9'b111111111;
assign micromatrizz[85][73] = 9'b111111111;
assign micromatrizz[85][74] = 9'b111111111;
assign micromatrizz[85][75] = 9'b111111111;
assign micromatrizz[85][76] = 9'b111111111;
assign micromatrizz[85][77] = 9'b111111111;
assign micromatrizz[85][78] = 9'b111111111;
assign micromatrizz[85][79] = 9'b111111111;
assign micromatrizz[85][80] = 9'b111111111;
assign micromatrizz[85][81] = 9'b111111111;
assign micromatrizz[85][82] = 9'b111111111;
assign micromatrizz[85][83] = 9'b111111111;
assign micromatrizz[85][84] = 9'b111111111;
assign micromatrizz[85][85] = 9'b111111111;
assign micromatrizz[85][86] = 9'b111111111;
assign micromatrizz[85][87] = 9'b111111111;
assign micromatrizz[85][88] = 9'b111111111;
assign micromatrizz[85][89] = 9'b111111111;
assign micromatrizz[85][90] = 9'b111111111;
assign micromatrizz[85][91] = 9'b111111111;
assign micromatrizz[85][92] = 9'b111111111;
assign micromatrizz[85][93] = 9'b111111111;
assign micromatrizz[85][94] = 9'b111111111;
assign micromatrizz[85][95] = 9'b111111111;
assign micromatrizz[85][96] = 9'b111111111;
assign micromatrizz[85][97] = 9'b111111111;
assign micromatrizz[85][98] = 9'b111111111;
assign micromatrizz[85][99] = 9'b111111111;
assign micromatrizz[85][100] = 9'b111111111;
assign micromatrizz[85][101] = 9'b111111111;
assign micromatrizz[85][102] = 9'b111111111;
assign micromatrizz[85][103] = 9'b111111111;
assign micromatrizz[85][104] = 9'b111111111;
assign micromatrizz[85][105] = 9'b111111111;
assign micromatrizz[85][106] = 9'b111111111;
assign micromatrizz[85][107] = 9'b111111111;
assign micromatrizz[85][108] = 9'b111111111;
assign micromatrizz[85][109] = 9'b111111111;
assign micromatrizz[85][110] = 9'b111111111;
assign micromatrizz[85][111] = 9'b111111111;
assign micromatrizz[85][112] = 9'b111111111;
assign micromatrizz[85][113] = 9'b111111111;
assign micromatrizz[85][114] = 9'b111111111;
assign micromatrizz[85][115] = 9'b111111111;
assign micromatrizz[85][116] = 9'b111111111;
assign micromatrizz[85][117] = 9'b111111111;
assign micromatrizz[85][118] = 9'b111111111;
assign micromatrizz[85][119] = 9'b111111111;
assign micromatrizz[85][120] = 9'b111111111;
assign micromatrizz[85][121] = 9'b111111111;
assign micromatrizz[85][122] = 9'b111111111;
assign micromatrizz[85][123] = 9'b111111111;
assign micromatrizz[85][124] = 9'b111111111;
assign micromatrizz[85][125] = 9'b111111111;
assign micromatrizz[85][126] = 9'b111111111;
assign micromatrizz[85][127] = 9'b111111111;
assign micromatrizz[85][128] = 9'b111111111;
assign micromatrizz[85][129] = 9'b111111111;
assign micromatrizz[85][130] = 9'b111111111;
assign micromatrizz[85][131] = 9'b111111111;
assign micromatrizz[85][132] = 9'b111111111;
assign micromatrizz[85][133] = 9'b111111111;
assign micromatrizz[85][134] = 9'b111111111;
assign micromatrizz[85][135] = 9'b111111111;
assign micromatrizz[85][136] = 9'b111111111;
assign micromatrizz[85][137] = 9'b111111111;
assign micromatrizz[85][138] = 9'b111111111;
assign micromatrizz[85][139] = 9'b111111111;
assign micromatrizz[85][140] = 9'b111111111;
assign micromatrizz[85][141] = 9'b111111111;
assign micromatrizz[85][142] = 9'b111111111;
assign micromatrizz[85][143] = 9'b111111111;
assign micromatrizz[85][144] = 9'b111111111;
assign micromatrizz[85][145] = 9'b111111111;
assign micromatrizz[85][146] = 9'b111111111;
assign micromatrizz[85][147] = 9'b111111111;
assign micromatrizz[85][148] = 9'b111111111;
assign micromatrizz[85][149] = 9'b111111111;
assign micromatrizz[85][150] = 9'b111111111;
assign micromatrizz[85][151] = 9'b111111111;
assign micromatrizz[85][152] = 9'b111111111;
assign micromatrizz[85][153] = 9'b111111111;
assign micromatrizz[85][154] = 9'b111111111;
assign micromatrizz[85][155] = 9'b111111111;
assign micromatrizz[85][156] = 9'b111111111;
assign micromatrizz[85][157] = 9'b111111111;
assign micromatrizz[85][158] = 9'b111111111;
assign micromatrizz[85][159] = 9'b111111111;
assign micromatrizz[85][160] = 9'b111111111;
assign micromatrizz[85][161] = 9'b111111111;
assign micromatrizz[85][162] = 9'b111111111;
assign micromatrizz[85][163] = 9'b111111111;
assign micromatrizz[85][164] = 9'b111111111;
assign micromatrizz[85][165] = 9'b111111111;
assign micromatrizz[85][166] = 9'b111111111;
assign micromatrizz[85][167] = 9'b111111111;
assign micromatrizz[85][168] = 9'b111111111;
assign micromatrizz[85][169] = 9'b111111111;
assign micromatrizz[85][170] = 9'b111111111;
assign micromatrizz[85][171] = 9'b111111111;
assign micromatrizz[85][172] = 9'b111111111;
assign micromatrizz[85][173] = 9'b111111111;
assign micromatrizz[85][174] = 9'b111111111;
assign micromatrizz[85][175] = 9'b111111111;
assign micromatrizz[85][176] = 9'b111111111;
assign micromatrizz[85][177] = 9'b111111111;
assign micromatrizz[85][178] = 9'b111111111;
assign micromatrizz[85][179] = 9'b111111111;
assign micromatrizz[85][180] = 9'b111111111;
assign micromatrizz[85][181] = 9'b111111111;
assign micromatrizz[85][182] = 9'b111111111;
assign micromatrizz[85][183] = 9'b111111111;
assign micromatrizz[85][184] = 9'b111111111;
assign micromatrizz[85][185] = 9'b111111111;
assign micromatrizz[85][186] = 9'b111111111;
assign micromatrizz[85][187] = 9'b111111111;
assign micromatrizz[85][188] = 9'b111111111;
assign micromatrizz[85][189] = 9'b111111111;
assign micromatrizz[85][190] = 9'b111111111;
assign micromatrizz[85][191] = 9'b111111111;
assign micromatrizz[85][192] = 9'b111111111;
assign micromatrizz[85][193] = 9'b111111111;
assign micromatrizz[85][194] = 9'b111111111;
assign micromatrizz[85][195] = 9'b111111111;
assign micromatrizz[85][196] = 9'b111111111;
assign micromatrizz[85][197] = 9'b111111111;
assign micromatrizz[85][198] = 9'b111111111;
assign micromatrizz[85][199] = 9'b111111111;
assign micromatrizz[85][200] = 9'b111111111;
assign micromatrizz[85][201] = 9'b111111111;
assign micromatrizz[85][202] = 9'b111111111;
assign micromatrizz[85][203] = 9'b111111111;
assign micromatrizz[85][204] = 9'b111111111;
assign micromatrizz[85][205] = 9'b111111111;
assign micromatrizz[85][206] = 9'b111111111;
assign micromatrizz[85][207] = 9'b111111111;
assign micromatrizz[85][208] = 9'b111111111;
assign micromatrizz[85][209] = 9'b111111111;
assign micromatrizz[85][210] = 9'b111111111;
assign micromatrizz[85][211] = 9'b111111111;
assign micromatrizz[85][212] = 9'b111111111;
assign micromatrizz[85][213] = 9'b111111111;
assign micromatrizz[85][214] = 9'b111111111;
assign micromatrizz[85][215] = 9'b111111111;
assign micromatrizz[85][216] = 9'b111111111;
assign micromatrizz[85][217] = 9'b111111111;
assign micromatrizz[85][218] = 9'b111111111;
assign micromatrizz[85][219] = 9'b111111111;
assign micromatrizz[85][220] = 9'b111111111;
assign micromatrizz[85][221] = 9'b111111111;
assign micromatrizz[85][222] = 9'b111111111;
assign micromatrizz[85][223] = 9'b111111111;
assign micromatrizz[85][224] = 9'b111111111;
assign micromatrizz[85][225] = 9'b111111111;
assign micromatrizz[85][226] = 9'b111111111;
assign micromatrizz[85][227] = 9'b111111111;
assign micromatrizz[85][228] = 9'b111111111;
assign micromatrizz[85][229] = 9'b111111111;
assign micromatrizz[85][230] = 9'b111111111;
assign micromatrizz[85][231] = 9'b111111111;
assign micromatrizz[85][232] = 9'b111111111;
assign micromatrizz[85][233] = 9'b111111111;
assign micromatrizz[85][234] = 9'b111111111;
assign micromatrizz[85][235] = 9'b111111111;
assign micromatrizz[85][236] = 9'b111111111;
assign micromatrizz[85][237] = 9'b111111111;
assign micromatrizz[85][238] = 9'b111111111;
assign micromatrizz[85][239] = 9'b111111111;
assign micromatrizz[85][240] = 9'b111111111;
assign micromatrizz[85][241] = 9'b111111111;
assign micromatrizz[85][242] = 9'b111111111;
assign micromatrizz[85][243] = 9'b111111111;
assign micromatrizz[85][244] = 9'b111111111;
assign micromatrizz[85][245] = 9'b111111111;
assign micromatrizz[85][246] = 9'b111111111;
assign micromatrizz[85][247] = 9'b111111111;
assign micromatrizz[85][248] = 9'b111111111;
assign micromatrizz[85][249] = 9'b111111111;
assign micromatrizz[85][250] = 9'b111111111;
assign micromatrizz[85][251] = 9'b111111111;
assign micromatrizz[85][252] = 9'b111111111;
assign micromatrizz[85][253] = 9'b111111111;
assign micromatrizz[85][254] = 9'b111111111;
assign micromatrizz[85][255] = 9'b111111111;
assign micromatrizz[85][256] = 9'b111111111;
assign micromatrizz[85][257] = 9'b111111111;
assign micromatrizz[85][258] = 9'b111111111;
assign micromatrizz[85][259] = 9'b111111111;
assign micromatrizz[85][260] = 9'b111111111;
assign micromatrizz[85][261] = 9'b111111111;
assign micromatrizz[85][262] = 9'b111111111;
assign micromatrizz[85][263] = 9'b111111111;
assign micromatrizz[85][264] = 9'b111111111;
assign micromatrizz[85][265] = 9'b111111111;
assign micromatrizz[85][266] = 9'b111111111;
assign micromatrizz[85][267] = 9'b111111111;
assign micromatrizz[85][268] = 9'b111111111;
assign micromatrizz[85][269] = 9'b111111111;
assign micromatrizz[85][270] = 9'b111111111;
assign micromatrizz[85][271] = 9'b111111111;
assign micromatrizz[85][272] = 9'b111111111;
assign micromatrizz[85][273] = 9'b111111111;
assign micromatrizz[85][274] = 9'b111111111;
assign micromatrizz[85][275] = 9'b111111111;
assign micromatrizz[85][276] = 9'b111111111;
assign micromatrizz[85][277] = 9'b111111111;
assign micromatrizz[85][278] = 9'b111111111;
assign micromatrizz[85][279] = 9'b111111111;
assign micromatrizz[85][280] = 9'b111111111;
assign micromatrizz[85][281] = 9'b111111111;
assign micromatrizz[85][282] = 9'b111111111;
assign micromatrizz[85][283] = 9'b111111111;
assign micromatrizz[85][284] = 9'b111111111;
assign micromatrizz[85][285] = 9'b111111111;
assign micromatrizz[85][286] = 9'b111111111;
assign micromatrizz[85][287] = 9'b111111111;
assign micromatrizz[85][288] = 9'b111111111;
assign micromatrizz[85][289] = 9'b111111111;
assign micromatrizz[85][290] = 9'b111111111;
assign micromatrizz[85][291] = 9'b111111111;
assign micromatrizz[85][292] = 9'b111111111;
assign micromatrizz[85][293] = 9'b111111111;
assign micromatrizz[85][294] = 9'b111111111;
assign micromatrizz[85][295] = 9'b111111111;
assign micromatrizz[85][296] = 9'b111111111;
assign micromatrizz[85][297] = 9'b111111111;
assign micromatrizz[85][298] = 9'b111111111;
assign micromatrizz[85][299] = 9'b111111111;
assign micromatrizz[85][300] = 9'b111111111;
assign micromatrizz[85][301] = 9'b111111111;
assign micromatrizz[85][302] = 9'b111111111;
assign micromatrizz[85][303] = 9'b111111111;
assign micromatrizz[85][304] = 9'b111111111;
assign micromatrizz[85][305] = 9'b111111111;
assign micromatrizz[85][306] = 9'b111111111;
assign micromatrizz[85][307] = 9'b111111111;
assign micromatrizz[85][308] = 9'b111111111;
assign micromatrizz[85][309] = 9'b111111111;
assign micromatrizz[85][310] = 9'b111111111;
assign micromatrizz[85][311] = 9'b111111111;
assign micromatrizz[85][312] = 9'b111111111;
assign micromatrizz[85][313] = 9'b111111111;
assign micromatrizz[85][314] = 9'b111111111;
assign micromatrizz[85][315] = 9'b111111111;
assign micromatrizz[85][316] = 9'b111111111;
assign micromatrizz[85][317] = 9'b111111111;
assign micromatrizz[85][318] = 9'b111111111;
assign micromatrizz[85][319] = 9'b111111111;
assign micromatrizz[85][320] = 9'b111111111;
assign micromatrizz[85][321] = 9'b111111111;
assign micromatrizz[85][322] = 9'b111111111;
assign micromatrizz[85][323] = 9'b111111111;
assign micromatrizz[85][324] = 9'b111111111;
assign micromatrizz[85][325] = 9'b111111111;
assign micromatrizz[85][326] = 9'b111111111;
assign micromatrizz[85][327] = 9'b111111111;
assign micromatrizz[85][328] = 9'b111111111;
assign micromatrizz[85][329] = 9'b111111111;
assign micromatrizz[85][330] = 9'b111111111;
assign micromatrizz[85][331] = 9'b111111111;
assign micromatrizz[85][332] = 9'b111111111;
assign micromatrizz[85][333] = 9'b111111111;
assign micromatrizz[85][334] = 9'b111111111;
assign micromatrizz[85][335] = 9'b111111111;
assign micromatrizz[85][336] = 9'b111111111;
assign micromatrizz[85][337] = 9'b111111111;
assign micromatrizz[85][338] = 9'b111111111;
assign micromatrizz[85][339] = 9'b111111111;
assign micromatrizz[85][340] = 9'b111111111;
assign micromatrizz[85][341] = 9'b111111111;
assign micromatrizz[85][342] = 9'b111111111;
assign micromatrizz[85][343] = 9'b111111111;
assign micromatrizz[85][344] = 9'b111111111;
assign micromatrizz[85][345] = 9'b111111111;
assign micromatrizz[85][346] = 9'b111111111;
assign micromatrizz[85][347] = 9'b111111111;
assign micromatrizz[85][348] = 9'b111111111;
assign micromatrizz[85][349] = 9'b111111111;
assign micromatrizz[85][350] = 9'b111111111;
assign micromatrizz[85][351] = 9'b111111111;
assign micromatrizz[85][352] = 9'b111111111;
assign micromatrizz[85][353] = 9'b111111111;
assign micromatrizz[85][354] = 9'b111111111;
assign micromatrizz[85][355] = 9'b111111111;
assign micromatrizz[85][356] = 9'b111111111;
assign micromatrizz[85][357] = 9'b111111111;
assign micromatrizz[85][358] = 9'b111111111;
assign micromatrizz[85][359] = 9'b111111111;
assign micromatrizz[85][360] = 9'b111111111;
assign micromatrizz[85][361] = 9'b111111111;
assign micromatrizz[85][362] = 9'b111111111;
assign micromatrizz[85][363] = 9'b111111111;
assign micromatrizz[85][364] = 9'b111111111;
assign micromatrizz[85][365] = 9'b111111111;
assign micromatrizz[85][366] = 9'b111111111;
assign micromatrizz[85][367] = 9'b111111111;
assign micromatrizz[85][368] = 9'b111111111;
assign micromatrizz[85][369] = 9'b111111111;
assign micromatrizz[85][370] = 9'b111111111;
assign micromatrizz[85][371] = 9'b111111111;
assign micromatrizz[85][372] = 9'b111111111;
assign micromatrizz[85][373] = 9'b111111111;
assign micromatrizz[85][374] = 9'b111111111;
assign micromatrizz[85][375] = 9'b111111111;
assign micromatrizz[85][376] = 9'b111111111;
assign micromatrizz[85][377] = 9'b111111111;
assign micromatrizz[85][378] = 9'b111111111;
assign micromatrizz[85][379] = 9'b111111111;
assign micromatrizz[85][380] = 9'b111111111;
assign micromatrizz[85][381] = 9'b111111111;
assign micromatrizz[85][382] = 9'b111111111;
assign micromatrizz[85][383] = 9'b111111111;
assign micromatrizz[85][384] = 9'b111111111;
assign micromatrizz[85][385] = 9'b111111111;
assign micromatrizz[85][386] = 9'b111111111;
assign micromatrizz[85][387] = 9'b111111111;
assign micromatrizz[85][388] = 9'b111111111;
assign micromatrizz[85][389] = 9'b111111111;
assign micromatrizz[85][390] = 9'b111111111;
assign micromatrizz[85][391] = 9'b111111111;
assign micromatrizz[85][392] = 9'b111111111;
assign micromatrizz[85][393] = 9'b111111111;
assign micromatrizz[85][394] = 9'b111111111;
assign micromatrizz[85][395] = 9'b111111111;
assign micromatrizz[85][396] = 9'b111111111;
assign micromatrizz[85][397] = 9'b111111111;
assign micromatrizz[85][398] = 9'b111111111;
assign micromatrizz[85][399] = 9'b111111111;
assign micromatrizz[85][400] = 9'b111111111;
assign micromatrizz[85][401] = 9'b111111111;
assign micromatrizz[85][402] = 9'b111111111;
assign micromatrizz[85][403] = 9'b111111111;
assign micromatrizz[85][404] = 9'b111111111;
assign micromatrizz[85][405] = 9'b111111111;
assign micromatrizz[85][406] = 9'b111111111;
assign micromatrizz[85][407] = 9'b111111111;
assign micromatrizz[85][408] = 9'b111111111;
assign micromatrizz[85][409] = 9'b111111111;
assign micromatrizz[85][410] = 9'b111111111;
assign micromatrizz[85][411] = 9'b111111111;
assign micromatrizz[85][412] = 9'b111111111;
assign micromatrizz[85][413] = 9'b111111111;
assign micromatrizz[85][414] = 9'b111111111;
assign micromatrizz[85][415] = 9'b111111111;
assign micromatrizz[85][416] = 9'b111111111;
assign micromatrizz[85][417] = 9'b111111111;
assign micromatrizz[85][418] = 9'b111111111;
assign micromatrizz[85][419] = 9'b111111111;
assign micromatrizz[85][420] = 9'b111111111;
assign micromatrizz[85][421] = 9'b111111111;
assign micromatrizz[85][422] = 9'b111111111;
assign micromatrizz[85][423] = 9'b111111111;
assign micromatrizz[85][424] = 9'b111111111;
assign micromatrizz[85][425] = 9'b111111111;
assign micromatrizz[85][426] = 9'b111111111;
assign micromatrizz[85][427] = 9'b111111111;
assign micromatrizz[85][428] = 9'b111111111;
assign micromatrizz[85][429] = 9'b111111111;
assign micromatrizz[85][430] = 9'b111111111;
assign micromatrizz[85][431] = 9'b111111111;
assign micromatrizz[85][432] = 9'b111111111;
assign micromatrizz[85][433] = 9'b111111111;
assign micromatrizz[85][434] = 9'b111111111;
assign micromatrizz[85][435] = 9'b111111111;
assign micromatrizz[85][436] = 9'b111111111;
assign micromatrizz[85][437] = 9'b111111111;
assign micromatrizz[85][438] = 9'b111111111;
assign micromatrizz[85][439] = 9'b111111111;
assign micromatrizz[85][440] = 9'b111111111;
assign micromatrizz[85][441] = 9'b111111111;
assign micromatrizz[85][442] = 9'b111111111;
assign micromatrizz[85][443] = 9'b111111111;
assign micromatrizz[85][444] = 9'b111111111;
assign micromatrizz[85][445] = 9'b111111111;
assign micromatrizz[85][446] = 9'b111111111;
assign micromatrizz[85][447] = 9'b111111111;
assign micromatrizz[85][448] = 9'b111111111;
assign micromatrizz[85][449] = 9'b111111111;
assign micromatrizz[85][450] = 9'b111111111;
assign micromatrizz[85][451] = 9'b111111111;
assign micromatrizz[85][452] = 9'b111111111;
assign micromatrizz[85][453] = 9'b111111111;
assign micromatrizz[85][454] = 9'b111111111;
assign micromatrizz[85][455] = 9'b111111111;
assign micromatrizz[85][456] = 9'b111111111;
assign micromatrizz[85][457] = 9'b111111111;
assign micromatrizz[85][458] = 9'b111111111;
assign micromatrizz[85][459] = 9'b111111111;
assign micromatrizz[85][460] = 9'b111111111;
assign micromatrizz[85][461] = 9'b111111111;
assign micromatrizz[85][462] = 9'b111111111;
assign micromatrizz[85][463] = 9'b111111111;
assign micromatrizz[85][464] = 9'b111111111;
assign micromatrizz[85][465] = 9'b111111111;
assign micromatrizz[85][466] = 9'b111111111;
assign micromatrizz[85][467] = 9'b111111111;
assign micromatrizz[85][468] = 9'b111111111;
assign micromatrizz[85][469] = 9'b111111111;
assign micromatrizz[85][470] = 9'b111111111;
assign micromatrizz[85][471] = 9'b111111111;
assign micromatrizz[85][472] = 9'b111111111;
assign micromatrizz[85][473] = 9'b111111111;
assign micromatrizz[85][474] = 9'b111111111;
assign micromatrizz[85][475] = 9'b111111111;
assign micromatrizz[85][476] = 9'b111111111;
assign micromatrizz[85][477] = 9'b111111111;
assign micromatrizz[85][478] = 9'b111111111;
assign micromatrizz[85][479] = 9'b111111111;
assign micromatrizz[85][480] = 9'b111111111;
assign micromatrizz[85][481] = 9'b111111111;
assign micromatrizz[85][482] = 9'b111111111;
assign micromatrizz[85][483] = 9'b111111111;
assign micromatrizz[85][484] = 9'b111111111;
assign micromatrizz[85][485] = 9'b111111111;
assign micromatrizz[85][486] = 9'b111111111;
assign micromatrizz[85][487] = 9'b111111111;
assign micromatrizz[85][488] = 9'b111111111;
assign micromatrizz[85][489] = 9'b111111111;
assign micromatrizz[85][490] = 9'b111111111;
assign micromatrizz[85][491] = 9'b111111111;
assign micromatrizz[85][492] = 9'b111111111;
assign micromatrizz[85][493] = 9'b111111111;
assign micromatrizz[85][494] = 9'b111111111;
assign micromatrizz[85][495] = 9'b111111111;
assign micromatrizz[85][496] = 9'b111111111;
assign micromatrizz[85][497] = 9'b111111111;
assign micromatrizz[85][498] = 9'b111111111;
assign micromatrizz[85][499] = 9'b111111111;
assign micromatrizz[85][500] = 9'b111111111;
assign micromatrizz[85][501] = 9'b111111111;
assign micromatrizz[85][502] = 9'b111111111;
assign micromatrizz[85][503] = 9'b111111111;
assign micromatrizz[85][504] = 9'b111111111;
assign micromatrizz[85][505] = 9'b111111111;
assign micromatrizz[85][506] = 9'b111111111;
assign micromatrizz[85][507] = 9'b111111111;
assign micromatrizz[85][508] = 9'b111111111;
assign micromatrizz[85][509] = 9'b111111111;
assign micromatrizz[85][510] = 9'b111111111;
assign micromatrizz[85][511] = 9'b111111111;
assign micromatrizz[85][512] = 9'b111111111;
assign micromatrizz[85][513] = 9'b111111111;
assign micromatrizz[85][514] = 9'b111111111;
assign micromatrizz[85][515] = 9'b111111111;
assign micromatrizz[85][516] = 9'b111111111;
assign micromatrizz[85][517] = 9'b111111111;
assign micromatrizz[85][518] = 9'b111111111;
assign micromatrizz[85][519] = 9'b111111111;
assign micromatrizz[85][520] = 9'b111111111;
assign micromatrizz[85][521] = 9'b111111111;
assign micromatrizz[85][522] = 9'b111111111;
assign micromatrizz[85][523] = 9'b111111111;
assign micromatrizz[85][524] = 9'b111111111;
assign micromatrizz[85][525] = 9'b111111111;
assign micromatrizz[85][526] = 9'b111111111;
assign micromatrizz[85][527] = 9'b111111111;
assign micromatrizz[85][528] = 9'b111111111;
assign micromatrizz[85][529] = 9'b111111111;
assign micromatrizz[85][530] = 9'b111111111;
assign micromatrizz[85][531] = 9'b111111111;
assign micromatrizz[85][532] = 9'b111111111;
assign micromatrizz[85][533] = 9'b111111111;
assign micromatrizz[85][534] = 9'b111111111;
assign micromatrizz[85][535] = 9'b111111111;
assign micromatrizz[85][536] = 9'b111111111;
assign micromatrizz[85][537] = 9'b111111111;
assign micromatrizz[85][538] = 9'b111111111;
assign micromatrizz[85][539] = 9'b111111111;
assign micromatrizz[85][540] = 9'b111111111;
assign micromatrizz[85][541] = 9'b111111111;
assign micromatrizz[85][542] = 9'b111111111;
assign micromatrizz[85][543] = 9'b111111111;
assign micromatrizz[85][544] = 9'b111111111;
assign micromatrizz[85][545] = 9'b111111111;
assign micromatrizz[85][546] = 9'b111111111;
assign micromatrizz[85][547] = 9'b111111111;
assign micromatrizz[85][548] = 9'b111111111;
assign micromatrizz[85][549] = 9'b111111111;
assign micromatrizz[85][550] = 9'b111111111;
assign micromatrizz[85][551] = 9'b111111111;
assign micromatrizz[85][552] = 9'b111111111;
assign micromatrizz[85][553] = 9'b111111111;
assign micromatrizz[85][554] = 9'b111111111;
assign micromatrizz[85][555] = 9'b111111111;
assign micromatrizz[85][556] = 9'b111111111;
assign micromatrizz[85][557] = 9'b111111111;
assign micromatrizz[85][558] = 9'b111111111;
assign micromatrizz[85][559] = 9'b111111111;
assign micromatrizz[85][560] = 9'b111111111;
assign micromatrizz[85][561] = 9'b111111111;
assign micromatrizz[85][562] = 9'b111111111;
assign micromatrizz[85][563] = 9'b111111111;
assign micromatrizz[85][564] = 9'b111111111;
assign micromatrizz[85][565] = 9'b111111111;
assign micromatrizz[85][566] = 9'b111111111;
assign micromatrizz[85][567] = 9'b111111111;
assign micromatrizz[85][568] = 9'b111111111;
assign micromatrizz[85][569] = 9'b111111111;
assign micromatrizz[85][570] = 9'b111111111;
assign micromatrizz[85][571] = 9'b111111111;
assign micromatrizz[85][572] = 9'b111111111;
assign micromatrizz[85][573] = 9'b111111111;
assign micromatrizz[85][574] = 9'b111111111;
assign micromatrizz[85][575] = 9'b111111111;
assign micromatrizz[85][576] = 9'b111111111;
assign micromatrizz[85][577] = 9'b111111111;
assign micromatrizz[85][578] = 9'b111111111;
assign micromatrizz[85][579] = 9'b111111111;
assign micromatrizz[85][580] = 9'b111111111;
assign micromatrizz[85][581] = 9'b111111111;
assign micromatrizz[85][582] = 9'b111111111;
assign micromatrizz[85][583] = 9'b111111111;
assign micromatrizz[85][584] = 9'b111111111;
assign micromatrizz[85][585] = 9'b111111111;
assign micromatrizz[85][586] = 9'b111111111;
assign micromatrizz[85][587] = 9'b111111111;
assign micromatrizz[85][588] = 9'b111111111;
assign micromatrizz[85][589] = 9'b111111111;
assign micromatrizz[85][590] = 9'b111111111;
assign micromatrizz[85][591] = 9'b111111111;
assign micromatrizz[85][592] = 9'b111111111;
assign micromatrizz[85][593] = 9'b111111111;
assign micromatrizz[85][594] = 9'b111111111;
assign micromatrizz[85][595] = 9'b111111111;
assign micromatrizz[85][596] = 9'b111111111;
assign micromatrizz[85][597] = 9'b111111111;
assign micromatrizz[85][598] = 9'b111111111;
assign micromatrizz[85][599] = 9'b111111111;
assign micromatrizz[85][600] = 9'b111111111;
assign micromatrizz[85][601] = 9'b111111111;
assign micromatrizz[85][602] = 9'b111111111;
assign micromatrizz[85][603] = 9'b111111111;
assign micromatrizz[85][604] = 9'b111111111;
assign micromatrizz[85][605] = 9'b111111111;
assign micromatrizz[85][606] = 9'b111111111;
assign micromatrizz[85][607] = 9'b111111111;
assign micromatrizz[85][608] = 9'b111111111;
assign micromatrizz[85][609] = 9'b111111111;
assign micromatrizz[85][610] = 9'b111111111;
assign micromatrizz[85][611] = 9'b111111111;
assign micromatrizz[85][612] = 9'b111111111;
assign micromatrizz[85][613] = 9'b111111111;
assign micromatrizz[85][614] = 9'b111111111;
assign micromatrizz[85][615] = 9'b111111111;
assign micromatrizz[85][616] = 9'b111111111;
assign micromatrizz[85][617] = 9'b111111111;
assign micromatrizz[85][618] = 9'b111111111;
assign micromatrizz[85][619] = 9'b111111111;
assign micromatrizz[85][620] = 9'b111111111;
assign micromatrizz[85][621] = 9'b111111111;
assign micromatrizz[85][622] = 9'b111111111;
assign micromatrizz[85][623] = 9'b111111111;
assign micromatrizz[85][624] = 9'b111111111;
assign micromatrizz[85][625] = 9'b111111111;
assign micromatrizz[85][626] = 9'b111111111;
assign micromatrizz[85][627] = 9'b111111111;
assign micromatrizz[85][628] = 9'b111111111;
assign micromatrizz[85][629] = 9'b111111111;
assign micromatrizz[85][630] = 9'b111111111;
assign micromatrizz[85][631] = 9'b111111111;
assign micromatrizz[85][632] = 9'b111111111;
assign micromatrizz[85][633] = 9'b111111111;
assign micromatrizz[85][634] = 9'b111111111;
assign micromatrizz[85][635] = 9'b111111111;
assign micromatrizz[85][636] = 9'b111111111;
assign micromatrizz[85][637] = 9'b111111111;
assign micromatrizz[85][638] = 9'b111111111;
assign micromatrizz[85][639] = 9'b111111111;
assign micromatrizz[86][0] = 9'b111111111;
assign micromatrizz[86][1] = 9'b111111111;
assign micromatrizz[86][2] = 9'b111111111;
assign micromatrizz[86][3] = 9'b111111111;
assign micromatrizz[86][4] = 9'b111111111;
assign micromatrizz[86][5] = 9'b111111111;
assign micromatrizz[86][6] = 9'b111111111;
assign micromatrizz[86][7] = 9'b111111111;
assign micromatrizz[86][8] = 9'b111111111;
assign micromatrizz[86][9] = 9'b111111111;
assign micromatrizz[86][10] = 9'b111111111;
assign micromatrizz[86][11] = 9'b111111111;
assign micromatrizz[86][12] = 9'b111111111;
assign micromatrizz[86][13] = 9'b111111111;
assign micromatrizz[86][14] = 9'b111111111;
assign micromatrizz[86][15] = 9'b111111111;
assign micromatrizz[86][16] = 9'b111111111;
assign micromatrizz[86][17] = 9'b111111111;
assign micromatrizz[86][18] = 9'b111111111;
assign micromatrizz[86][19] = 9'b111111111;
assign micromatrizz[86][20] = 9'b111111111;
assign micromatrizz[86][21] = 9'b111111111;
assign micromatrizz[86][22] = 9'b111111111;
assign micromatrizz[86][23] = 9'b111111111;
assign micromatrizz[86][24] = 9'b111111111;
assign micromatrizz[86][25] = 9'b111111111;
assign micromatrizz[86][26] = 9'b111111111;
assign micromatrizz[86][27] = 9'b111111111;
assign micromatrizz[86][28] = 9'b111111111;
assign micromatrizz[86][29] = 9'b111111111;
assign micromatrizz[86][30] = 9'b111111111;
assign micromatrizz[86][31] = 9'b111111111;
assign micromatrizz[86][32] = 9'b111111111;
assign micromatrizz[86][33] = 9'b111111111;
assign micromatrizz[86][34] = 9'b111111111;
assign micromatrizz[86][35] = 9'b111111111;
assign micromatrizz[86][36] = 9'b111111111;
assign micromatrizz[86][37] = 9'b111111111;
assign micromatrizz[86][38] = 9'b111111111;
assign micromatrizz[86][39] = 9'b111111111;
assign micromatrizz[86][40] = 9'b111111111;
assign micromatrizz[86][41] = 9'b111111111;
assign micromatrizz[86][42] = 9'b111111111;
assign micromatrizz[86][43] = 9'b111111111;
assign micromatrizz[86][44] = 9'b111111111;
assign micromatrizz[86][45] = 9'b111111111;
assign micromatrizz[86][46] = 9'b111111111;
assign micromatrizz[86][47] = 9'b111111111;
assign micromatrizz[86][48] = 9'b111111111;
assign micromatrizz[86][49] = 9'b111111111;
assign micromatrizz[86][50] = 9'b111111111;
assign micromatrizz[86][51] = 9'b111111111;
assign micromatrizz[86][52] = 9'b111111111;
assign micromatrizz[86][53] = 9'b111111111;
assign micromatrizz[86][54] = 9'b111111111;
assign micromatrizz[86][55] = 9'b111111111;
assign micromatrizz[86][56] = 9'b111111111;
assign micromatrizz[86][57] = 9'b111111111;
assign micromatrizz[86][58] = 9'b111111111;
assign micromatrizz[86][59] = 9'b111111111;
assign micromatrizz[86][60] = 9'b111111111;
assign micromatrizz[86][61] = 9'b111111111;
assign micromatrizz[86][62] = 9'b111111111;
assign micromatrizz[86][63] = 9'b111111111;
assign micromatrizz[86][64] = 9'b111111111;
assign micromatrizz[86][65] = 9'b111111111;
assign micromatrizz[86][66] = 9'b111111111;
assign micromatrizz[86][67] = 9'b111111111;
assign micromatrizz[86][68] = 9'b111111111;
assign micromatrizz[86][69] = 9'b111111111;
assign micromatrizz[86][70] = 9'b111111111;
assign micromatrizz[86][71] = 9'b111111111;
assign micromatrizz[86][72] = 9'b111111111;
assign micromatrizz[86][73] = 9'b111111111;
assign micromatrizz[86][74] = 9'b111111111;
assign micromatrizz[86][75] = 9'b111111111;
assign micromatrizz[86][76] = 9'b111111111;
assign micromatrizz[86][77] = 9'b111111111;
assign micromatrizz[86][78] = 9'b111111111;
assign micromatrizz[86][79] = 9'b111111111;
assign micromatrizz[86][80] = 9'b111111111;
assign micromatrizz[86][81] = 9'b111111111;
assign micromatrizz[86][82] = 9'b111111111;
assign micromatrizz[86][83] = 9'b111111111;
assign micromatrizz[86][84] = 9'b111111111;
assign micromatrizz[86][85] = 9'b111111111;
assign micromatrizz[86][86] = 9'b111111111;
assign micromatrizz[86][87] = 9'b111111111;
assign micromatrizz[86][88] = 9'b111111111;
assign micromatrizz[86][89] = 9'b111111111;
assign micromatrizz[86][90] = 9'b111111111;
assign micromatrizz[86][91] = 9'b111111111;
assign micromatrizz[86][92] = 9'b111111111;
assign micromatrizz[86][93] = 9'b111111111;
assign micromatrizz[86][94] = 9'b111111111;
assign micromatrizz[86][95] = 9'b111111111;
assign micromatrizz[86][96] = 9'b111111111;
assign micromatrizz[86][97] = 9'b111111111;
assign micromatrizz[86][98] = 9'b111111111;
assign micromatrizz[86][99] = 9'b111111111;
assign micromatrizz[86][100] = 9'b111111111;
assign micromatrizz[86][101] = 9'b111111111;
assign micromatrizz[86][102] = 9'b111111111;
assign micromatrizz[86][103] = 9'b111111111;
assign micromatrizz[86][104] = 9'b111111111;
assign micromatrizz[86][105] = 9'b111111111;
assign micromatrizz[86][106] = 9'b111111111;
assign micromatrizz[86][107] = 9'b111111111;
assign micromatrizz[86][108] = 9'b111111111;
assign micromatrizz[86][109] = 9'b111111111;
assign micromatrizz[86][110] = 9'b111111111;
assign micromatrizz[86][111] = 9'b111111111;
assign micromatrizz[86][112] = 9'b111111111;
assign micromatrizz[86][113] = 9'b111111111;
assign micromatrizz[86][114] = 9'b111111111;
assign micromatrizz[86][115] = 9'b111111111;
assign micromatrizz[86][116] = 9'b111111111;
assign micromatrizz[86][117] = 9'b111111111;
assign micromatrizz[86][118] = 9'b111111111;
assign micromatrizz[86][119] = 9'b111111111;
assign micromatrizz[86][120] = 9'b111111111;
assign micromatrizz[86][121] = 9'b111111111;
assign micromatrizz[86][122] = 9'b111111111;
assign micromatrizz[86][123] = 9'b111111111;
assign micromatrizz[86][124] = 9'b111111111;
assign micromatrizz[86][125] = 9'b111111111;
assign micromatrizz[86][126] = 9'b111111111;
assign micromatrizz[86][127] = 9'b111111111;
assign micromatrizz[86][128] = 9'b111111111;
assign micromatrizz[86][129] = 9'b111111111;
assign micromatrizz[86][130] = 9'b111111111;
assign micromatrizz[86][131] = 9'b111111111;
assign micromatrizz[86][132] = 9'b111111111;
assign micromatrizz[86][133] = 9'b111111111;
assign micromatrizz[86][134] = 9'b111111111;
assign micromatrizz[86][135] = 9'b111111111;
assign micromatrizz[86][136] = 9'b111111111;
assign micromatrizz[86][137] = 9'b111111111;
assign micromatrizz[86][138] = 9'b111111111;
assign micromatrizz[86][139] = 9'b111111111;
assign micromatrizz[86][140] = 9'b111111111;
assign micromatrizz[86][141] = 9'b111111111;
assign micromatrizz[86][142] = 9'b111111111;
assign micromatrizz[86][143] = 9'b111111111;
assign micromatrizz[86][144] = 9'b111111111;
assign micromatrizz[86][145] = 9'b111111111;
assign micromatrizz[86][146] = 9'b111111111;
assign micromatrizz[86][147] = 9'b111111111;
assign micromatrizz[86][148] = 9'b111111111;
assign micromatrizz[86][149] = 9'b111111111;
assign micromatrizz[86][150] = 9'b111111111;
assign micromatrizz[86][151] = 9'b111111111;
assign micromatrizz[86][152] = 9'b111111111;
assign micromatrizz[86][153] = 9'b111111111;
assign micromatrizz[86][154] = 9'b111111111;
assign micromatrizz[86][155] = 9'b111111111;
assign micromatrizz[86][156] = 9'b111111111;
assign micromatrizz[86][157] = 9'b111111111;
assign micromatrizz[86][158] = 9'b111111111;
assign micromatrizz[86][159] = 9'b111111111;
assign micromatrizz[86][160] = 9'b111111111;
assign micromatrizz[86][161] = 9'b111111111;
assign micromatrizz[86][162] = 9'b111111111;
assign micromatrizz[86][163] = 9'b111111111;
assign micromatrizz[86][164] = 9'b111111111;
assign micromatrizz[86][165] = 9'b111111111;
assign micromatrizz[86][166] = 9'b111111111;
assign micromatrizz[86][167] = 9'b111111111;
assign micromatrizz[86][168] = 9'b111111111;
assign micromatrizz[86][169] = 9'b111111111;
assign micromatrizz[86][170] = 9'b111111111;
assign micromatrizz[86][171] = 9'b111111111;
assign micromatrizz[86][172] = 9'b111111111;
assign micromatrizz[86][173] = 9'b111111111;
assign micromatrizz[86][174] = 9'b111111111;
assign micromatrizz[86][175] = 9'b111111111;
assign micromatrizz[86][176] = 9'b111111111;
assign micromatrizz[86][177] = 9'b111111111;
assign micromatrizz[86][178] = 9'b111111111;
assign micromatrizz[86][179] = 9'b111111111;
assign micromatrizz[86][180] = 9'b111111111;
assign micromatrizz[86][181] = 9'b111111111;
assign micromatrizz[86][182] = 9'b111111111;
assign micromatrizz[86][183] = 9'b111111111;
assign micromatrizz[86][184] = 9'b111111111;
assign micromatrizz[86][185] = 9'b111111111;
assign micromatrizz[86][186] = 9'b111111111;
assign micromatrizz[86][187] = 9'b111111111;
assign micromatrizz[86][188] = 9'b111111111;
assign micromatrizz[86][189] = 9'b111111111;
assign micromatrizz[86][190] = 9'b111111111;
assign micromatrizz[86][191] = 9'b111111111;
assign micromatrizz[86][192] = 9'b111111111;
assign micromatrizz[86][193] = 9'b111111111;
assign micromatrizz[86][194] = 9'b111111111;
assign micromatrizz[86][195] = 9'b111111111;
assign micromatrizz[86][196] = 9'b111111111;
assign micromatrizz[86][197] = 9'b111111111;
assign micromatrizz[86][198] = 9'b111111111;
assign micromatrizz[86][199] = 9'b111111111;
assign micromatrizz[86][200] = 9'b111111111;
assign micromatrizz[86][201] = 9'b111111111;
assign micromatrizz[86][202] = 9'b111111111;
assign micromatrizz[86][203] = 9'b111111111;
assign micromatrizz[86][204] = 9'b111111111;
assign micromatrizz[86][205] = 9'b111111111;
assign micromatrizz[86][206] = 9'b111111111;
assign micromatrizz[86][207] = 9'b111111111;
assign micromatrizz[86][208] = 9'b111111111;
assign micromatrizz[86][209] = 9'b111111111;
assign micromatrizz[86][210] = 9'b111111111;
assign micromatrizz[86][211] = 9'b111111111;
assign micromatrizz[86][212] = 9'b111111111;
assign micromatrizz[86][213] = 9'b111111111;
assign micromatrizz[86][214] = 9'b111111111;
assign micromatrizz[86][215] = 9'b111111111;
assign micromatrizz[86][216] = 9'b111111111;
assign micromatrizz[86][217] = 9'b111111111;
assign micromatrizz[86][218] = 9'b111111111;
assign micromatrizz[86][219] = 9'b111111111;
assign micromatrizz[86][220] = 9'b111111111;
assign micromatrizz[86][221] = 9'b111111111;
assign micromatrizz[86][222] = 9'b111111111;
assign micromatrizz[86][223] = 9'b111111111;
assign micromatrizz[86][224] = 9'b111111111;
assign micromatrizz[86][225] = 9'b111111111;
assign micromatrizz[86][226] = 9'b111111111;
assign micromatrizz[86][227] = 9'b111111111;
assign micromatrizz[86][228] = 9'b111111111;
assign micromatrizz[86][229] = 9'b111111111;
assign micromatrizz[86][230] = 9'b111111111;
assign micromatrizz[86][231] = 9'b111111111;
assign micromatrizz[86][232] = 9'b111111111;
assign micromatrizz[86][233] = 9'b111111111;
assign micromatrizz[86][234] = 9'b111111111;
assign micromatrizz[86][235] = 9'b111111111;
assign micromatrizz[86][236] = 9'b111111111;
assign micromatrizz[86][237] = 9'b111111111;
assign micromatrizz[86][238] = 9'b111111111;
assign micromatrizz[86][239] = 9'b111111111;
assign micromatrizz[86][240] = 9'b111111111;
assign micromatrizz[86][241] = 9'b111111111;
assign micromatrizz[86][242] = 9'b111111111;
assign micromatrizz[86][243] = 9'b111111111;
assign micromatrizz[86][244] = 9'b111111111;
assign micromatrizz[86][245] = 9'b111111111;
assign micromatrizz[86][246] = 9'b111111111;
assign micromatrizz[86][247] = 9'b111111111;
assign micromatrizz[86][248] = 9'b111111111;
assign micromatrizz[86][249] = 9'b111111111;
assign micromatrizz[86][250] = 9'b111111111;
assign micromatrizz[86][251] = 9'b111111111;
assign micromatrizz[86][252] = 9'b111111111;
assign micromatrizz[86][253] = 9'b111111111;
assign micromatrizz[86][254] = 9'b111111111;
assign micromatrizz[86][255] = 9'b111111111;
assign micromatrizz[86][256] = 9'b111111111;
assign micromatrizz[86][257] = 9'b111111111;
assign micromatrizz[86][258] = 9'b111111111;
assign micromatrizz[86][259] = 9'b111111111;
assign micromatrizz[86][260] = 9'b111111111;
assign micromatrizz[86][261] = 9'b111111111;
assign micromatrizz[86][262] = 9'b111111111;
assign micromatrizz[86][263] = 9'b111111111;
assign micromatrizz[86][264] = 9'b111111111;
assign micromatrizz[86][265] = 9'b111111111;
assign micromatrizz[86][266] = 9'b111111111;
assign micromatrizz[86][267] = 9'b111111111;
assign micromatrizz[86][268] = 9'b111111111;
assign micromatrizz[86][269] = 9'b111111111;
assign micromatrizz[86][270] = 9'b111111111;
assign micromatrizz[86][271] = 9'b111111111;
assign micromatrizz[86][272] = 9'b111111111;
assign micromatrizz[86][273] = 9'b111111111;
assign micromatrizz[86][274] = 9'b111111111;
assign micromatrizz[86][275] = 9'b111111111;
assign micromatrizz[86][276] = 9'b111111111;
assign micromatrizz[86][277] = 9'b111111111;
assign micromatrizz[86][278] = 9'b111111111;
assign micromatrizz[86][279] = 9'b111111111;
assign micromatrizz[86][280] = 9'b111111111;
assign micromatrizz[86][281] = 9'b111111111;
assign micromatrizz[86][282] = 9'b111111111;
assign micromatrizz[86][283] = 9'b111111111;
assign micromatrizz[86][284] = 9'b111111111;
assign micromatrizz[86][285] = 9'b111111111;
assign micromatrizz[86][286] = 9'b111111111;
assign micromatrizz[86][287] = 9'b111111111;
assign micromatrizz[86][288] = 9'b111111111;
assign micromatrizz[86][289] = 9'b111111111;
assign micromatrizz[86][290] = 9'b111111111;
assign micromatrizz[86][291] = 9'b111111111;
assign micromatrizz[86][292] = 9'b111111111;
assign micromatrizz[86][293] = 9'b111111111;
assign micromatrizz[86][294] = 9'b111111111;
assign micromatrizz[86][295] = 9'b111111111;
assign micromatrizz[86][296] = 9'b111111111;
assign micromatrizz[86][297] = 9'b111111111;
assign micromatrizz[86][298] = 9'b111111111;
assign micromatrizz[86][299] = 9'b111111111;
assign micromatrizz[86][300] = 9'b111111111;
assign micromatrizz[86][301] = 9'b111111111;
assign micromatrizz[86][302] = 9'b111111111;
assign micromatrizz[86][303] = 9'b111111111;
assign micromatrizz[86][304] = 9'b111111111;
assign micromatrizz[86][305] = 9'b111111111;
assign micromatrizz[86][306] = 9'b111111111;
assign micromatrizz[86][307] = 9'b111111111;
assign micromatrizz[86][308] = 9'b111111111;
assign micromatrizz[86][309] = 9'b111111111;
assign micromatrizz[86][310] = 9'b111111111;
assign micromatrizz[86][311] = 9'b111111111;
assign micromatrizz[86][312] = 9'b111111111;
assign micromatrizz[86][313] = 9'b111111111;
assign micromatrizz[86][314] = 9'b111111111;
assign micromatrizz[86][315] = 9'b111111111;
assign micromatrizz[86][316] = 9'b111111111;
assign micromatrizz[86][317] = 9'b111111111;
assign micromatrizz[86][318] = 9'b111111111;
assign micromatrizz[86][319] = 9'b111111111;
assign micromatrizz[86][320] = 9'b111111111;
assign micromatrizz[86][321] = 9'b111111111;
assign micromatrizz[86][322] = 9'b111111111;
assign micromatrizz[86][323] = 9'b111111111;
assign micromatrizz[86][324] = 9'b111111111;
assign micromatrizz[86][325] = 9'b111111111;
assign micromatrizz[86][326] = 9'b111111111;
assign micromatrizz[86][327] = 9'b111111111;
assign micromatrizz[86][328] = 9'b111111111;
assign micromatrizz[86][329] = 9'b111111111;
assign micromatrizz[86][330] = 9'b111111111;
assign micromatrizz[86][331] = 9'b111111111;
assign micromatrizz[86][332] = 9'b111111111;
assign micromatrizz[86][333] = 9'b111111111;
assign micromatrizz[86][334] = 9'b111111111;
assign micromatrizz[86][335] = 9'b111111111;
assign micromatrizz[86][336] = 9'b111111111;
assign micromatrizz[86][337] = 9'b111111111;
assign micromatrizz[86][338] = 9'b111111111;
assign micromatrizz[86][339] = 9'b111111111;
assign micromatrizz[86][340] = 9'b111111111;
assign micromatrizz[86][341] = 9'b111111111;
assign micromatrizz[86][342] = 9'b111111111;
assign micromatrizz[86][343] = 9'b111111111;
assign micromatrizz[86][344] = 9'b111111111;
assign micromatrizz[86][345] = 9'b111111111;
assign micromatrizz[86][346] = 9'b111111111;
assign micromatrizz[86][347] = 9'b111111111;
assign micromatrizz[86][348] = 9'b111111111;
assign micromatrizz[86][349] = 9'b111111111;
assign micromatrizz[86][350] = 9'b111111111;
assign micromatrizz[86][351] = 9'b111111111;
assign micromatrizz[86][352] = 9'b111111111;
assign micromatrizz[86][353] = 9'b111111111;
assign micromatrizz[86][354] = 9'b111111111;
assign micromatrizz[86][355] = 9'b111111111;
assign micromatrizz[86][356] = 9'b111111111;
assign micromatrizz[86][357] = 9'b111111111;
assign micromatrizz[86][358] = 9'b111111111;
assign micromatrizz[86][359] = 9'b111111111;
assign micromatrizz[86][360] = 9'b111111111;
assign micromatrizz[86][361] = 9'b111111111;
assign micromatrizz[86][362] = 9'b111111111;
assign micromatrizz[86][363] = 9'b111111111;
assign micromatrizz[86][364] = 9'b111111111;
assign micromatrizz[86][365] = 9'b111111111;
assign micromatrizz[86][366] = 9'b111111111;
assign micromatrizz[86][367] = 9'b111111111;
assign micromatrizz[86][368] = 9'b111111111;
assign micromatrizz[86][369] = 9'b111111111;
assign micromatrizz[86][370] = 9'b111111111;
assign micromatrizz[86][371] = 9'b111111111;
assign micromatrizz[86][372] = 9'b111111111;
assign micromatrizz[86][373] = 9'b111111111;
assign micromatrizz[86][374] = 9'b111111111;
assign micromatrizz[86][375] = 9'b111111111;
assign micromatrizz[86][376] = 9'b111111111;
assign micromatrizz[86][377] = 9'b111111111;
assign micromatrizz[86][378] = 9'b111111111;
assign micromatrizz[86][379] = 9'b111111111;
assign micromatrizz[86][380] = 9'b111111111;
assign micromatrizz[86][381] = 9'b111111111;
assign micromatrizz[86][382] = 9'b111111111;
assign micromatrizz[86][383] = 9'b111111111;
assign micromatrizz[86][384] = 9'b111111111;
assign micromatrizz[86][385] = 9'b111111111;
assign micromatrizz[86][386] = 9'b111111111;
assign micromatrizz[86][387] = 9'b111111111;
assign micromatrizz[86][388] = 9'b111111111;
assign micromatrizz[86][389] = 9'b111111111;
assign micromatrizz[86][390] = 9'b111111111;
assign micromatrizz[86][391] = 9'b111111111;
assign micromatrizz[86][392] = 9'b111111111;
assign micromatrizz[86][393] = 9'b111111111;
assign micromatrizz[86][394] = 9'b111111111;
assign micromatrizz[86][395] = 9'b111111111;
assign micromatrizz[86][396] = 9'b111111111;
assign micromatrizz[86][397] = 9'b111111111;
assign micromatrizz[86][398] = 9'b111111111;
assign micromatrizz[86][399] = 9'b111111111;
assign micromatrizz[86][400] = 9'b111111111;
assign micromatrizz[86][401] = 9'b111111111;
assign micromatrizz[86][402] = 9'b111111111;
assign micromatrizz[86][403] = 9'b111111111;
assign micromatrizz[86][404] = 9'b111111111;
assign micromatrizz[86][405] = 9'b111111111;
assign micromatrizz[86][406] = 9'b111111111;
assign micromatrizz[86][407] = 9'b111111111;
assign micromatrizz[86][408] = 9'b111111111;
assign micromatrizz[86][409] = 9'b111111111;
assign micromatrizz[86][410] = 9'b111111111;
assign micromatrizz[86][411] = 9'b111111111;
assign micromatrizz[86][412] = 9'b111111111;
assign micromatrizz[86][413] = 9'b111111111;
assign micromatrizz[86][414] = 9'b111111111;
assign micromatrizz[86][415] = 9'b111111111;
assign micromatrizz[86][416] = 9'b111111111;
assign micromatrizz[86][417] = 9'b111111111;
assign micromatrizz[86][418] = 9'b111111111;
assign micromatrizz[86][419] = 9'b111111111;
assign micromatrizz[86][420] = 9'b111111111;
assign micromatrizz[86][421] = 9'b111111111;
assign micromatrizz[86][422] = 9'b111111111;
assign micromatrizz[86][423] = 9'b111111111;
assign micromatrizz[86][424] = 9'b111111111;
assign micromatrizz[86][425] = 9'b111111111;
assign micromatrizz[86][426] = 9'b111111111;
assign micromatrizz[86][427] = 9'b111111111;
assign micromatrizz[86][428] = 9'b111111111;
assign micromatrizz[86][429] = 9'b111111111;
assign micromatrizz[86][430] = 9'b111111111;
assign micromatrizz[86][431] = 9'b111111111;
assign micromatrizz[86][432] = 9'b111111111;
assign micromatrizz[86][433] = 9'b111111111;
assign micromatrizz[86][434] = 9'b111111111;
assign micromatrizz[86][435] = 9'b111111111;
assign micromatrizz[86][436] = 9'b111111111;
assign micromatrizz[86][437] = 9'b111111111;
assign micromatrizz[86][438] = 9'b111111111;
assign micromatrizz[86][439] = 9'b111111111;
assign micromatrizz[86][440] = 9'b111111111;
assign micromatrizz[86][441] = 9'b111111111;
assign micromatrizz[86][442] = 9'b111111111;
assign micromatrizz[86][443] = 9'b111111111;
assign micromatrizz[86][444] = 9'b111111111;
assign micromatrizz[86][445] = 9'b111111111;
assign micromatrizz[86][446] = 9'b111111111;
assign micromatrizz[86][447] = 9'b111111111;
assign micromatrizz[86][448] = 9'b111111111;
assign micromatrizz[86][449] = 9'b111111111;
assign micromatrizz[86][450] = 9'b111111111;
assign micromatrizz[86][451] = 9'b111111111;
assign micromatrizz[86][452] = 9'b111111111;
assign micromatrizz[86][453] = 9'b111111111;
assign micromatrizz[86][454] = 9'b111111111;
assign micromatrizz[86][455] = 9'b111111111;
assign micromatrizz[86][456] = 9'b111111111;
assign micromatrizz[86][457] = 9'b111111111;
assign micromatrizz[86][458] = 9'b111111111;
assign micromatrizz[86][459] = 9'b111111111;
assign micromatrizz[86][460] = 9'b111111111;
assign micromatrizz[86][461] = 9'b111111111;
assign micromatrizz[86][462] = 9'b111111111;
assign micromatrizz[86][463] = 9'b111111111;
assign micromatrizz[86][464] = 9'b111111111;
assign micromatrizz[86][465] = 9'b111111111;
assign micromatrizz[86][466] = 9'b111111111;
assign micromatrizz[86][467] = 9'b111111111;
assign micromatrizz[86][468] = 9'b111111111;
assign micromatrizz[86][469] = 9'b111111111;
assign micromatrizz[86][470] = 9'b111111111;
assign micromatrizz[86][471] = 9'b111111111;
assign micromatrizz[86][472] = 9'b111111111;
assign micromatrizz[86][473] = 9'b111111111;
assign micromatrizz[86][474] = 9'b111111111;
assign micromatrizz[86][475] = 9'b111111111;
assign micromatrizz[86][476] = 9'b111111111;
assign micromatrizz[86][477] = 9'b111111111;
assign micromatrizz[86][478] = 9'b111111111;
assign micromatrizz[86][479] = 9'b111111111;
assign micromatrizz[86][480] = 9'b111111111;
assign micromatrizz[86][481] = 9'b111111111;
assign micromatrizz[86][482] = 9'b111111111;
assign micromatrizz[86][483] = 9'b111111111;
assign micromatrizz[86][484] = 9'b111111111;
assign micromatrizz[86][485] = 9'b111111111;
assign micromatrizz[86][486] = 9'b111111111;
assign micromatrizz[86][487] = 9'b111111111;
assign micromatrizz[86][488] = 9'b111111111;
assign micromatrizz[86][489] = 9'b111111111;
assign micromatrizz[86][490] = 9'b111111111;
assign micromatrizz[86][491] = 9'b111111111;
assign micromatrizz[86][492] = 9'b111111111;
assign micromatrizz[86][493] = 9'b111111111;
assign micromatrizz[86][494] = 9'b111111111;
assign micromatrizz[86][495] = 9'b111111111;
assign micromatrizz[86][496] = 9'b111111111;
assign micromatrizz[86][497] = 9'b111111111;
assign micromatrizz[86][498] = 9'b111111111;
assign micromatrizz[86][499] = 9'b111111111;
assign micromatrizz[86][500] = 9'b111111111;
assign micromatrizz[86][501] = 9'b111111111;
assign micromatrizz[86][502] = 9'b111111111;
assign micromatrizz[86][503] = 9'b111111111;
assign micromatrizz[86][504] = 9'b111111111;
assign micromatrizz[86][505] = 9'b111111111;
assign micromatrizz[86][506] = 9'b111111111;
assign micromatrizz[86][507] = 9'b111111111;
assign micromatrizz[86][508] = 9'b111111111;
assign micromatrizz[86][509] = 9'b111111111;
assign micromatrizz[86][510] = 9'b111111111;
assign micromatrizz[86][511] = 9'b111111111;
assign micromatrizz[86][512] = 9'b111111111;
assign micromatrizz[86][513] = 9'b111111111;
assign micromatrizz[86][514] = 9'b111111111;
assign micromatrizz[86][515] = 9'b111111111;
assign micromatrizz[86][516] = 9'b111111111;
assign micromatrizz[86][517] = 9'b111111111;
assign micromatrizz[86][518] = 9'b111111111;
assign micromatrizz[86][519] = 9'b111111111;
assign micromatrizz[86][520] = 9'b111111111;
assign micromatrizz[86][521] = 9'b111111111;
assign micromatrizz[86][522] = 9'b111111111;
assign micromatrizz[86][523] = 9'b111111111;
assign micromatrizz[86][524] = 9'b111111111;
assign micromatrizz[86][525] = 9'b111111111;
assign micromatrizz[86][526] = 9'b111111111;
assign micromatrizz[86][527] = 9'b111111111;
assign micromatrizz[86][528] = 9'b111111111;
assign micromatrizz[86][529] = 9'b111111111;
assign micromatrizz[86][530] = 9'b111111111;
assign micromatrizz[86][531] = 9'b111111111;
assign micromatrizz[86][532] = 9'b111111111;
assign micromatrizz[86][533] = 9'b111111111;
assign micromatrizz[86][534] = 9'b111111111;
assign micromatrizz[86][535] = 9'b111111111;
assign micromatrizz[86][536] = 9'b111111111;
assign micromatrizz[86][537] = 9'b111111111;
assign micromatrizz[86][538] = 9'b111111111;
assign micromatrizz[86][539] = 9'b111111111;
assign micromatrizz[86][540] = 9'b111111111;
assign micromatrizz[86][541] = 9'b111111111;
assign micromatrizz[86][542] = 9'b111111111;
assign micromatrizz[86][543] = 9'b111111111;
assign micromatrizz[86][544] = 9'b111111111;
assign micromatrizz[86][545] = 9'b111111111;
assign micromatrizz[86][546] = 9'b111111111;
assign micromatrizz[86][547] = 9'b111111111;
assign micromatrizz[86][548] = 9'b111111111;
assign micromatrizz[86][549] = 9'b111111111;
assign micromatrizz[86][550] = 9'b111111111;
assign micromatrizz[86][551] = 9'b111111111;
assign micromatrizz[86][552] = 9'b111111111;
assign micromatrizz[86][553] = 9'b111111111;
assign micromatrizz[86][554] = 9'b111111111;
assign micromatrizz[86][555] = 9'b111111111;
assign micromatrizz[86][556] = 9'b111111111;
assign micromatrizz[86][557] = 9'b111111111;
assign micromatrizz[86][558] = 9'b111111111;
assign micromatrizz[86][559] = 9'b111111111;
assign micromatrizz[86][560] = 9'b111111111;
assign micromatrizz[86][561] = 9'b111111111;
assign micromatrizz[86][562] = 9'b111111111;
assign micromatrizz[86][563] = 9'b111111111;
assign micromatrizz[86][564] = 9'b111111111;
assign micromatrizz[86][565] = 9'b111111111;
assign micromatrizz[86][566] = 9'b111111111;
assign micromatrizz[86][567] = 9'b111111111;
assign micromatrizz[86][568] = 9'b111111111;
assign micromatrizz[86][569] = 9'b111111111;
assign micromatrizz[86][570] = 9'b111111111;
assign micromatrizz[86][571] = 9'b111111111;
assign micromatrizz[86][572] = 9'b111111111;
assign micromatrizz[86][573] = 9'b111111111;
assign micromatrizz[86][574] = 9'b111111111;
assign micromatrizz[86][575] = 9'b111111111;
assign micromatrizz[86][576] = 9'b111111111;
assign micromatrizz[86][577] = 9'b111111111;
assign micromatrizz[86][578] = 9'b111111111;
assign micromatrizz[86][579] = 9'b111111111;
assign micromatrizz[86][580] = 9'b111111111;
assign micromatrizz[86][581] = 9'b111111111;
assign micromatrizz[86][582] = 9'b111111111;
assign micromatrizz[86][583] = 9'b111111111;
assign micromatrizz[86][584] = 9'b111111111;
assign micromatrizz[86][585] = 9'b111111111;
assign micromatrizz[86][586] = 9'b111111111;
assign micromatrizz[86][587] = 9'b111111111;
assign micromatrizz[86][588] = 9'b111111111;
assign micromatrizz[86][589] = 9'b111111111;
assign micromatrizz[86][590] = 9'b111111111;
assign micromatrizz[86][591] = 9'b111111111;
assign micromatrizz[86][592] = 9'b111111111;
assign micromatrizz[86][593] = 9'b111111111;
assign micromatrizz[86][594] = 9'b111111111;
assign micromatrizz[86][595] = 9'b111111111;
assign micromatrizz[86][596] = 9'b111111111;
assign micromatrizz[86][597] = 9'b111111111;
assign micromatrizz[86][598] = 9'b111111111;
assign micromatrizz[86][599] = 9'b111111111;
assign micromatrizz[86][600] = 9'b111111111;
assign micromatrizz[86][601] = 9'b111111111;
assign micromatrizz[86][602] = 9'b111111111;
assign micromatrizz[86][603] = 9'b111111111;
assign micromatrizz[86][604] = 9'b111111111;
assign micromatrizz[86][605] = 9'b111111111;
assign micromatrizz[86][606] = 9'b111111111;
assign micromatrizz[86][607] = 9'b111111111;
assign micromatrizz[86][608] = 9'b111111111;
assign micromatrizz[86][609] = 9'b111111111;
assign micromatrizz[86][610] = 9'b111111111;
assign micromatrizz[86][611] = 9'b111111111;
assign micromatrizz[86][612] = 9'b111111111;
assign micromatrizz[86][613] = 9'b111111111;
assign micromatrizz[86][614] = 9'b111111111;
assign micromatrizz[86][615] = 9'b111111111;
assign micromatrizz[86][616] = 9'b111111111;
assign micromatrizz[86][617] = 9'b111111111;
assign micromatrizz[86][618] = 9'b111111111;
assign micromatrizz[86][619] = 9'b111111111;
assign micromatrizz[86][620] = 9'b111111111;
assign micromatrizz[86][621] = 9'b111111111;
assign micromatrizz[86][622] = 9'b111111111;
assign micromatrizz[86][623] = 9'b111111111;
assign micromatrizz[86][624] = 9'b111111111;
assign micromatrizz[86][625] = 9'b111111111;
assign micromatrizz[86][626] = 9'b111111111;
assign micromatrizz[86][627] = 9'b111111111;
assign micromatrizz[86][628] = 9'b111111111;
assign micromatrizz[86][629] = 9'b111111111;
assign micromatrizz[86][630] = 9'b111111111;
assign micromatrizz[86][631] = 9'b111111111;
assign micromatrizz[86][632] = 9'b111111111;
assign micromatrizz[86][633] = 9'b111111111;
assign micromatrizz[86][634] = 9'b111111111;
assign micromatrizz[86][635] = 9'b111111111;
assign micromatrizz[86][636] = 9'b111111111;
assign micromatrizz[86][637] = 9'b111111111;
assign micromatrizz[86][638] = 9'b111111111;
assign micromatrizz[86][639] = 9'b111111111;
assign micromatrizz[87][0] = 9'b111111111;
assign micromatrizz[87][1] = 9'b111111111;
assign micromatrizz[87][2] = 9'b111111111;
assign micromatrizz[87][3] = 9'b111111111;
assign micromatrizz[87][4] = 9'b111111111;
assign micromatrizz[87][5] = 9'b111111111;
assign micromatrizz[87][6] = 9'b111111111;
assign micromatrizz[87][7] = 9'b111111111;
assign micromatrizz[87][8] = 9'b111111111;
assign micromatrizz[87][9] = 9'b111111111;
assign micromatrizz[87][10] = 9'b111111111;
assign micromatrizz[87][11] = 9'b111111111;
assign micromatrizz[87][12] = 9'b111111111;
assign micromatrizz[87][13] = 9'b111111111;
assign micromatrizz[87][14] = 9'b111111111;
assign micromatrizz[87][15] = 9'b111111111;
assign micromatrizz[87][16] = 9'b111111111;
assign micromatrizz[87][17] = 9'b111111111;
assign micromatrizz[87][18] = 9'b111111111;
assign micromatrizz[87][19] = 9'b111111111;
assign micromatrizz[87][20] = 9'b111111111;
assign micromatrizz[87][21] = 9'b111111111;
assign micromatrizz[87][22] = 9'b111111111;
assign micromatrizz[87][23] = 9'b111111111;
assign micromatrizz[87][24] = 9'b111111111;
assign micromatrizz[87][25] = 9'b111111111;
assign micromatrizz[87][26] = 9'b111111111;
assign micromatrizz[87][27] = 9'b111111111;
assign micromatrizz[87][28] = 9'b111111111;
assign micromatrizz[87][29] = 9'b111111111;
assign micromatrizz[87][30] = 9'b111111111;
assign micromatrizz[87][31] = 9'b111111111;
assign micromatrizz[87][32] = 9'b111111111;
assign micromatrizz[87][33] = 9'b111111111;
assign micromatrizz[87][34] = 9'b111111111;
assign micromatrizz[87][35] = 9'b111111111;
assign micromatrizz[87][36] = 9'b111111111;
assign micromatrizz[87][37] = 9'b111111111;
assign micromatrizz[87][38] = 9'b111111111;
assign micromatrizz[87][39] = 9'b111111111;
assign micromatrizz[87][40] = 9'b111111111;
assign micromatrizz[87][41] = 9'b111111111;
assign micromatrizz[87][42] = 9'b111111111;
assign micromatrizz[87][43] = 9'b111111111;
assign micromatrizz[87][44] = 9'b111111111;
assign micromatrizz[87][45] = 9'b111111111;
assign micromatrizz[87][46] = 9'b111111111;
assign micromatrizz[87][47] = 9'b111111111;
assign micromatrizz[87][48] = 9'b111111111;
assign micromatrizz[87][49] = 9'b111111111;
assign micromatrizz[87][50] = 9'b111111111;
assign micromatrizz[87][51] = 9'b111111111;
assign micromatrizz[87][52] = 9'b111111111;
assign micromatrizz[87][53] = 9'b111111111;
assign micromatrizz[87][54] = 9'b111111111;
assign micromatrizz[87][55] = 9'b111111111;
assign micromatrizz[87][56] = 9'b111111111;
assign micromatrizz[87][57] = 9'b111111111;
assign micromatrizz[87][58] = 9'b111111111;
assign micromatrizz[87][59] = 9'b111111111;
assign micromatrizz[87][60] = 9'b111111111;
assign micromatrizz[87][61] = 9'b111111111;
assign micromatrizz[87][62] = 9'b111111111;
assign micromatrizz[87][63] = 9'b111111111;
assign micromatrizz[87][64] = 9'b111111111;
assign micromatrizz[87][65] = 9'b111111111;
assign micromatrizz[87][66] = 9'b111111111;
assign micromatrizz[87][67] = 9'b111111111;
assign micromatrizz[87][68] = 9'b111111111;
assign micromatrizz[87][69] = 9'b111111111;
assign micromatrizz[87][70] = 9'b111111111;
assign micromatrizz[87][71] = 9'b111111111;
assign micromatrizz[87][72] = 9'b111111111;
assign micromatrizz[87][73] = 9'b111111111;
assign micromatrizz[87][74] = 9'b111111111;
assign micromatrizz[87][75] = 9'b111111111;
assign micromatrizz[87][76] = 9'b111111111;
assign micromatrizz[87][77] = 9'b111111111;
assign micromatrizz[87][78] = 9'b111111111;
assign micromatrizz[87][79] = 9'b111111111;
assign micromatrizz[87][80] = 9'b111111111;
assign micromatrizz[87][81] = 9'b111111111;
assign micromatrizz[87][82] = 9'b111111111;
assign micromatrizz[87][83] = 9'b111111111;
assign micromatrizz[87][84] = 9'b111111111;
assign micromatrizz[87][85] = 9'b111111111;
assign micromatrizz[87][86] = 9'b111111111;
assign micromatrizz[87][87] = 9'b111111111;
assign micromatrizz[87][88] = 9'b111111111;
assign micromatrizz[87][89] = 9'b111111111;
assign micromatrizz[87][90] = 9'b111111111;
assign micromatrizz[87][91] = 9'b111111111;
assign micromatrizz[87][92] = 9'b111111111;
assign micromatrizz[87][93] = 9'b111111111;
assign micromatrizz[87][94] = 9'b111111111;
assign micromatrizz[87][95] = 9'b111111111;
assign micromatrizz[87][96] = 9'b111111111;
assign micromatrizz[87][97] = 9'b111111111;
assign micromatrizz[87][98] = 9'b111111111;
assign micromatrizz[87][99] = 9'b111111111;
assign micromatrizz[87][100] = 9'b111111111;
assign micromatrizz[87][101] = 9'b111111111;
assign micromatrizz[87][102] = 9'b111111111;
assign micromatrizz[87][103] = 9'b111111111;
assign micromatrizz[87][104] = 9'b111111111;
assign micromatrizz[87][105] = 9'b111111111;
assign micromatrizz[87][106] = 9'b111111111;
assign micromatrizz[87][107] = 9'b111111111;
assign micromatrizz[87][108] = 9'b111111111;
assign micromatrizz[87][109] = 9'b111111111;
assign micromatrizz[87][110] = 9'b111111111;
assign micromatrizz[87][111] = 9'b111111111;
assign micromatrizz[87][112] = 9'b111111111;
assign micromatrizz[87][113] = 9'b111111111;
assign micromatrizz[87][114] = 9'b111111111;
assign micromatrizz[87][115] = 9'b111111111;
assign micromatrizz[87][116] = 9'b111111111;
assign micromatrizz[87][117] = 9'b111111111;
assign micromatrizz[87][118] = 9'b111111111;
assign micromatrizz[87][119] = 9'b111111111;
assign micromatrizz[87][120] = 9'b111111111;
assign micromatrizz[87][121] = 9'b111111111;
assign micromatrizz[87][122] = 9'b111111111;
assign micromatrizz[87][123] = 9'b111111111;
assign micromatrizz[87][124] = 9'b111111111;
assign micromatrizz[87][125] = 9'b111111111;
assign micromatrizz[87][126] = 9'b111111111;
assign micromatrizz[87][127] = 9'b111111111;
assign micromatrizz[87][128] = 9'b111111111;
assign micromatrizz[87][129] = 9'b111111111;
assign micromatrizz[87][130] = 9'b111111111;
assign micromatrizz[87][131] = 9'b111111111;
assign micromatrizz[87][132] = 9'b111111111;
assign micromatrizz[87][133] = 9'b111111111;
assign micromatrizz[87][134] = 9'b111111111;
assign micromatrizz[87][135] = 9'b111111111;
assign micromatrizz[87][136] = 9'b111111111;
assign micromatrizz[87][137] = 9'b111111111;
assign micromatrizz[87][138] = 9'b111111111;
assign micromatrizz[87][139] = 9'b111111111;
assign micromatrizz[87][140] = 9'b111111111;
assign micromatrizz[87][141] = 9'b111111111;
assign micromatrizz[87][142] = 9'b111111111;
assign micromatrizz[87][143] = 9'b111111111;
assign micromatrizz[87][144] = 9'b111111111;
assign micromatrizz[87][145] = 9'b111111111;
assign micromatrizz[87][146] = 9'b111111111;
assign micromatrizz[87][147] = 9'b111111111;
assign micromatrizz[87][148] = 9'b111111111;
assign micromatrizz[87][149] = 9'b111111111;
assign micromatrizz[87][150] = 9'b111111111;
assign micromatrizz[87][151] = 9'b111111111;
assign micromatrizz[87][152] = 9'b111111111;
assign micromatrizz[87][153] = 9'b111111111;
assign micromatrizz[87][154] = 9'b111111111;
assign micromatrizz[87][155] = 9'b111111111;
assign micromatrizz[87][156] = 9'b111111111;
assign micromatrizz[87][157] = 9'b111111111;
assign micromatrizz[87][158] = 9'b111111111;
assign micromatrizz[87][159] = 9'b111111111;
assign micromatrizz[87][160] = 9'b111111111;
assign micromatrizz[87][161] = 9'b111111111;
assign micromatrizz[87][162] = 9'b111111111;
assign micromatrizz[87][163] = 9'b111111111;
assign micromatrizz[87][164] = 9'b111111111;
assign micromatrizz[87][165] = 9'b111111111;
assign micromatrizz[87][166] = 9'b111111111;
assign micromatrizz[87][167] = 9'b111111111;
assign micromatrizz[87][168] = 9'b111111111;
assign micromatrizz[87][169] = 9'b111111111;
assign micromatrizz[87][170] = 9'b111111111;
assign micromatrizz[87][171] = 9'b111111111;
assign micromatrizz[87][172] = 9'b111111111;
assign micromatrizz[87][173] = 9'b111111111;
assign micromatrizz[87][174] = 9'b111111111;
assign micromatrizz[87][175] = 9'b111111111;
assign micromatrizz[87][176] = 9'b111111111;
assign micromatrizz[87][177] = 9'b111111111;
assign micromatrizz[87][178] = 9'b111111111;
assign micromatrizz[87][179] = 9'b111111111;
assign micromatrizz[87][180] = 9'b111111111;
assign micromatrizz[87][181] = 9'b111111111;
assign micromatrizz[87][182] = 9'b111111111;
assign micromatrizz[87][183] = 9'b111111111;
assign micromatrizz[87][184] = 9'b111111111;
assign micromatrizz[87][185] = 9'b111111111;
assign micromatrizz[87][186] = 9'b111111111;
assign micromatrizz[87][187] = 9'b111111111;
assign micromatrizz[87][188] = 9'b111111111;
assign micromatrizz[87][189] = 9'b111111111;
assign micromatrizz[87][190] = 9'b111111111;
assign micromatrizz[87][191] = 9'b111111111;
assign micromatrizz[87][192] = 9'b111111111;
assign micromatrizz[87][193] = 9'b111111111;
assign micromatrizz[87][194] = 9'b111111111;
assign micromatrizz[87][195] = 9'b111111111;
assign micromatrizz[87][196] = 9'b111111111;
assign micromatrizz[87][197] = 9'b111111111;
assign micromatrizz[87][198] = 9'b111111111;
assign micromatrizz[87][199] = 9'b111111111;
assign micromatrizz[87][200] = 9'b111111111;
assign micromatrizz[87][201] = 9'b111111111;
assign micromatrizz[87][202] = 9'b111111111;
assign micromatrizz[87][203] = 9'b111111111;
assign micromatrizz[87][204] = 9'b111111111;
assign micromatrizz[87][205] = 9'b111111111;
assign micromatrizz[87][206] = 9'b111111111;
assign micromatrizz[87][207] = 9'b111111111;
assign micromatrizz[87][208] = 9'b111111111;
assign micromatrizz[87][209] = 9'b111111111;
assign micromatrizz[87][210] = 9'b111111111;
assign micromatrizz[87][211] = 9'b111111111;
assign micromatrizz[87][212] = 9'b111111111;
assign micromatrizz[87][213] = 9'b111111111;
assign micromatrizz[87][214] = 9'b111111111;
assign micromatrizz[87][215] = 9'b111111111;
assign micromatrizz[87][216] = 9'b111111111;
assign micromatrizz[87][217] = 9'b111111111;
assign micromatrizz[87][218] = 9'b111111111;
assign micromatrizz[87][219] = 9'b111111111;
assign micromatrizz[87][220] = 9'b111111111;
assign micromatrizz[87][221] = 9'b111111111;
assign micromatrizz[87][222] = 9'b111111111;
assign micromatrizz[87][223] = 9'b111111111;
assign micromatrizz[87][224] = 9'b111111111;
assign micromatrizz[87][225] = 9'b111111111;
assign micromatrizz[87][226] = 9'b111111111;
assign micromatrizz[87][227] = 9'b111111111;
assign micromatrizz[87][228] = 9'b111111111;
assign micromatrizz[87][229] = 9'b111111111;
assign micromatrizz[87][230] = 9'b111111111;
assign micromatrizz[87][231] = 9'b111111111;
assign micromatrizz[87][232] = 9'b111111111;
assign micromatrizz[87][233] = 9'b111111111;
assign micromatrizz[87][234] = 9'b111111111;
assign micromatrizz[87][235] = 9'b111111111;
assign micromatrizz[87][236] = 9'b111111111;
assign micromatrizz[87][237] = 9'b111111111;
assign micromatrizz[87][238] = 9'b111111111;
assign micromatrizz[87][239] = 9'b111111111;
assign micromatrizz[87][240] = 9'b111111111;
assign micromatrizz[87][241] = 9'b111111111;
assign micromatrizz[87][242] = 9'b111111111;
assign micromatrizz[87][243] = 9'b111111111;
assign micromatrizz[87][244] = 9'b111111111;
assign micromatrizz[87][245] = 9'b111111111;
assign micromatrizz[87][246] = 9'b111111111;
assign micromatrizz[87][247] = 9'b111111111;
assign micromatrizz[87][248] = 9'b111111111;
assign micromatrizz[87][249] = 9'b111111111;
assign micromatrizz[87][250] = 9'b111111111;
assign micromatrizz[87][251] = 9'b111111111;
assign micromatrizz[87][252] = 9'b111111111;
assign micromatrizz[87][253] = 9'b111111111;
assign micromatrizz[87][254] = 9'b111111111;
assign micromatrizz[87][255] = 9'b111111111;
assign micromatrizz[87][256] = 9'b111111111;
assign micromatrizz[87][257] = 9'b111111111;
assign micromatrizz[87][258] = 9'b111111111;
assign micromatrizz[87][259] = 9'b111111111;
assign micromatrizz[87][260] = 9'b111111111;
assign micromatrizz[87][261] = 9'b111111111;
assign micromatrizz[87][262] = 9'b111111111;
assign micromatrizz[87][263] = 9'b111111111;
assign micromatrizz[87][264] = 9'b111111111;
assign micromatrizz[87][265] = 9'b111111111;
assign micromatrizz[87][266] = 9'b111111111;
assign micromatrizz[87][267] = 9'b111111111;
assign micromatrizz[87][268] = 9'b111111111;
assign micromatrizz[87][269] = 9'b111111111;
assign micromatrizz[87][270] = 9'b111111111;
assign micromatrizz[87][271] = 9'b111111111;
assign micromatrizz[87][272] = 9'b111111111;
assign micromatrizz[87][273] = 9'b111111111;
assign micromatrizz[87][274] = 9'b111111111;
assign micromatrizz[87][275] = 9'b111111111;
assign micromatrizz[87][276] = 9'b111111111;
assign micromatrizz[87][277] = 9'b111111111;
assign micromatrizz[87][278] = 9'b111111111;
assign micromatrizz[87][279] = 9'b111111111;
assign micromatrizz[87][280] = 9'b111111111;
assign micromatrizz[87][281] = 9'b111111111;
assign micromatrizz[87][282] = 9'b111111111;
assign micromatrizz[87][283] = 9'b111111111;
assign micromatrizz[87][284] = 9'b111111111;
assign micromatrizz[87][285] = 9'b111111111;
assign micromatrizz[87][286] = 9'b111111111;
assign micromatrizz[87][287] = 9'b111111111;
assign micromatrizz[87][288] = 9'b111111111;
assign micromatrizz[87][289] = 9'b111111111;
assign micromatrizz[87][290] = 9'b111111111;
assign micromatrizz[87][291] = 9'b111111111;
assign micromatrizz[87][292] = 9'b111111111;
assign micromatrizz[87][293] = 9'b111111111;
assign micromatrizz[87][294] = 9'b111111111;
assign micromatrizz[87][295] = 9'b111111111;
assign micromatrizz[87][296] = 9'b111111111;
assign micromatrizz[87][297] = 9'b111111111;
assign micromatrizz[87][298] = 9'b111111111;
assign micromatrizz[87][299] = 9'b111111111;
assign micromatrizz[87][300] = 9'b111111111;
assign micromatrizz[87][301] = 9'b111111111;
assign micromatrizz[87][302] = 9'b111111111;
assign micromatrizz[87][303] = 9'b111111111;
assign micromatrizz[87][304] = 9'b111111111;
assign micromatrizz[87][305] = 9'b111111111;
assign micromatrizz[87][306] = 9'b111111111;
assign micromatrizz[87][307] = 9'b111111111;
assign micromatrizz[87][308] = 9'b111111111;
assign micromatrizz[87][309] = 9'b111111111;
assign micromatrizz[87][310] = 9'b111111111;
assign micromatrizz[87][311] = 9'b111111111;
assign micromatrizz[87][312] = 9'b111111111;
assign micromatrizz[87][313] = 9'b111111111;
assign micromatrizz[87][314] = 9'b111111111;
assign micromatrizz[87][315] = 9'b111111111;
assign micromatrizz[87][316] = 9'b111111111;
assign micromatrizz[87][317] = 9'b111111111;
assign micromatrizz[87][318] = 9'b111111111;
assign micromatrizz[87][319] = 9'b111111111;
assign micromatrizz[87][320] = 9'b111111111;
assign micromatrizz[87][321] = 9'b111111111;
assign micromatrizz[87][322] = 9'b111111111;
assign micromatrizz[87][323] = 9'b111111111;
assign micromatrizz[87][324] = 9'b111111111;
assign micromatrizz[87][325] = 9'b111111111;
assign micromatrizz[87][326] = 9'b111111111;
assign micromatrizz[87][327] = 9'b111111111;
assign micromatrizz[87][328] = 9'b111111111;
assign micromatrizz[87][329] = 9'b111111111;
assign micromatrizz[87][330] = 9'b111111111;
assign micromatrizz[87][331] = 9'b111111111;
assign micromatrizz[87][332] = 9'b111111111;
assign micromatrizz[87][333] = 9'b111111111;
assign micromatrizz[87][334] = 9'b111111111;
assign micromatrizz[87][335] = 9'b111111111;
assign micromatrizz[87][336] = 9'b111111111;
assign micromatrizz[87][337] = 9'b111111111;
assign micromatrizz[87][338] = 9'b111111111;
assign micromatrizz[87][339] = 9'b111111111;
assign micromatrizz[87][340] = 9'b111111111;
assign micromatrizz[87][341] = 9'b111111111;
assign micromatrizz[87][342] = 9'b111111111;
assign micromatrizz[87][343] = 9'b111111111;
assign micromatrizz[87][344] = 9'b111111111;
assign micromatrizz[87][345] = 9'b111111111;
assign micromatrizz[87][346] = 9'b111111111;
assign micromatrizz[87][347] = 9'b111111111;
assign micromatrizz[87][348] = 9'b111111111;
assign micromatrizz[87][349] = 9'b111111111;
assign micromatrizz[87][350] = 9'b111111111;
assign micromatrizz[87][351] = 9'b111111111;
assign micromatrizz[87][352] = 9'b111111111;
assign micromatrizz[87][353] = 9'b111111111;
assign micromatrizz[87][354] = 9'b111111111;
assign micromatrizz[87][355] = 9'b111111111;
assign micromatrizz[87][356] = 9'b111111111;
assign micromatrizz[87][357] = 9'b111111111;
assign micromatrizz[87][358] = 9'b111111111;
assign micromatrizz[87][359] = 9'b111111111;
assign micromatrizz[87][360] = 9'b111111111;
assign micromatrizz[87][361] = 9'b111111111;
assign micromatrizz[87][362] = 9'b111111111;
assign micromatrizz[87][363] = 9'b111111111;
assign micromatrizz[87][364] = 9'b111111111;
assign micromatrizz[87][365] = 9'b111111111;
assign micromatrizz[87][366] = 9'b111111111;
assign micromatrizz[87][367] = 9'b111111111;
assign micromatrizz[87][368] = 9'b111111111;
assign micromatrizz[87][369] = 9'b111111111;
assign micromatrizz[87][370] = 9'b111111111;
assign micromatrizz[87][371] = 9'b111111111;
assign micromatrizz[87][372] = 9'b111111111;
assign micromatrizz[87][373] = 9'b111111111;
assign micromatrizz[87][374] = 9'b111111111;
assign micromatrizz[87][375] = 9'b111111111;
assign micromatrizz[87][376] = 9'b111111111;
assign micromatrizz[87][377] = 9'b111111111;
assign micromatrizz[87][378] = 9'b111111111;
assign micromatrizz[87][379] = 9'b111111111;
assign micromatrizz[87][380] = 9'b111111111;
assign micromatrizz[87][381] = 9'b111111111;
assign micromatrizz[87][382] = 9'b111111111;
assign micromatrizz[87][383] = 9'b111111111;
assign micromatrizz[87][384] = 9'b111111111;
assign micromatrizz[87][385] = 9'b111111111;
assign micromatrizz[87][386] = 9'b111111111;
assign micromatrizz[87][387] = 9'b111111111;
assign micromatrizz[87][388] = 9'b111111111;
assign micromatrizz[87][389] = 9'b111111111;
assign micromatrizz[87][390] = 9'b111111111;
assign micromatrizz[87][391] = 9'b111111111;
assign micromatrizz[87][392] = 9'b111111111;
assign micromatrizz[87][393] = 9'b111111111;
assign micromatrizz[87][394] = 9'b111111111;
assign micromatrizz[87][395] = 9'b111111111;
assign micromatrizz[87][396] = 9'b111111111;
assign micromatrizz[87][397] = 9'b111111111;
assign micromatrizz[87][398] = 9'b111111111;
assign micromatrizz[87][399] = 9'b111111111;
assign micromatrizz[87][400] = 9'b111111111;
assign micromatrizz[87][401] = 9'b111111111;
assign micromatrizz[87][402] = 9'b111111111;
assign micromatrizz[87][403] = 9'b111111111;
assign micromatrizz[87][404] = 9'b111111111;
assign micromatrizz[87][405] = 9'b111111111;
assign micromatrizz[87][406] = 9'b111111111;
assign micromatrizz[87][407] = 9'b111111111;
assign micromatrizz[87][408] = 9'b111111111;
assign micromatrizz[87][409] = 9'b111111111;
assign micromatrizz[87][410] = 9'b111111111;
assign micromatrizz[87][411] = 9'b111111111;
assign micromatrizz[87][412] = 9'b111111111;
assign micromatrizz[87][413] = 9'b111111111;
assign micromatrizz[87][414] = 9'b111111111;
assign micromatrizz[87][415] = 9'b111111111;
assign micromatrizz[87][416] = 9'b111111111;
assign micromatrizz[87][417] = 9'b111111111;
assign micromatrizz[87][418] = 9'b111111111;
assign micromatrizz[87][419] = 9'b111111111;
assign micromatrizz[87][420] = 9'b111111111;
assign micromatrizz[87][421] = 9'b111111111;
assign micromatrizz[87][422] = 9'b111111111;
assign micromatrizz[87][423] = 9'b111111111;
assign micromatrizz[87][424] = 9'b111111111;
assign micromatrizz[87][425] = 9'b111111111;
assign micromatrizz[87][426] = 9'b111111111;
assign micromatrizz[87][427] = 9'b111111111;
assign micromatrizz[87][428] = 9'b111111111;
assign micromatrizz[87][429] = 9'b111111111;
assign micromatrizz[87][430] = 9'b111111111;
assign micromatrizz[87][431] = 9'b111111111;
assign micromatrizz[87][432] = 9'b111111111;
assign micromatrizz[87][433] = 9'b111111111;
assign micromatrizz[87][434] = 9'b111111111;
assign micromatrizz[87][435] = 9'b111111111;
assign micromatrizz[87][436] = 9'b111111111;
assign micromatrizz[87][437] = 9'b111111111;
assign micromatrizz[87][438] = 9'b111111111;
assign micromatrizz[87][439] = 9'b111111111;
assign micromatrizz[87][440] = 9'b111111111;
assign micromatrizz[87][441] = 9'b111111111;
assign micromatrizz[87][442] = 9'b111111111;
assign micromatrizz[87][443] = 9'b111111111;
assign micromatrizz[87][444] = 9'b111111111;
assign micromatrizz[87][445] = 9'b111111111;
assign micromatrizz[87][446] = 9'b111111111;
assign micromatrizz[87][447] = 9'b111111111;
assign micromatrizz[87][448] = 9'b111111111;
assign micromatrizz[87][449] = 9'b111111111;
assign micromatrizz[87][450] = 9'b111111111;
assign micromatrizz[87][451] = 9'b111111111;
assign micromatrizz[87][452] = 9'b111111111;
assign micromatrizz[87][453] = 9'b111111111;
assign micromatrizz[87][454] = 9'b111111111;
assign micromatrizz[87][455] = 9'b111111111;
assign micromatrizz[87][456] = 9'b111111111;
assign micromatrizz[87][457] = 9'b111111111;
assign micromatrizz[87][458] = 9'b111111111;
assign micromatrizz[87][459] = 9'b111111111;
assign micromatrizz[87][460] = 9'b111111111;
assign micromatrizz[87][461] = 9'b111111111;
assign micromatrizz[87][462] = 9'b111111111;
assign micromatrizz[87][463] = 9'b111111111;
assign micromatrizz[87][464] = 9'b111111111;
assign micromatrizz[87][465] = 9'b111111111;
assign micromatrizz[87][466] = 9'b111111111;
assign micromatrizz[87][467] = 9'b111111111;
assign micromatrizz[87][468] = 9'b111111111;
assign micromatrizz[87][469] = 9'b111111111;
assign micromatrizz[87][470] = 9'b111111111;
assign micromatrizz[87][471] = 9'b111111111;
assign micromatrizz[87][472] = 9'b111111111;
assign micromatrizz[87][473] = 9'b111111111;
assign micromatrizz[87][474] = 9'b111111111;
assign micromatrizz[87][475] = 9'b111111111;
assign micromatrizz[87][476] = 9'b111111111;
assign micromatrizz[87][477] = 9'b111111111;
assign micromatrizz[87][478] = 9'b111111111;
assign micromatrizz[87][479] = 9'b111111111;
assign micromatrizz[87][480] = 9'b111111111;
assign micromatrizz[87][481] = 9'b111111111;
assign micromatrizz[87][482] = 9'b111111111;
assign micromatrizz[87][483] = 9'b111111111;
assign micromatrizz[87][484] = 9'b111111111;
assign micromatrizz[87][485] = 9'b111111111;
assign micromatrizz[87][486] = 9'b111111111;
assign micromatrizz[87][487] = 9'b111111111;
assign micromatrizz[87][488] = 9'b111111111;
assign micromatrizz[87][489] = 9'b111111111;
assign micromatrizz[87][490] = 9'b111111111;
assign micromatrizz[87][491] = 9'b111111111;
assign micromatrizz[87][492] = 9'b111111111;
assign micromatrizz[87][493] = 9'b111111111;
assign micromatrizz[87][494] = 9'b111111111;
assign micromatrizz[87][495] = 9'b111111111;
assign micromatrizz[87][496] = 9'b111111111;
assign micromatrizz[87][497] = 9'b111111111;
assign micromatrizz[87][498] = 9'b111111111;
assign micromatrizz[87][499] = 9'b111111111;
assign micromatrizz[87][500] = 9'b111111111;
assign micromatrizz[87][501] = 9'b111111111;
assign micromatrizz[87][502] = 9'b111111111;
assign micromatrizz[87][503] = 9'b111111111;
assign micromatrizz[87][504] = 9'b111111111;
assign micromatrizz[87][505] = 9'b111111111;
assign micromatrizz[87][506] = 9'b111111111;
assign micromatrizz[87][507] = 9'b111111111;
assign micromatrizz[87][508] = 9'b111111111;
assign micromatrizz[87][509] = 9'b111111111;
assign micromatrizz[87][510] = 9'b111111111;
assign micromatrizz[87][511] = 9'b111111111;
assign micromatrizz[87][512] = 9'b111111111;
assign micromatrizz[87][513] = 9'b111111111;
assign micromatrizz[87][514] = 9'b111111111;
assign micromatrizz[87][515] = 9'b111111111;
assign micromatrizz[87][516] = 9'b111111111;
assign micromatrizz[87][517] = 9'b111111111;
assign micromatrizz[87][518] = 9'b111111111;
assign micromatrizz[87][519] = 9'b111111111;
assign micromatrizz[87][520] = 9'b111111111;
assign micromatrizz[87][521] = 9'b111111111;
assign micromatrizz[87][522] = 9'b111111111;
assign micromatrizz[87][523] = 9'b111111111;
assign micromatrizz[87][524] = 9'b111111111;
assign micromatrizz[87][525] = 9'b111111111;
assign micromatrizz[87][526] = 9'b111111111;
assign micromatrizz[87][527] = 9'b111111111;
assign micromatrizz[87][528] = 9'b111111111;
assign micromatrizz[87][529] = 9'b111111111;
assign micromatrizz[87][530] = 9'b111111111;
assign micromatrizz[87][531] = 9'b111111111;
assign micromatrizz[87][532] = 9'b111111111;
assign micromatrizz[87][533] = 9'b111111111;
assign micromatrizz[87][534] = 9'b111111111;
assign micromatrizz[87][535] = 9'b111111111;
assign micromatrizz[87][536] = 9'b111111111;
assign micromatrizz[87][537] = 9'b111111111;
assign micromatrizz[87][538] = 9'b111111111;
assign micromatrizz[87][539] = 9'b111111111;
assign micromatrizz[87][540] = 9'b111111111;
assign micromatrizz[87][541] = 9'b111111111;
assign micromatrizz[87][542] = 9'b111111111;
assign micromatrizz[87][543] = 9'b111111111;
assign micromatrizz[87][544] = 9'b111111111;
assign micromatrizz[87][545] = 9'b111111111;
assign micromatrizz[87][546] = 9'b111111111;
assign micromatrizz[87][547] = 9'b111111111;
assign micromatrizz[87][548] = 9'b111111111;
assign micromatrizz[87][549] = 9'b111111111;
assign micromatrizz[87][550] = 9'b111111111;
assign micromatrizz[87][551] = 9'b111111111;
assign micromatrizz[87][552] = 9'b111111111;
assign micromatrizz[87][553] = 9'b111111111;
assign micromatrizz[87][554] = 9'b111111111;
assign micromatrizz[87][555] = 9'b111111111;
assign micromatrizz[87][556] = 9'b111111111;
assign micromatrizz[87][557] = 9'b111111111;
assign micromatrizz[87][558] = 9'b111111111;
assign micromatrizz[87][559] = 9'b111111111;
assign micromatrizz[87][560] = 9'b111111111;
assign micromatrizz[87][561] = 9'b111111111;
assign micromatrizz[87][562] = 9'b111111111;
assign micromatrizz[87][563] = 9'b111111111;
assign micromatrizz[87][564] = 9'b111111111;
assign micromatrizz[87][565] = 9'b111111111;
assign micromatrizz[87][566] = 9'b111111111;
assign micromatrizz[87][567] = 9'b111111111;
assign micromatrizz[87][568] = 9'b111111111;
assign micromatrizz[87][569] = 9'b111111111;
assign micromatrizz[87][570] = 9'b111111111;
assign micromatrizz[87][571] = 9'b111111111;
assign micromatrizz[87][572] = 9'b111111111;
assign micromatrizz[87][573] = 9'b111111111;
assign micromatrizz[87][574] = 9'b111111111;
assign micromatrizz[87][575] = 9'b111111111;
assign micromatrizz[87][576] = 9'b111111111;
assign micromatrizz[87][577] = 9'b111111111;
assign micromatrizz[87][578] = 9'b111111111;
assign micromatrizz[87][579] = 9'b111111111;
assign micromatrizz[87][580] = 9'b111111111;
assign micromatrizz[87][581] = 9'b111111111;
assign micromatrizz[87][582] = 9'b111111111;
assign micromatrizz[87][583] = 9'b111111111;
assign micromatrizz[87][584] = 9'b111111111;
assign micromatrizz[87][585] = 9'b111111111;
assign micromatrizz[87][586] = 9'b111111111;
assign micromatrizz[87][587] = 9'b111111111;
assign micromatrizz[87][588] = 9'b111111111;
assign micromatrizz[87][589] = 9'b111111111;
assign micromatrizz[87][590] = 9'b111111111;
assign micromatrizz[87][591] = 9'b111111111;
assign micromatrizz[87][592] = 9'b111111111;
assign micromatrizz[87][593] = 9'b111111111;
assign micromatrizz[87][594] = 9'b111111111;
assign micromatrizz[87][595] = 9'b111111111;
assign micromatrizz[87][596] = 9'b111111111;
assign micromatrizz[87][597] = 9'b111111111;
assign micromatrizz[87][598] = 9'b111111111;
assign micromatrizz[87][599] = 9'b111111111;
assign micromatrizz[87][600] = 9'b111111111;
assign micromatrizz[87][601] = 9'b111111111;
assign micromatrizz[87][602] = 9'b111111111;
assign micromatrizz[87][603] = 9'b111111111;
assign micromatrizz[87][604] = 9'b111111111;
assign micromatrizz[87][605] = 9'b111111111;
assign micromatrizz[87][606] = 9'b111111111;
assign micromatrizz[87][607] = 9'b111111111;
assign micromatrizz[87][608] = 9'b111111111;
assign micromatrizz[87][609] = 9'b111111111;
assign micromatrizz[87][610] = 9'b111111111;
assign micromatrizz[87][611] = 9'b111111111;
assign micromatrizz[87][612] = 9'b111111111;
assign micromatrizz[87][613] = 9'b111111111;
assign micromatrizz[87][614] = 9'b111111111;
assign micromatrizz[87][615] = 9'b111111111;
assign micromatrizz[87][616] = 9'b111111111;
assign micromatrizz[87][617] = 9'b111111111;
assign micromatrizz[87][618] = 9'b111111111;
assign micromatrizz[87][619] = 9'b111111111;
assign micromatrizz[87][620] = 9'b111111111;
assign micromatrizz[87][621] = 9'b111111111;
assign micromatrizz[87][622] = 9'b111111111;
assign micromatrizz[87][623] = 9'b111111111;
assign micromatrizz[87][624] = 9'b111111111;
assign micromatrizz[87][625] = 9'b111111111;
assign micromatrizz[87][626] = 9'b111111111;
assign micromatrizz[87][627] = 9'b111111111;
assign micromatrizz[87][628] = 9'b111111111;
assign micromatrizz[87][629] = 9'b111111111;
assign micromatrizz[87][630] = 9'b111111111;
assign micromatrizz[87][631] = 9'b111111111;
assign micromatrizz[87][632] = 9'b111111111;
assign micromatrizz[87][633] = 9'b111111111;
assign micromatrizz[87][634] = 9'b111111111;
assign micromatrizz[87][635] = 9'b111111111;
assign micromatrizz[87][636] = 9'b111111111;
assign micromatrizz[87][637] = 9'b111111111;
assign micromatrizz[87][638] = 9'b111111111;
assign micromatrizz[87][639] = 9'b111111111;
assign micromatrizz[88][0] = 9'b111111111;
assign micromatrizz[88][1] = 9'b111111111;
assign micromatrizz[88][2] = 9'b111111111;
assign micromatrizz[88][3] = 9'b111111111;
assign micromatrizz[88][4] = 9'b111111111;
assign micromatrizz[88][5] = 9'b111111111;
assign micromatrizz[88][6] = 9'b111111111;
assign micromatrizz[88][7] = 9'b111111111;
assign micromatrizz[88][8] = 9'b111111111;
assign micromatrizz[88][9] = 9'b111111111;
assign micromatrizz[88][10] = 9'b111111111;
assign micromatrizz[88][11] = 9'b111111111;
assign micromatrizz[88][12] = 9'b111111111;
assign micromatrizz[88][13] = 9'b111111111;
assign micromatrizz[88][14] = 9'b111111111;
assign micromatrizz[88][15] = 9'b111111111;
assign micromatrizz[88][16] = 9'b111111111;
assign micromatrizz[88][17] = 9'b111111111;
assign micromatrizz[88][18] = 9'b111111111;
assign micromatrizz[88][19] = 9'b111111111;
assign micromatrizz[88][20] = 9'b111111111;
assign micromatrizz[88][21] = 9'b111111111;
assign micromatrizz[88][22] = 9'b111111111;
assign micromatrizz[88][23] = 9'b111111111;
assign micromatrizz[88][24] = 9'b111111111;
assign micromatrizz[88][25] = 9'b111111111;
assign micromatrizz[88][26] = 9'b111111111;
assign micromatrizz[88][27] = 9'b111111111;
assign micromatrizz[88][28] = 9'b111111111;
assign micromatrizz[88][29] = 9'b111111111;
assign micromatrizz[88][30] = 9'b111111111;
assign micromatrizz[88][31] = 9'b111111111;
assign micromatrizz[88][32] = 9'b111111111;
assign micromatrizz[88][33] = 9'b111111111;
assign micromatrizz[88][34] = 9'b111111111;
assign micromatrizz[88][35] = 9'b111111111;
assign micromatrizz[88][36] = 9'b111111111;
assign micromatrizz[88][37] = 9'b111111111;
assign micromatrizz[88][38] = 9'b111111111;
assign micromatrizz[88][39] = 9'b111111111;
assign micromatrizz[88][40] = 9'b111111111;
assign micromatrizz[88][41] = 9'b111111111;
assign micromatrizz[88][42] = 9'b111111111;
assign micromatrizz[88][43] = 9'b111111111;
assign micromatrizz[88][44] = 9'b111111111;
assign micromatrizz[88][45] = 9'b111111111;
assign micromatrizz[88][46] = 9'b111111111;
assign micromatrizz[88][47] = 9'b111111111;
assign micromatrizz[88][48] = 9'b111111111;
assign micromatrizz[88][49] = 9'b111111111;
assign micromatrizz[88][50] = 9'b111111111;
assign micromatrizz[88][51] = 9'b111111111;
assign micromatrizz[88][52] = 9'b111111111;
assign micromatrizz[88][53] = 9'b111111111;
assign micromatrizz[88][54] = 9'b111111111;
assign micromatrizz[88][55] = 9'b111111111;
assign micromatrizz[88][56] = 9'b111111111;
assign micromatrizz[88][57] = 9'b111111111;
assign micromatrizz[88][58] = 9'b111111111;
assign micromatrizz[88][59] = 9'b111111111;
assign micromatrizz[88][60] = 9'b111111111;
assign micromatrizz[88][61] = 9'b111111111;
assign micromatrizz[88][62] = 9'b111111111;
assign micromatrizz[88][63] = 9'b111111111;
assign micromatrizz[88][64] = 9'b111111111;
assign micromatrizz[88][65] = 9'b111111111;
assign micromatrizz[88][66] = 9'b111111111;
assign micromatrizz[88][67] = 9'b111111111;
assign micromatrizz[88][68] = 9'b111111111;
assign micromatrizz[88][69] = 9'b111111111;
assign micromatrizz[88][70] = 9'b111111111;
assign micromatrizz[88][71] = 9'b111111111;
assign micromatrizz[88][72] = 9'b111111111;
assign micromatrizz[88][73] = 9'b111111111;
assign micromatrizz[88][74] = 9'b111111111;
assign micromatrizz[88][75] = 9'b111111111;
assign micromatrizz[88][76] = 9'b111111111;
assign micromatrizz[88][77] = 9'b111111111;
assign micromatrizz[88][78] = 9'b111111111;
assign micromatrizz[88][79] = 9'b111111111;
assign micromatrizz[88][80] = 9'b111111111;
assign micromatrizz[88][81] = 9'b111111111;
assign micromatrizz[88][82] = 9'b111111111;
assign micromatrizz[88][83] = 9'b111111111;
assign micromatrizz[88][84] = 9'b111111111;
assign micromatrizz[88][85] = 9'b111111111;
assign micromatrizz[88][86] = 9'b111111111;
assign micromatrizz[88][87] = 9'b111111111;
assign micromatrizz[88][88] = 9'b111111111;
assign micromatrizz[88][89] = 9'b111111111;
assign micromatrizz[88][90] = 9'b111111111;
assign micromatrizz[88][91] = 9'b111111111;
assign micromatrizz[88][92] = 9'b111111111;
assign micromatrizz[88][93] = 9'b111111111;
assign micromatrizz[88][94] = 9'b111111111;
assign micromatrizz[88][95] = 9'b111111111;
assign micromatrizz[88][96] = 9'b111111111;
assign micromatrizz[88][97] = 9'b111111111;
assign micromatrizz[88][98] = 9'b111111111;
assign micromatrizz[88][99] = 9'b111111111;
assign micromatrizz[88][100] = 9'b111111111;
assign micromatrizz[88][101] = 9'b111111111;
assign micromatrizz[88][102] = 9'b111111111;
assign micromatrizz[88][103] = 9'b111111111;
assign micromatrizz[88][104] = 9'b111111111;
assign micromatrizz[88][105] = 9'b111111111;
assign micromatrizz[88][106] = 9'b111111111;
assign micromatrizz[88][107] = 9'b111111111;
assign micromatrizz[88][108] = 9'b111111111;
assign micromatrizz[88][109] = 9'b111111111;
assign micromatrizz[88][110] = 9'b111111111;
assign micromatrizz[88][111] = 9'b111111111;
assign micromatrizz[88][112] = 9'b111111111;
assign micromatrizz[88][113] = 9'b111111111;
assign micromatrizz[88][114] = 9'b111111111;
assign micromatrizz[88][115] = 9'b111111111;
assign micromatrizz[88][116] = 9'b111111111;
assign micromatrizz[88][117] = 9'b111111111;
assign micromatrizz[88][118] = 9'b111111111;
assign micromatrizz[88][119] = 9'b111111111;
assign micromatrizz[88][120] = 9'b111111111;
assign micromatrizz[88][121] = 9'b111111111;
assign micromatrizz[88][122] = 9'b111111111;
assign micromatrizz[88][123] = 9'b111111111;
assign micromatrizz[88][124] = 9'b111111111;
assign micromatrizz[88][125] = 9'b111111111;
assign micromatrizz[88][126] = 9'b111111111;
assign micromatrizz[88][127] = 9'b111111111;
assign micromatrizz[88][128] = 9'b111111111;
assign micromatrizz[88][129] = 9'b111111111;
assign micromatrizz[88][130] = 9'b111111111;
assign micromatrizz[88][131] = 9'b111111111;
assign micromatrizz[88][132] = 9'b111111111;
assign micromatrizz[88][133] = 9'b111111111;
assign micromatrizz[88][134] = 9'b111111111;
assign micromatrizz[88][135] = 9'b111111111;
assign micromatrizz[88][136] = 9'b111111111;
assign micromatrizz[88][137] = 9'b111111111;
assign micromatrizz[88][138] = 9'b111111111;
assign micromatrizz[88][139] = 9'b111111111;
assign micromatrizz[88][140] = 9'b111111111;
assign micromatrizz[88][141] = 9'b111111111;
assign micromatrizz[88][142] = 9'b111111111;
assign micromatrizz[88][143] = 9'b111111111;
assign micromatrizz[88][144] = 9'b111111111;
assign micromatrizz[88][145] = 9'b111111111;
assign micromatrizz[88][146] = 9'b111111111;
assign micromatrizz[88][147] = 9'b111111111;
assign micromatrizz[88][148] = 9'b111111111;
assign micromatrizz[88][149] = 9'b111111111;
assign micromatrizz[88][150] = 9'b111111111;
assign micromatrizz[88][151] = 9'b111111111;
assign micromatrizz[88][152] = 9'b111111111;
assign micromatrizz[88][153] = 9'b111111111;
assign micromatrizz[88][154] = 9'b111111111;
assign micromatrizz[88][155] = 9'b111111111;
assign micromatrizz[88][156] = 9'b111111111;
assign micromatrizz[88][157] = 9'b111111111;
assign micromatrizz[88][158] = 9'b111111111;
assign micromatrizz[88][159] = 9'b111111111;
assign micromatrizz[88][160] = 9'b111111111;
assign micromatrizz[88][161] = 9'b111111111;
assign micromatrizz[88][162] = 9'b111111111;
assign micromatrizz[88][163] = 9'b111111111;
assign micromatrizz[88][164] = 9'b111111111;
assign micromatrizz[88][165] = 9'b111111111;
assign micromatrizz[88][166] = 9'b111111111;
assign micromatrizz[88][167] = 9'b111111111;
assign micromatrizz[88][168] = 9'b111111111;
assign micromatrizz[88][169] = 9'b111111111;
assign micromatrizz[88][170] = 9'b111111111;
assign micromatrizz[88][171] = 9'b111111111;
assign micromatrizz[88][172] = 9'b111111111;
assign micromatrizz[88][173] = 9'b111111111;
assign micromatrizz[88][174] = 9'b111111111;
assign micromatrizz[88][175] = 9'b111111111;
assign micromatrizz[88][176] = 9'b111111111;
assign micromatrizz[88][177] = 9'b111111111;
assign micromatrizz[88][178] = 9'b111111111;
assign micromatrizz[88][179] = 9'b111111111;
assign micromatrizz[88][180] = 9'b111111111;
assign micromatrizz[88][181] = 9'b111111111;
assign micromatrizz[88][182] = 9'b111111111;
assign micromatrizz[88][183] = 9'b111111111;
assign micromatrizz[88][184] = 9'b111111111;
assign micromatrizz[88][185] = 9'b111111111;
assign micromatrizz[88][186] = 9'b111111111;
assign micromatrizz[88][187] = 9'b111111111;
assign micromatrizz[88][188] = 9'b111111111;
assign micromatrizz[88][189] = 9'b111111111;
assign micromatrizz[88][190] = 9'b111111111;
assign micromatrizz[88][191] = 9'b111111111;
assign micromatrizz[88][192] = 9'b111111111;
assign micromatrizz[88][193] = 9'b111111111;
assign micromatrizz[88][194] = 9'b111111111;
assign micromatrizz[88][195] = 9'b111111111;
assign micromatrizz[88][196] = 9'b111111111;
assign micromatrizz[88][197] = 9'b111111111;
assign micromatrizz[88][198] = 9'b111111111;
assign micromatrizz[88][199] = 9'b111111111;
assign micromatrizz[88][200] = 9'b111111111;
assign micromatrizz[88][201] = 9'b111111111;
assign micromatrizz[88][202] = 9'b111111111;
assign micromatrizz[88][203] = 9'b111111111;
assign micromatrizz[88][204] = 9'b111111111;
assign micromatrizz[88][205] = 9'b111111111;
assign micromatrizz[88][206] = 9'b111111111;
assign micromatrizz[88][207] = 9'b111111111;
assign micromatrizz[88][208] = 9'b111111111;
assign micromatrizz[88][209] = 9'b111111111;
assign micromatrizz[88][210] = 9'b111111111;
assign micromatrizz[88][211] = 9'b111111111;
assign micromatrizz[88][212] = 9'b111111111;
assign micromatrizz[88][213] = 9'b111111111;
assign micromatrizz[88][214] = 9'b111111111;
assign micromatrizz[88][215] = 9'b111111111;
assign micromatrizz[88][216] = 9'b111111111;
assign micromatrizz[88][217] = 9'b111111111;
assign micromatrizz[88][218] = 9'b111111111;
assign micromatrizz[88][219] = 9'b111111111;
assign micromatrizz[88][220] = 9'b111111111;
assign micromatrizz[88][221] = 9'b111111111;
assign micromatrizz[88][222] = 9'b111111111;
assign micromatrizz[88][223] = 9'b111111111;
assign micromatrizz[88][224] = 9'b111111111;
assign micromatrizz[88][225] = 9'b111111111;
assign micromatrizz[88][226] = 9'b111111111;
assign micromatrizz[88][227] = 9'b111111111;
assign micromatrizz[88][228] = 9'b111111111;
assign micromatrizz[88][229] = 9'b111111111;
assign micromatrizz[88][230] = 9'b111111111;
assign micromatrizz[88][231] = 9'b111111111;
assign micromatrizz[88][232] = 9'b111111111;
assign micromatrizz[88][233] = 9'b111111111;
assign micromatrizz[88][234] = 9'b111111111;
assign micromatrizz[88][235] = 9'b111111111;
assign micromatrizz[88][236] = 9'b111111111;
assign micromatrizz[88][237] = 9'b111111111;
assign micromatrizz[88][238] = 9'b111111111;
assign micromatrizz[88][239] = 9'b111111111;
assign micromatrizz[88][240] = 9'b111111111;
assign micromatrizz[88][241] = 9'b111111111;
assign micromatrizz[88][242] = 9'b111111111;
assign micromatrizz[88][243] = 9'b111111111;
assign micromatrizz[88][244] = 9'b111111111;
assign micromatrizz[88][245] = 9'b111111111;
assign micromatrizz[88][246] = 9'b111111111;
assign micromatrizz[88][247] = 9'b111111111;
assign micromatrizz[88][248] = 9'b111111111;
assign micromatrizz[88][249] = 9'b111111111;
assign micromatrizz[88][250] = 9'b111111111;
assign micromatrizz[88][251] = 9'b111111111;
assign micromatrizz[88][252] = 9'b111111111;
assign micromatrizz[88][253] = 9'b111111111;
assign micromatrizz[88][254] = 9'b111111111;
assign micromatrizz[88][255] = 9'b111111111;
assign micromatrizz[88][256] = 9'b111111111;
assign micromatrizz[88][257] = 9'b111111111;
assign micromatrizz[88][258] = 9'b111111111;
assign micromatrizz[88][259] = 9'b111111111;
assign micromatrizz[88][260] = 9'b111111111;
assign micromatrizz[88][261] = 9'b111111111;
assign micromatrizz[88][262] = 9'b111111111;
assign micromatrizz[88][263] = 9'b111111111;
assign micromatrizz[88][264] = 9'b111111111;
assign micromatrizz[88][265] = 9'b111111111;
assign micromatrizz[88][266] = 9'b111111111;
assign micromatrizz[88][267] = 9'b111111111;
assign micromatrizz[88][268] = 9'b111111111;
assign micromatrizz[88][269] = 9'b111111111;
assign micromatrizz[88][270] = 9'b111111111;
assign micromatrizz[88][271] = 9'b111111111;
assign micromatrizz[88][272] = 9'b111111111;
assign micromatrizz[88][273] = 9'b111111111;
assign micromatrizz[88][274] = 9'b111111111;
assign micromatrizz[88][275] = 9'b111111111;
assign micromatrizz[88][276] = 9'b111111111;
assign micromatrizz[88][277] = 9'b111111111;
assign micromatrizz[88][278] = 9'b111111111;
assign micromatrizz[88][279] = 9'b111111111;
assign micromatrizz[88][280] = 9'b111111111;
assign micromatrizz[88][281] = 9'b111111111;
assign micromatrizz[88][282] = 9'b111111111;
assign micromatrizz[88][283] = 9'b111111111;
assign micromatrizz[88][284] = 9'b111111111;
assign micromatrizz[88][285] = 9'b111111111;
assign micromatrizz[88][286] = 9'b111111111;
assign micromatrizz[88][287] = 9'b111111111;
assign micromatrizz[88][288] = 9'b111111111;
assign micromatrizz[88][289] = 9'b111111111;
assign micromatrizz[88][290] = 9'b111111111;
assign micromatrizz[88][291] = 9'b111111111;
assign micromatrizz[88][292] = 9'b111111111;
assign micromatrizz[88][293] = 9'b111111111;
assign micromatrizz[88][294] = 9'b111111111;
assign micromatrizz[88][295] = 9'b111111111;
assign micromatrizz[88][296] = 9'b111111111;
assign micromatrizz[88][297] = 9'b111111111;
assign micromatrizz[88][298] = 9'b111111111;
assign micromatrizz[88][299] = 9'b111111111;
assign micromatrizz[88][300] = 9'b111111111;
assign micromatrizz[88][301] = 9'b111111111;
assign micromatrizz[88][302] = 9'b111111111;
assign micromatrizz[88][303] = 9'b111111111;
assign micromatrizz[88][304] = 9'b111111111;
assign micromatrizz[88][305] = 9'b111111111;
assign micromatrizz[88][306] = 9'b111111111;
assign micromatrizz[88][307] = 9'b111111111;
assign micromatrizz[88][308] = 9'b111111111;
assign micromatrizz[88][309] = 9'b111111111;
assign micromatrizz[88][310] = 9'b111111111;
assign micromatrizz[88][311] = 9'b111111111;
assign micromatrizz[88][312] = 9'b111111111;
assign micromatrizz[88][313] = 9'b111111111;
assign micromatrizz[88][314] = 9'b111111111;
assign micromatrizz[88][315] = 9'b111111111;
assign micromatrizz[88][316] = 9'b111111111;
assign micromatrizz[88][317] = 9'b111111111;
assign micromatrizz[88][318] = 9'b111111111;
assign micromatrizz[88][319] = 9'b111111111;
assign micromatrizz[88][320] = 9'b111111111;
assign micromatrizz[88][321] = 9'b111111111;
assign micromatrizz[88][322] = 9'b111111111;
assign micromatrizz[88][323] = 9'b111111111;
assign micromatrizz[88][324] = 9'b111111111;
assign micromatrizz[88][325] = 9'b111111111;
assign micromatrizz[88][326] = 9'b111111111;
assign micromatrizz[88][327] = 9'b111111111;
assign micromatrizz[88][328] = 9'b111111111;
assign micromatrizz[88][329] = 9'b111111111;
assign micromatrizz[88][330] = 9'b111111111;
assign micromatrizz[88][331] = 9'b111111111;
assign micromatrizz[88][332] = 9'b111111111;
assign micromatrizz[88][333] = 9'b111111111;
assign micromatrizz[88][334] = 9'b111111111;
assign micromatrizz[88][335] = 9'b111111111;
assign micromatrizz[88][336] = 9'b111111111;
assign micromatrizz[88][337] = 9'b111111111;
assign micromatrizz[88][338] = 9'b111111111;
assign micromatrizz[88][339] = 9'b111111111;
assign micromatrizz[88][340] = 9'b111111111;
assign micromatrizz[88][341] = 9'b111111111;
assign micromatrizz[88][342] = 9'b111111111;
assign micromatrizz[88][343] = 9'b111111111;
assign micromatrizz[88][344] = 9'b111111111;
assign micromatrizz[88][345] = 9'b111111111;
assign micromatrizz[88][346] = 9'b111111111;
assign micromatrizz[88][347] = 9'b111111111;
assign micromatrizz[88][348] = 9'b111111111;
assign micromatrizz[88][349] = 9'b111111111;
assign micromatrizz[88][350] = 9'b111111111;
assign micromatrizz[88][351] = 9'b111111111;
assign micromatrizz[88][352] = 9'b111111111;
assign micromatrizz[88][353] = 9'b111111111;
assign micromatrizz[88][354] = 9'b111111111;
assign micromatrizz[88][355] = 9'b111111111;
assign micromatrizz[88][356] = 9'b111111111;
assign micromatrizz[88][357] = 9'b111111111;
assign micromatrizz[88][358] = 9'b111111111;
assign micromatrizz[88][359] = 9'b111111111;
assign micromatrizz[88][360] = 9'b111111111;
assign micromatrizz[88][361] = 9'b111111111;
assign micromatrizz[88][362] = 9'b111111111;
assign micromatrizz[88][363] = 9'b111111111;
assign micromatrizz[88][364] = 9'b111111111;
assign micromatrizz[88][365] = 9'b111111111;
assign micromatrizz[88][366] = 9'b111111111;
assign micromatrizz[88][367] = 9'b111111111;
assign micromatrizz[88][368] = 9'b111111111;
assign micromatrizz[88][369] = 9'b111111111;
assign micromatrizz[88][370] = 9'b111111111;
assign micromatrizz[88][371] = 9'b111111111;
assign micromatrizz[88][372] = 9'b111111111;
assign micromatrizz[88][373] = 9'b111111111;
assign micromatrizz[88][374] = 9'b111111111;
assign micromatrizz[88][375] = 9'b111111111;
assign micromatrizz[88][376] = 9'b111111111;
assign micromatrizz[88][377] = 9'b111111111;
assign micromatrizz[88][378] = 9'b111111111;
assign micromatrizz[88][379] = 9'b111111111;
assign micromatrizz[88][380] = 9'b111111111;
assign micromatrizz[88][381] = 9'b111111111;
assign micromatrizz[88][382] = 9'b111111111;
assign micromatrizz[88][383] = 9'b111111111;
assign micromatrizz[88][384] = 9'b111111111;
assign micromatrizz[88][385] = 9'b111111111;
assign micromatrizz[88][386] = 9'b111111111;
assign micromatrizz[88][387] = 9'b111111111;
assign micromatrizz[88][388] = 9'b111111111;
assign micromatrizz[88][389] = 9'b111111111;
assign micromatrizz[88][390] = 9'b111111111;
assign micromatrizz[88][391] = 9'b111111111;
assign micromatrizz[88][392] = 9'b111111111;
assign micromatrizz[88][393] = 9'b111111111;
assign micromatrizz[88][394] = 9'b111111111;
assign micromatrizz[88][395] = 9'b111111111;
assign micromatrizz[88][396] = 9'b111111111;
assign micromatrizz[88][397] = 9'b111111111;
assign micromatrizz[88][398] = 9'b111111111;
assign micromatrizz[88][399] = 9'b111111111;
assign micromatrizz[88][400] = 9'b111111111;
assign micromatrizz[88][401] = 9'b111111111;
assign micromatrizz[88][402] = 9'b111111111;
assign micromatrizz[88][403] = 9'b111111111;
assign micromatrizz[88][404] = 9'b111111111;
assign micromatrizz[88][405] = 9'b111111111;
assign micromatrizz[88][406] = 9'b111111111;
assign micromatrizz[88][407] = 9'b111111111;
assign micromatrizz[88][408] = 9'b111111111;
assign micromatrizz[88][409] = 9'b111111111;
assign micromatrizz[88][410] = 9'b111111111;
assign micromatrizz[88][411] = 9'b111111111;
assign micromatrizz[88][412] = 9'b111111111;
assign micromatrizz[88][413] = 9'b111111111;
assign micromatrizz[88][414] = 9'b111111111;
assign micromatrizz[88][415] = 9'b111111111;
assign micromatrizz[88][416] = 9'b111111111;
assign micromatrizz[88][417] = 9'b111111111;
assign micromatrizz[88][418] = 9'b111111111;
assign micromatrizz[88][419] = 9'b111111111;
assign micromatrizz[88][420] = 9'b111111111;
assign micromatrizz[88][421] = 9'b111111111;
assign micromatrizz[88][422] = 9'b111111111;
assign micromatrizz[88][423] = 9'b111111111;
assign micromatrizz[88][424] = 9'b111111111;
assign micromatrizz[88][425] = 9'b111111111;
assign micromatrizz[88][426] = 9'b111111111;
assign micromatrizz[88][427] = 9'b111111111;
assign micromatrizz[88][428] = 9'b111111111;
assign micromatrizz[88][429] = 9'b111111111;
assign micromatrizz[88][430] = 9'b111111111;
assign micromatrizz[88][431] = 9'b111111111;
assign micromatrizz[88][432] = 9'b111111111;
assign micromatrizz[88][433] = 9'b111111111;
assign micromatrizz[88][434] = 9'b111111111;
assign micromatrizz[88][435] = 9'b111111111;
assign micromatrizz[88][436] = 9'b111111111;
assign micromatrizz[88][437] = 9'b111111111;
assign micromatrizz[88][438] = 9'b111111111;
assign micromatrizz[88][439] = 9'b111111111;
assign micromatrizz[88][440] = 9'b111111111;
assign micromatrizz[88][441] = 9'b111111111;
assign micromatrizz[88][442] = 9'b111111111;
assign micromatrizz[88][443] = 9'b111111111;
assign micromatrizz[88][444] = 9'b111111111;
assign micromatrizz[88][445] = 9'b111111111;
assign micromatrizz[88][446] = 9'b111111111;
assign micromatrizz[88][447] = 9'b111111111;
assign micromatrizz[88][448] = 9'b111111111;
assign micromatrizz[88][449] = 9'b111111111;
assign micromatrizz[88][450] = 9'b111111111;
assign micromatrizz[88][451] = 9'b111111111;
assign micromatrizz[88][452] = 9'b111111111;
assign micromatrizz[88][453] = 9'b111111111;
assign micromatrizz[88][454] = 9'b111111111;
assign micromatrizz[88][455] = 9'b111111111;
assign micromatrizz[88][456] = 9'b111111111;
assign micromatrizz[88][457] = 9'b111111111;
assign micromatrizz[88][458] = 9'b111111111;
assign micromatrizz[88][459] = 9'b111111111;
assign micromatrizz[88][460] = 9'b111111111;
assign micromatrizz[88][461] = 9'b111111111;
assign micromatrizz[88][462] = 9'b111111111;
assign micromatrizz[88][463] = 9'b111111111;
assign micromatrizz[88][464] = 9'b111111111;
assign micromatrizz[88][465] = 9'b111111111;
assign micromatrizz[88][466] = 9'b111111111;
assign micromatrizz[88][467] = 9'b111111111;
assign micromatrizz[88][468] = 9'b111111111;
assign micromatrizz[88][469] = 9'b111111111;
assign micromatrizz[88][470] = 9'b111111111;
assign micromatrizz[88][471] = 9'b111111111;
assign micromatrizz[88][472] = 9'b111111111;
assign micromatrizz[88][473] = 9'b111111111;
assign micromatrizz[88][474] = 9'b111111111;
assign micromatrizz[88][475] = 9'b111111111;
assign micromatrizz[88][476] = 9'b111111111;
assign micromatrizz[88][477] = 9'b111111111;
assign micromatrizz[88][478] = 9'b111111111;
assign micromatrizz[88][479] = 9'b111111111;
assign micromatrizz[88][480] = 9'b111111111;
assign micromatrizz[88][481] = 9'b111111111;
assign micromatrizz[88][482] = 9'b111111111;
assign micromatrizz[88][483] = 9'b111111111;
assign micromatrizz[88][484] = 9'b111111111;
assign micromatrizz[88][485] = 9'b111111111;
assign micromatrizz[88][486] = 9'b111111111;
assign micromatrizz[88][487] = 9'b111111111;
assign micromatrizz[88][488] = 9'b111111111;
assign micromatrizz[88][489] = 9'b111111111;
assign micromatrizz[88][490] = 9'b111111111;
assign micromatrizz[88][491] = 9'b111111111;
assign micromatrizz[88][492] = 9'b111111111;
assign micromatrizz[88][493] = 9'b111111111;
assign micromatrizz[88][494] = 9'b111111111;
assign micromatrizz[88][495] = 9'b111111111;
assign micromatrizz[88][496] = 9'b111111111;
assign micromatrizz[88][497] = 9'b111111111;
assign micromatrizz[88][498] = 9'b111111111;
assign micromatrizz[88][499] = 9'b111111111;
assign micromatrizz[88][500] = 9'b111111111;
assign micromatrizz[88][501] = 9'b111111111;
assign micromatrizz[88][502] = 9'b111111111;
assign micromatrizz[88][503] = 9'b111111111;
assign micromatrizz[88][504] = 9'b111111111;
assign micromatrizz[88][505] = 9'b111111111;
assign micromatrizz[88][506] = 9'b111111111;
assign micromatrizz[88][507] = 9'b111111111;
assign micromatrizz[88][508] = 9'b111111111;
assign micromatrizz[88][509] = 9'b111111111;
assign micromatrizz[88][510] = 9'b111111111;
assign micromatrizz[88][511] = 9'b111111111;
assign micromatrizz[88][512] = 9'b111111111;
assign micromatrizz[88][513] = 9'b111111111;
assign micromatrizz[88][514] = 9'b111111111;
assign micromatrizz[88][515] = 9'b111111111;
assign micromatrizz[88][516] = 9'b111111111;
assign micromatrizz[88][517] = 9'b111111111;
assign micromatrizz[88][518] = 9'b111111111;
assign micromatrizz[88][519] = 9'b111111111;
assign micromatrizz[88][520] = 9'b111111111;
assign micromatrizz[88][521] = 9'b111111111;
assign micromatrizz[88][522] = 9'b111111111;
assign micromatrizz[88][523] = 9'b111111111;
assign micromatrizz[88][524] = 9'b111111111;
assign micromatrizz[88][525] = 9'b111111111;
assign micromatrizz[88][526] = 9'b111111111;
assign micromatrizz[88][527] = 9'b111111111;
assign micromatrizz[88][528] = 9'b111111111;
assign micromatrizz[88][529] = 9'b111111111;
assign micromatrizz[88][530] = 9'b111111111;
assign micromatrizz[88][531] = 9'b111111111;
assign micromatrizz[88][532] = 9'b111111111;
assign micromatrizz[88][533] = 9'b111111111;
assign micromatrizz[88][534] = 9'b111111111;
assign micromatrizz[88][535] = 9'b111111111;
assign micromatrizz[88][536] = 9'b111111111;
assign micromatrizz[88][537] = 9'b111111111;
assign micromatrizz[88][538] = 9'b111111111;
assign micromatrizz[88][539] = 9'b111111111;
assign micromatrizz[88][540] = 9'b111111111;
assign micromatrizz[88][541] = 9'b111111111;
assign micromatrizz[88][542] = 9'b111111111;
assign micromatrizz[88][543] = 9'b111111111;
assign micromatrizz[88][544] = 9'b111111111;
assign micromatrizz[88][545] = 9'b111111111;
assign micromatrizz[88][546] = 9'b111111111;
assign micromatrizz[88][547] = 9'b111111111;
assign micromatrizz[88][548] = 9'b111111111;
assign micromatrizz[88][549] = 9'b111111111;
assign micromatrizz[88][550] = 9'b111111111;
assign micromatrizz[88][551] = 9'b111111111;
assign micromatrizz[88][552] = 9'b111111111;
assign micromatrizz[88][553] = 9'b111111111;
assign micromatrizz[88][554] = 9'b111111111;
assign micromatrizz[88][555] = 9'b111111111;
assign micromatrizz[88][556] = 9'b111111111;
assign micromatrizz[88][557] = 9'b111111111;
assign micromatrizz[88][558] = 9'b111111111;
assign micromatrizz[88][559] = 9'b111111111;
assign micromatrizz[88][560] = 9'b111111111;
assign micromatrizz[88][561] = 9'b111111111;
assign micromatrizz[88][562] = 9'b111111111;
assign micromatrizz[88][563] = 9'b111111111;
assign micromatrizz[88][564] = 9'b111111111;
assign micromatrizz[88][565] = 9'b111111111;
assign micromatrizz[88][566] = 9'b111111111;
assign micromatrizz[88][567] = 9'b111111111;
assign micromatrizz[88][568] = 9'b111111111;
assign micromatrizz[88][569] = 9'b111111111;
assign micromatrizz[88][570] = 9'b111111111;
assign micromatrizz[88][571] = 9'b111111111;
assign micromatrizz[88][572] = 9'b111111111;
assign micromatrizz[88][573] = 9'b111111111;
assign micromatrizz[88][574] = 9'b111111111;
assign micromatrizz[88][575] = 9'b111111111;
assign micromatrizz[88][576] = 9'b111111111;
assign micromatrizz[88][577] = 9'b111111111;
assign micromatrizz[88][578] = 9'b111111111;
assign micromatrizz[88][579] = 9'b111111111;
assign micromatrizz[88][580] = 9'b111111111;
assign micromatrizz[88][581] = 9'b111111111;
assign micromatrizz[88][582] = 9'b111111111;
assign micromatrizz[88][583] = 9'b111111111;
assign micromatrizz[88][584] = 9'b111111111;
assign micromatrizz[88][585] = 9'b111111111;
assign micromatrizz[88][586] = 9'b111111111;
assign micromatrizz[88][587] = 9'b111111111;
assign micromatrizz[88][588] = 9'b111111111;
assign micromatrizz[88][589] = 9'b111111111;
assign micromatrizz[88][590] = 9'b111111111;
assign micromatrizz[88][591] = 9'b111111111;
assign micromatrizz[88][592] = 9'b111111111;
assign micromatrizz[88][593] = 9'b111111111;
assign micromatrizz[88][594] = 9'b111111111;
assign micromatrizz[88][595] = 9'b111111111;
assign micromatrizz[88][596] = 9'b111111111;
assign micromatrizz[88][597] = 9'b111111111;
assign micromatrizz[88][598] = 9'b111111111;
assign micromatrizz[88][599] = 9'b111111111;
assign micromatrizz[88][600] = 9'b111111111;
assign micromatrizz[88][601] = 9'b111111111;
assign micromatrizz[88][602] = 9'b111111111;
assign micromatrizz[88][603] = 9'b111111111;
assign micromatrizz[88][604] = 9'b111111111;
assign micromatrizz[88][605] = 9'b111111111;
assign micromatrizz[88][606] = 9'b111111111;
assign micromatrizz[88][607] = 9'b111111111;
assign micromatrizz[88][608] = 9'b111111111;
assign micromatrizz[88][609] = 9'b111111111;
assign micromatrizz[88][610] = 9'b111111111;
assign micromatrizz[88][611] = 9'b111111111;
assign micromatrizz[88][612] = 9'b111111111;
assign micromatrizz[88][613] = 9'b111111111;
assign micromatrizz[88][614] = 9'b111111111;
assign micromatrizz[88][615] = 9'b111111111;
assign micromatrizz[88][616] = 9'b111111111;
assign micromatrizz[88][617] = 9'b111111111;
assign micromatrizz[88][618] = 9'b111111111;
assign micromatrizz[88][619] = 9'b111111111;
assign micromatrizz[88][620] = 9'b111111111;
assign micromatrizz[88][621] = 9'b111111111;
assign micromatrizz[88][622] = 9'b111111111;
assign micromatrizz[88][623] = 9'b111111111;
assign micromatrizz[88][624] = 9'b111111111;
assign micromatrizz[88][625] = 9'b111111111;
assign micromatrizz[88][626] = 9'b111111111;
assign micromatrizz[88][627] = 9'b111111111;
assign micromatrizz[88][628] = 9'b111111111;
assign micromatrizz[88][629] = 9'b111111111;
assign micromatrizz[88][630] = 9'b111111111;
assign micromatrizz[88][631] = 9'b111111111;
assign micromatrizz[88][632] = 9'b111111111;
assign micromatrizz[88][633] = 9'b111111111;
assign micromatrizz[88][634] = 9'b111111111;
assign micromatrizz[88][635] = 9'b111111111;
assign micromatrizz[88][636] = 9'b111111111;
assign micromatrizz[88][637] = 9'b111111111;
assign micromatrizz[88][638] = 9'b111111111;
assign micromatrizz[88][639] = 9'b111111111;
assign micromatrizz[89][0] = 9'b111111111;
assign micromatrizz[89][1] = 9'b111111111;
assign micromatrizz[89][2] = 9'b111111111;
assign micromatrizz[89][3] = 9'b111111111;
assign micromatrizz[89][4] = 9'b111111111;
assign micromatrizz[89][5] = 9'b111111111;
assign micromatrizz[89][6] = 9'b111111111;
assign micromatrizz[89][7] = 9'b111111111;
assign micromatrizz[89][8] = 9'b111111111;
assign micromatrizz[89][9] = 9'b111111111;
assign micromatrizz[89][10] = 9'b111111111;
assign micromatrizz[89][11] = 9'b111111111;
assign micromatrizz[89][12] = 9'b111111111;
assign micromatrizz[89][13] = 9'b111111111;
assign micromatrizz[89][14] = 9'b111111111;
assign micromatrizz[89][15] = 9'b111111111;
assign micromatrizz[89][16] = 9'b111111111;
assign micromatrizz[89][17] = 9'b111111111;
assign micromatrizz[89][18] = 9'b111111111;
assign micromatrizz[89][19] = 9'b111111111;
assign micromatrizz[89][20] = 9'b111111111;
assign micromatrizz[89][21] = 9'b111111111;
assign micromatrizz[89][22] = 9'b111111111;
assign micromatrizz[89][23] = 9'b111111111;
assign micromatrizz[89][24] = 9'b111111111;
assign micromatrizz[89][25] = 9'b111111111;
assign micromatrizz[89][26] = 9'b111111111;
assign micromatrizz[89][27] = 9'b111111111;
assign micromatrizz[89][28] = 9'b111111111;
assign micromatrizz[89][29] = 9'b111111111;
assign micromatrizz[89][30] = 9'b111111111;
assign micromatrizz[89][31] = 9'b111111111;
assign micromatrizz[89][32] = 9'b111111111;
assign micromatrizz[89][33] = 9'b111111111;
assign micromatrizz[89][34] = 9'b111111111;
assign micromatrizz[89][35] = 9'b111111111;
assign micromatrizz[89][36] = 9'b111111111;
assign micromatrizz[89][37] = 9'b111111111;
assign micromatrizz[89][38] = 9'b111111111;
assign micromatrizz[89][39] = 9'b111111111;
assign micromatrizz[89][40] = 9'b111111111;
assign micromatrizz[89][41] = 9'b111111111;
assign micromatrizz[89][42] = 9'b111111111;
assign micromatrizz[89][43] = 9'b111111111;
assign micromatrizz[89][44] = 9'b111111111;
assign micromatrizz[89][45] = 9'b111111111;
assign micromatrizz[89][46] = 9'b111111111;
assign micromatrizz[89][47] = 9'b111111111;
assign micromatrizz[89][48] = 9'b111111111;
assign micromatrizz[89][49] = 9'b111111111;
assign micromatrizz[89][50] = 9'b111111111;
assign micromatrizz[89][51] = 9'b111111111;
assign micromatrizz[89][52] = 9'b111111111;
assign micromatrizz[89][53] = 9'b111111111;
assign micromatrizz[89][54] = 9'b111111111;
assign micromatrizz[89][55] = 9'b111111111;
assign micromatrizz[89][56] = 9'b111111111;
assign micromatrizz[89][57] = 9'b111111111;
assign micromatrizz[89][58] = 9'b111111111;
assign micromatrizz[89][59] = 9'b111111111;
assign micromatrizz[89][60] = 9'b111111111;
assign micromatrizz[89][61] = 9'b111111111;
assign micromatrizz[89][62] = 9'b111111111;
assign micromatrizz[89][63] = 9'b111111111;
assign micromatrizz[89][64] = 9'b111111111;
assign micromatrizz[89][65] = 9'b111111111;
assign micromatrizz[89][66] = 9'b111111111;
assign micromatrizz[89][67] = 9'b111111111;
assign micromatrizz[89][68] = 9'b111111111;
assign micromatrizz[89][69] = 9'b111111111;
assign micromatrizz[89][70] = 9'b111111111;
assign micromatrizz[89][71] = 9'b111111111;
assign micromatrizz[89][72] = 9'b111111111;
assign micromatrizz[89][73] = 9'b111111111;
assign micromatrizz[89][74] = 9'b111111111;
assign micromatrizz[89][75] = 9'b111111111;
assign micromatrizz[89][76] = 9'b111111111;
assign micromatrizz[89][77] = 9'b111111111;
assign micromatrizz[89][78] = 9'b111111111;
assign micromatrizz[89][79] = 9'b111111111;
assign micromatrizz[89][80] = 9'b111111111;
assign micromatrizz[89][81] = 9'b111111111;
assign micromatrizz[89][82] = 9'b111111111;
assign micromatrizz[89][83] = 9'b111111111;
assign micromatrizz[89][84] = 9'b111111111;
assign micromatrizz[89][85] = 9'b111111111;
assign micromatrizz[89][86] = 9'b111111111;
assign micromatrizz[89][87] = 9'b111111111;
assign micromatrizz[89][88] = 9'b111111111;
assign micromatrizz[89][89] = 9'b111111111;
assign micromatrizz[89][90] = 9'b111111111;
assign micromatrizz[89][91] = 9'b111111111;
assign micromatrizz[89][92] = 9'b111111111;
assign micromatrizz[89][93] = 9'b111111111;
assign micromatrizz[89][94] = 9'b111111111;
assign micromatrizz[89][95] = 9'b111111111;
assign micromatrizz[89][96] = 9'b111111111;
assign micromatrizz[89][97] = 9'b111111111;
assign micromatrizz[89][98] = 9'b111111111;
assign micromatrizz[89][99] = 9'b111111111;
assign micromatrizz[89][100] = 9'b111111111;
assign micromatrizz[89][101] = 9'b111111111;
assign micromatrizz[89][102] = 9'b111111111;
assign micromatrizz[89][103] = 9'b111111111;
assign micromatrizz[89][104] = 9'b111111111;
assign micromatrizz[89][105] = 9'b111111111;
assign micromatrizz[89][106] = 9'b111111111;
assign micromatrizz[89][107] = 9'b111111111;
assign micromatrizz[89][108] = 9'b111111111;
assign micromatrizz[89][109] = 9'b111111111;
assign micromatrizz[89][110] = 9'b111111111;
assign micromatrizz[89][111] = 9'b111111111;
assign micromatrizz[89][112] = 9'b111111111;
assign micromatrizz[89][113] = 9'b111111111;
assign micromatrizz[89][114] = 9'b111111111;
assign micromatrizz[89][115] = 9'b111111111;
assign micromatrizz[89][116] = 9'b111111111;
assign micromatrizz[89][117] = 9'b111111111;
assign micromatrizz[89][118] = 9'b111111111;
assign micromatrizz[89][119] = 9'b111111111;
assign micromatrizz[89][120] = 9'b111111111;
assign micromatrizz[89][121] = 9'b111111111;
assign micromatrizz[89][122] = 9'b111111111;
assign micromatrizz[89][123] = 9'b111111111;
assign micromatrizz[89][124] = 9'b111111111;
assign micromatrizz[89][125] = 9'b111111111;
assign micromatrizz[89][126] = 9'b111111111;
assign micromatrizz[89][127] = 9'b111111111;
assign micromatrizz[89][128] = 9'b111111111;
assign micromatrizz[89][129] = 9'b111111111;
assign micromatrizz[89][130] = 9'b111111111;
assign micromatrizz[89][131] = 9'b111111111;
assign micromatrizz[89][132] = 9'b111111111;
assign micromatrizz[89][133] = 9'b111111111;
assign micromatrizz[89][134] = 9'b111111111;
assign micromatrizz[89][135] = 9'b111111111;
assign micromatrizz[89][136] = 9'b111111111;
assign micromatrizz[89][137] = 9'b111111111;
assign micromatrizz[89][138] = 9'b111111111;
assign micromatrizz[89][139] = 9'b111111111;
assign micromatrizz[89][140] = 9'b111111111;
assign micromatrizz[89][141] = 9'b111111111;
assign micromatrizz[89][142] = 9'b111111111;
assign micromatrizz[89][143] = 9'b111111111;
assign micromatrizz[89][144] = 9'b111111111;
assign micromatrizz[89][145] = 9'b111111111;
assign micromatrizz[89][146] = 9'b111111111;
assign micromatrizz[89][147] = 9'b111111111;
assign micromatrizz[89][148] = 9'b111111111;
assign micromatrizz[89][149] = 9'b111111111;
assign micromatrizz[89][150] = 9'b111111111;
assign micromatrizz[89][151] = 9'b111111111;
assign micromatrizz[89][152] = 9'b111111111;
assign micromatrizz[89][153] = 9'b111111111;
assign micromatrizz[89][154] = 9'b111111111;
assign micromatrizz[89][155] = 9'b111111111;
assign micromatrizz[89][156] = 9'b111111111;
assign micromatrizz[89][157] = 9'b111111111;
assign micromatrizz[89][158] = 9'b111111111;
assign micromatrizz[89][159] = 9'b111111111;
assign micromatrizz[89][160] = 9'b111111111;
assign micromatrizz[89][161] = 9'b111111111;
assign micromatrizz[89][162] = 9'b111111111;
assign micromatrizz[89][163] = 9'b111111111;
assign micromatrizz[89][164] = 9'b111111111;
assign micromatrizz[89][165] = 9'b111111111;
assign micromatrizz[89][166] = 9'b111111111;
assign micromatrizz[89][167] = 9'b111111111;
assign micromatrizz[89][168] = 9'b111111111;
assign micromatrizz[89][169] = 9'b111111111;
assign micromatrizz[89][170] = 9'b111111111;
assign micromatrizz[89][171] = 9'b111111111;
assign micromatrizz[89][172] = 9'b111111111;
assign micromatrizz[89][173] = 9'b111111111;
assign micromatrizz[89][174] = 9'b111111111;
assign micromatrizz[89][175] = 9'b111111111;
assign micromatrizz[89][176] = 9'b111111111;
assign micromatrizz[89][177] = 9'b111111111;
assign micromatrizz[89][178] = 9'b111111111;
assign micromatrizz[89][179] = 9'b111111111;
assign micromatrizz[89][180] = 9'b111111111;
assign micromatrizz[89][181] = 9'b111111111;
assign micromatrizz[89][182] = 9'b111111111;
assign micromatrizz[89][183] = 9'b111111111;
assign micromatrizz[89][184] = 9'b111111111;
assign micromatrizz[89][185] = 9'b111111111;
assign micromatrizz[89][186] = 9'b111111111;
assign micromatrizz[89][187] = 9'b111111111;
assign micromatrizz[89][188] = 9'b111111111;
assign micromatrizz[89][189] = 9'b111111111;
assign micromatrizz[89][190] = 9'b111111111;
assign micromatrizz[89][191] = 9'b111111111;
assign micromatrizz[89][192] = 9'b111111111;
assign micromatrizz[89][193] = 9'b111111111;
assign micromatrizz[89][194] = 9'b111111111;
assign micromatrizz[89][195] = 9'b111111111;
assign micromatrizz[89][196] = 9'b111111111;
assign micromatrizz[89][197] = 9'b111111111;
assign micromatrizz[89][198] = 9'b111111111;
assign micromatrizz[89][199] = 9'b111111111;
assign micromatrizz[89][200] = 9'b111111111;
assign micromatrizz[89][201] = 9'b111111111;
assign micromatrizz[89][202] = 9'b111111111;
assign micromatrizz[89][203] = 9'b111111111;
assign micromatrizz[89][204] = 9'b111111111;
assign micromatrizz[89][205] = 9'b111111111;
assign micromatrizz[89][206] = 9'b111111111;
assign micromatrizz[89][207] = 9'b111111111;
assign micromatrizz[89][208] = 9'b111111111;
assign micromatrizz[89][209] = 9'b111111111;
assign micromatrizz[89][210] = 9'b111111111;
assign micromatrizz[89][211] = 9'b111111111;
assign micromatrizz[89][212] = 9'b111111111;
assign micromatrizz[89][213] = 9'b111111111;
assign micromatrizz[89][214] = 9'b111111111;
assign micromatrizz[89][215] = 9'b111111111;
assign micromatrizz[89][216] = 9'b111111111;
assign micromatrizz[89][217] = 9'b111111111;
assign micromatrizz[89][218] = 9'b111111111;
assign micromatrizz[89][219] = 9'b111111111;
assign micromatrizz[89][220] = 9'b111111111;
assign micromatrizz[89][221] = 9'b111111111;
assign micromatrizz[89][222] = 9'b111111111;
assign micromatrizz[89][223] = 9'b111111111;
assign micromatrizz[89][224] = 9'b111111111;
assign micromatrizz[89][225] = 9'b111111111;
assign micromatrizz[89][226] = 9'b111111111;
assign micromatrizz[89][227] = 9'b111111111;
assign micromatrizz[89][228] = 9'b111111111;
assign micromatrizz[89][229] = 9'b111111111;
assign micromatrizz[89][230] = 9'b111111111;
assign micromatrizz[89][231] = 9'b111111111;
assign micromatrizz[89][232] = 9'b111111111;
assign micromatrizz[89][233] = 9'b111111111;
assign micromatrizz[89][234] = 9'b111111111;
assign micromatrizz[89][235] = 9'b111111111;
assign micromatrizz[89][236] = 9'b111111111;
assign micromatrizz[89][237] = 9'b111111111;
assign micromatrizz[89][238] = 9'b111111111;
assign micromatrizz[89][239] = 9'b111111111;
assign micromatrizz[89][240] = 9'b111111111;
assign micromatrizz[89][241] = 9'b111111111;
assign micromatrizz[89][242] = 9'b111111111;
assign micromatrizz[89][243] = 9'b111111111;
assign micromatrizz[89][244] = 9'b111111111;
assign micromatrizz[89][245] = 9'b111111111;
assign micromatrizz[89][246] = 9'b111111111;
assign micromatrizz[89][247] = 9'b111111111;
assign micromatrizz[89][248] = 9'b111111111;
assign micromatrizz[89][249] = 9'b111111111;
assign micromatrizz[89][250] = 9'b111111111;
assign micromatrizz[89][251] = 9'b111111111;
assign micromatrizz[89][252] = 9'b111111111;
assign micromatrizz[89][253] = 9'b111111111;
assign micromatrizz[89][254] = 9'b111111111;
assign micromatrizz[89][255] = 9'b111111111;
assign micromatrizz[89][256] = 9'b111111111;
assign micromatrizz[89][257] = 9'b111111111;
assign micromatrizz[89][258] = 9'b111111111;
assign micromatrizz[89][259] = 9'b111111111;
assign micromatrizz[89][260] = 9'b111111111;
assign micromatrizz[89][261] = 9'b111111111;
assign micromatrizz[89][262] = 9'b111111111;
assign micromatrizz[89][263] = 9'b111111111;
assign micromatrizz[89][264] = 9'b111111111;
assign micromatrizz[89][265] = 9'b111111111;
assign micromatrizz[89][266] = 9'b111111111;
assign micromatrizz[89][267] = 9'b111111111;
assign micromatrizz[89][268] = 9'b111111111;
assign micromatrizz[89][269] = 9'b111111111;
assign micromatrizz[89][270] = 9'b111111111;
assign micromatrizz[89][271] = 9'b111111111;
assign micromatrizz[89][272] = 9'b111111111;
assign micromatrizz[89][273] = 9'b111111111;
assign micromatrizz[89][274] = 9'b111111111;
assign micromatrizz[89][275] = 9'b111111111;
assign micromatrizz[89][276] = 9'b111111111;
assign micromatrizz[89][277] = 9'b111111111;
assign micromatrizz[89][278] = 9'b111111111;
assign micromatrizz[89][279] = 9'b111111111;
assign micromatrizz[89][280] = 9'b111111111;
assign micromatrizz[89][281] = 9'b111111111;
assign micromatrizz[89][282] = 9'b111111111;
assign micromatrizz[89][283] = 9'b111111111;
assign micromatrizz[89][284] = 9'b111111111;
assign micromatrizz[89][285] = 9'b111111111;
assign micromatrizz[89][286] = 9'b111111111;
assign micromatrizz[89][287] = 9'b111111111;
assign micromatrizz[89][288] = 9'b111111111;
assign micromatrizz[89][289] = 9'b111111111;
assign micromatrizz[89][290] = 9'b111111111;
assign micromatrizz[89][291] = 9'b111111111;
assign micromatrizz[89][292] = 9'b111111111;
assign micromatrizz[89][293] = 9'b111111111;
assign micromatrizz[89][294] = 9'b111111111;
assign micromatrizz[89][295] = 9'b111111111;
assign micromatrizz[89][296] = 9'b111111111;
assign micromatrizz[89][297] = 9'b111111111;
assign micromatrizz[89][298] = 9'b111111111;
assign micromatrizz[89][299] = 9'b111111111;
assign micromatrizz[89][300] = 9'b111111111;
assign micromatrizz[89][301] = 9'b111111111;
assign micromatrizz[89][302] = 9'b111111111;
assign micromatrizz[89][303] = 9'b111111111;
assign micromatrizz[89][304] = 9'b111111111;
assign micromatrizz[89][305] = 9'b111111111;
assign micromatrizz[89][306] = 9'b111111111;
assign micromatrizz[89][307] = 9'b111111111;
assign micromatrizz[89][308] = 9'b111111111;
assign micromatrizz[89][309] = 9'b111111111;
assign micromatrizz[89][310] = 9'b111111111;
assign micromatrizz[89][311] = 9'b111111111;
assign micromatrizz[89][312] = 9'b111111111;
assign micromatrizz[89][313] = 9'b111111111;
assign micromatrizz[89][314] = 9'b111111111;
assign micromatrizz[89][315] = 9'b111111111;
assign micromatrizz[89][316] = 9'b111111111;
assign micromatrizz[89][317] = 9'b111111111;
assign micromatrizz[89][318] = 9'b111111111;
assign micromatrizz[89][319] = 9'b111111111;
assign micromatrizz[89][320] = 9'b111111111;
assign micromatrizz[89][321] = 9'b111111111;
assign micromatrizz[89][322] = 9'b111111111;
assign micromatrizz[89][323] = 9'b111111111;
assign micromatrizz[89][324] = 9'b111111111;
assign micromatrizz[89][325] = 9'b111111111;
assign micromatrizz[89][326] = 9'b111111111;
assign micromatrizz[89][327] = 9'b111111111;
assign micromatrizz[89][328] = 9'b111111111;
assign micromatrizz[89][329] = 9'b111111111;
assign micromatrizz[89][330] = 9'b111111111;
assign micromatrizz[89][331] = 9'b111111111;
assign micromatrizz[89][332] = 9'b111111111;
assign micromatrizz[89][333] = 9'b111111111;
assign micromatrizz[89][334] = 9'b111111111;
assign micromatrizz[89][335] = 9'b111111111;
assign micromatrizz[89][336] = 9'b111111111;
assign micromatrizz[89][337] = 9'b111111111;
assign micromatrizz[89][338] = 9'b111111111;
assign micromatrizz[89][339] = 9'b111111111;
assign micromatrizz[89][340] = 9'b111111111;
assign micromatrizz[89][341] = 9'b111111111;
assign micromatrizz[89][342] = 9'b111111111;
assign micromatrizz[89][343] = 9'b111111111;
assign micromatrizz[89][344] = 9'b111111111;
assign micromatrizz[89][345] = 9'b111111111;
assign micromatrizz[89][346] = 9'b111111111;
assign micromatrizz[89][347] = 9'b111111111;
assign micromatrizz[89][348] = 9'b111111111;
assign micromatrizz[89][349] = 9'b111111111;
assign micromatrizz[89][350] = 9'b111111111;
assign micromatrizz[89][351] = 9'b111111111;
assign micromatrizz[89][352] = 9'b111111111;
assign micromatrizz[89][353] = 9'b111111111;
assign micromatrizz[89][354] = 9'b111111111;
assign micromatrizz[89][355] = 9'b111111111;
assign micromatrizz[89][356] = 9'b111111111;
assign micromatrizz[89][357] = 9'b111111111;
assign micromatrizz[89][358] = 9'b111111111;
assign micromatrizz[89][359] = 9'b111111111;
assign micromatrizz[89][360] = 9'b111111111;
assign micromatrizz[89][361] = 9'b111111111;
assign micromatrizz[89][362] = 9'b111111111;
assign micromatrizz[89][363] = 9'b111111111;
assign micromatrizz[89][364] = 9'b111111111;
assign micromatrizz[89][365] = 9'b111111111;
assign micromatrizz[89][366] = 9'b111111111;
assign micromatrizz[89][367] = 9'b111111111;
assign micromatrizz[89][368] = 9'b111111111;
assign micromatrizz[89][369] = 9'b111111111;
assign micromatrizz[89][370] = 9'b111111111;
assign micromatrizz[89][371] = 9'b111111111;
assign micromatrizz[89][372] = 9'b111111111;
assign micromatrizz[89][373] = 9'b111111111;
assign micromatrizz[89][374] = 9'b111111111;
assign micromatrizz[89][375] = 9'b111111111;
assign micromatrizz[89][376] = 9'b111111111;
assign micromatrizz[89][377] = 9'b111111111;
assign micromatrizz[89][378] = 9'b111111111;
assign micromatrizz[89][379] = 9'b111111111;
assign micromatrizz[89][380] = 9'b111111111;
assign micromatrizz[89][381] = 9'b111111111;
assign micromatrizz[89][382] = 9'b111111111;
assign micromatrizz[89][383] = 9'b111111111;
assign micromatrizz[89][384] = 9'b111111111;
assign micromatrizz[89][385] = 9'b111111111;
assign micromatrizz[89][386] = 9'b111111111;
assign micromatrizz[89][387] = 9'b111111111;
assign micromatrizz[89][388] = 9'b111111111;
assign micromatrizz[89][389] = 9'b111111111;
assign micromatrizz[89][390] = 9'b111111111;
assign micromatrizz[89][391] = 9'b111111111;
assign micromatrizz[89][392] = 9'b111111111;
assign micromatrizz[89][393] = 9'b111111111;
assign micromatrizz[89][394] = 9'b111111111;
assign micromatrizz[89][395] = 9'b111111111;
assign micromatrizz[89][396] = 9'b111111111;
assign micromatrizz[89][397] = 9'b111111111;
assign micromatrizz[89][398] = 9'b111111111;
assign micromatrizz[89][399] = 9'b111111111;
assign micromatrizz[89][400] = 9'b111111111;
assign micromatrizz[89][401] = 9'b111111111;
assign micromatrizz[89][402] = 9'b111111111;
assign micromatrizz[89][403] = 9'b111111111;
assign micromatrizz[89][404] = 9'b111111111;
assign micromatrizz[89][405] = 9'b111111111;
assign micromatrizz[89][406] = 9'b111111111;
assign micromatrizz[89][407] = 9'b111111111;
assign micromatrizz[89][408] = 9'b111111111;
assign micromatrizz[89][409] = 9'b111111111;
assign micromatrizz[89][410] = 9'b111111111;
assign micromatrizz[89][411] = 9'b111111111;
assign micromatrizz[89][412] = 9'b111111111;
assign micromatrizz[89][413] = 9'b111111111;
assign micromatrizz[89][414] = 9'b111111111;
assign micromatrizz[89][415] = 9'b111111111;
assign micromatrizz[89][416] = 9'b111111111;
assign micromatrizz[89][417] = 9'b111111111;
assign micromatrizz[89][418] = 9'b111111111;
assign micromatrizz[89][419] = 9'b111111111;
assign micromatrizz[89][420] = 9'b111111111;
assign micromatrizz[89][421] = 9'b111111111;
assign micromatrizz[89][422] = 9'b111111111;
assign micromatrizz[89][423] = 9'b111111111;
assign micromatrizz[89][424] = 9'b111111111;
assign micromatrizz[89][425] = 9'b111111111;
assign micromatrizz[89][426] = 9'b111111111;
assign micromatrizz[89][427] = 9'b111111111;
assign micromatrizz[89][428] = 9'b111111111;
assign micromatrizz[89][429] = 9'b111111111;
assign micromatrizz[89][430] = 9'b111111111;
assign micromatrizz[89][431] = 9'b111111111;
assign micromatrizz[89][432] = 9'b111111111;
assign micromatrizz[89][433] = 9'b111111111;
assign micromatrizz[89][434] = 9'b111111111;
assign micromatrizz[89][435] = 9'b111111111;
assign micromatrizz[89][436] = 9'b111111111;
assign micromatrizz[89][437] = 9'b111111111;
assign micromatrizz[89][438] = 9'b111111111;
assign micromatrizz[89][439] = 9'b111111111;
assign micromatrizz[89][440] = 9'b111111111;
assign micromatrizz[89][441] = 9'b111111111;
assign micromatrizz[89][442] = 9'b111111111;
assign micromatrizz[89][443] = 9'b111111111;
assign micromatrizz[89][444] = 9'b111111111;
assign micromatrizz[89][445] = 9'b111111111;
assign micromatrizz[89][446] = 9'b111111111;
assign micromatrizz[89][447] = 9'b111111111;
assign micromatrizz[89][448] = 9'b111111111;
assign micromatrizz[89][449] = 9'b111111111;
assign micromatrizz[89][450] = 9'b111111111;
assign micromatrizz[89][451] = 9'b111111111;
assign micromatrizz[89][452] = 9'b111111111;
assign micromatrizz[89][453] = 9'b111111111;
assign micromatrizz[89][454] = 9'b111111111;
assign micromatrizz[89][455] = 9'b111111111;
assign micromatrizz[89][456] = 9'b111111111;
assign micromatrizz[89][457] = 9'b111111111;
assign micromatrizz[89][458] = 9'b111111111;
assign micromatrizz[89][459] = 9'b111111111;
assign micromatrizz[89][460] = 9'b111111111;
assign micromatrizz[89][461] = 9'b111111111;
assign micromatrizz[89][462] = 9'b111111111;
assign micromatrizz[89][463] = 9'b111111111;
assign micromatrizz[89][464] = 9'b111111111;
assign micromatrizz[89][465] = 9'b111111111;
assign micromatrizz[89][466] = 9'b111111111;
assign micromatrizz[89][467] = 9'b111111111;
assign micromatrizz[89][468] = 9'b111111111;
assign micromatrizz[89][469] = 9'b111111111;
assign micromatrizz[89][470] = 9'b111111111;
assign micromatrizz[89][471] = 9'b111111111;
assign micromatrizz[89][472] = 9'b111111111;
assign micromatrizz[89][473] = 9'b111111111;
assign micromatrizz[89][474] = 9'b111111111;
assign micromatrizz[89][475] = 9'b111111111;
assign micromatrizz[89][476] = 9'b111111111;
assign micromatrizz[89][477] = 9'b111111111;
assign micromatrizz[89][478] = 9'b111111111;
assign micromatrizz[89][479] = 9'b111111111;
assign micromatrizz[89][480] = 9'b111111111;
assign micromatrizz[89][481] = 9'b111111111;
assign micromatrizz[89][482] = 9'b111111111;
assign micromatrizz[89][483] = 9'b111111111;
assign micromatrizz[89][484] = 9'b111111111;
assign micromatrizz[89][485] = 9'b111111111;
assign micromatrizz[89][486] = 9'b111111111;
assign micromatrizz[89][487] = 9'b111111111;
assign micromatrizz[89][488] = 9'b111111111;
assign micromatrizz[89][489] = 9'b111111111;
assign micromatrizz[89][490] = 9'b111111111;
assign micromatrizz[89][491] = 9'b111111111;
assign micromatrizz[89][492] = 9'b111111111;
assign micromatrizz[89][493] = 9'b111111111;
assign micromatrizz[89][494] = 9'b111111111;
assign micromatrizz[89][495] = 9'b111111111;
assign micromatrizz[89][496] = 9'b111111111;
assign micromatrizz[89][497] = 9'b111111111;
assign micromatrizz[89][498] = 9'b111111111;
assign micromatrizz[89][499] = 9'b111111111;
assign micromatrizz[89][500] = 9'b111111111;
assign micromatrizz[89][501] = 9'b111111111;
assign micromatrizz[89][502] = 9'b111111111;
assign micromatrizz[89][503] = 9'b111111111;
assign micromatrizz[89][504] = 9'b111111111;
assign micromatrizz[89][505] = 9'b111111111;
assign micromatrizz[89][506] = 9'b111111111;
assign micromatrizz[89][507] = 9'b111111111;
assign micromatrizz[89][508] = 9'b111111111;
assign micromatrizz[89][509] = 9'b111111111;
assign micromatrizz[89][510] = 9'b111111111;
assign micromatrizz[89][511] = 9'b111111111;
assign micromatrizz[89][512] = 9'b111111111;
assign micromatrizz[89][513] = 9'b111111111;
assign micromatrizz[89][514] = 9'b111111111;
assign micromatrizz[89][515] = 9'b111111111;
assign micromatrizz[89][516] = 9'b111111111;
assign micromatrizz[89][517] = 9'b111111111;
assign micromatrizz[89][518] = 9'b111111111;
assign micromatrizz[89][519] = 9'b111111111;
assign micromatrizz[89][520] = 9'b111111111;
assign micromatrizz[89][521] = 9'b111111111;
assign micromatrizz[89][522] = 9'b111111111;
assign micromatrizz[89][523] = 9'b111111111;
assign micromatrizz[89][524] = 9'b111111111;
assign micromatrizz[89][525] = 9'b111111111;
assign micromatrizz[89][526] = 9'b111111111;
assign micromatrizz[89][527] = 9'b111111111;
assign micromatrizz[89][528] = 9'b111111111;
assign micromatrizz[89][529] = 9'b111111111;
assign micromatrizz[89][530] = 9'b111111111;
assign micromatrizz[89][531] = 9'b111111111;
assign micromatrizz[89][532] = 9'b111111111;
assign micromatrizz[89][533] = 9'b111111111;
assign micromatrizz[89][534] = 9'b111111111;
assign micromatrizz[89][535] = 9'b111111111;
assign micromatrizz[89][536] = 9'b111111111;
assign micromatrizz[89][537] = 9'b111111111;
assign micromatrizz[89][538] = 9'b111111111;
assign micromatrizz[89][539] = 9'b111111111;
assign micromatrizz[89][540] = 9'b111111111;
assign micromatrizz[89][541] = 9'b111111111;
assign micromatrizz[89][542] = 9'b111111111;
assign micromatrizz[89][543] = 9'b111111111;
assign micromatrizz[89][544] = 9'b111111111;
assign micromatrizz[89][545] = 9'b111111111;
assign micromatrizz[89][546] = 9'b111111111;
assign micromatrizz[89][547] = 9'b111111111;
assign micromatrizz[89][548] = 9'b111111111;
assign micromatrizz[89][549] = 9'b111111111;
assign micromatrizz[89][550] = 9'b111111111;
assign micromatrizz[89][551] = 9'b111111111;
assign micromatrizz[89][552] = 9'b111111111;
assign micromatrizz[89][553] = 9'b111111111;
assign micromatrizz[89][554] = 9'b111111111;
assign micromatrizz[89][555] = 9'b111111111;
assign micromatrizz[89][556] = 9'b111111111;
assign micromatrizz[89][557] = 9'b111111111;
assign micromatrizz[89][558] = 9'b111111111;
assign micromatrizz[89][559] = 9'b111111111;
assign micromatrizz[89][560] = 9'b111111111;
assign micromatrizz[89][561] = 9'b111111111;
assign micromatrizz[89][562] = 9'b111111111;
assign micromatrizz[89][563] = 9'b111111111;
assign micromatrizz[89][564] = 9'b111111111;
assign micromatrizz[89][565] = 9'b111111111;
assign micromatrizz[89][566] = 9'b111111111;
assign micromatrizz[89][567] = 9'b111111111;
assign micromatrizz[89][568] = 9'b111111111;
assign micromatrizz[89][569] = 9'b111111111;
assign micromatrizz[89][570] = 9'b111111111;
assign micromatrizz[89][571] = 9'b111111111;
assign micromatrizz[89][572] = 9'b111111111;
assign micromatrizz[89][573] = 9'b111111111;
assign micromatrizz[89][574] = 9'b111111111;
assign micromatrizz[89][575] = 9'b111111111;
assign micromatrizz[89][576] = 9'b111111111;
assign micromatrizz[89][577] = 9'b111111111;
assign micromatrizz[89][578] = 9'b111111111;
assign micromatrizz[89][579] = 9'b111111111;
assign micromatrizz[89][580] = 9'b111111111;
assign micromatrizz[89][581] = 9'b111111111;
assign micromatrizz[89][582] = 9'b111111111;
assign micromatrizz[89][583] = 9'b111111111;
assign micromatrizz[89][584] = 9'b111111111;
assign micromatrizz[89][585] = 9'b111111111;
assign micromatrizz[89][586] = 9'b111111111;
assign micromatrizz[89][587] = 9'b111111111;
assign micromatrizz[89][588] = 9'b111111111;
assign micromatrizz[89][589] = 9'b111111111;
assign micromatrizz[89][590] = 9'b111111111;
assign micromatrizz[89][591] = 9'b111111111;
assign micromatrizz[89][592] = 9'b111111111;
assign micromatrizz[89][593] = 9'b111111111;
assign micromatrizz[89][594] = 9'b111111111;
assign micromatrizz[89][595] = 9'b111111111;
assign micromatrizz[89][596] = 9'b111111111;
assign micromatrizz[89][597] = 9'b111111111;
assign micromatrizz[89][598] = 9'b111111111;
assign micromatrizz[89][599] = 9'b111111111;
assign micromatrizz[89][600] = 9'b111111111;
assign micromatrizz[89][601] = 9'b111111111;
assign micromatrizz[89][602] = 9'b111111111;
assign micromatrizz[89][603] = 9'b111111111;
assign micromatrizz[89][604] = 9'b111111111;
assign micromatrizz[89][605] = 9'b111111111;
assign micromatrizz[89][606] = 9'b111111111;
assign micromatrizz[89][607] = 9'b111111111;
assign micromatrizz[89][608] = 9'b111111111;
assign micromatrizz[89][609] = 9'b111111111;
assign micromatrizz[89][610] = 9'b111111111;
assign micromatrizz[89][611] = 9'b111111111;
assign micromatrizz[89][612] = 9'b111111111;
assign micromatrizz[89][613] = 9'b111111111;
assign micromatrizz[89][614] = 9'b111111111;
assign micromatrizz[89][615] = 9'b111111111;
assign micromatrizz[89][616] = 9'b111111111;
assign micromatrizz[89][617] = 9'b111111111;
assign micromatrizz[89][618] = 9'b111111111;
assign micromatrizz[89][619] = 9'b111111111;
assign micromatrizz[89][620] = 9'b111111111;
assign micromatrizz[89][621] = 9'b111111111;
assign micromatrizz[89][622] = 9'b111111111;
assign micromatrizz[89][623] = 9'b111111111;
assign micromatrizz[89][624] = 9'b111111111;
assign micromatrizz[89][625] = 9'b111111111;
assign micromatrizz[89][626] = 9'b111111111;
assign micromatrizz[89][627] = 9'b111111111;
assign micromatrizz[89][628] = 9'b111111111;
assign micromatrizz[89][629] = 9'b111111111;
assign micromatrizz[89][630] = 9'b111111111;
assign micromatrizz[89][631] = 9'b111111111;
assign micromatrizz[89][632] = 9'b111111111;
assign micromatrizz[89][633] = 9'b111111111;
assign micromatrizz[89][634] = 9'b111111111;
assign micromatrizz[89][635] = 9'b111111111;
assign micromatrizz[89][636] = 9'b111111111;
assign micromatrizz[89][637] = 9'b111111111;
assign micromatrizz[89][638] = 9'b111111111;
assign micromatrizz[89][639] = 9'b111111111;
assign micromatrizz[90][0] = 9'b111111111;
assign micromatrizz[90][1] = 9'b111111111;
assign micromatrizz[90][2] = 9'b111111111;
assign micromatrizz[90][3] = 9'b111111111;
assign micromatrizz[90][4] = 9'b111111111;
assign micromatrizz[90][5] = 9'b111111111;
assign micromatrizz[90][6] = 9'b111111111;
assign micromatrizz[90][7] = 9'b111111111;
assign micromatrizz[90][8] = 9'b111111111;
assign micromatrizz[90][9] = 9'b111111111;
assign micromatrizz[90][10] = 9'b111111111;
assign micromatrizz[90][11] = 9'b111111111;
assign micromatrizz[90][12] = 9'b111111111;
assign micromatrizz[90][13] = 9'b111111111;
assign micromatrizz[90][14] = 9'b111111111;
assign micromatrizz[90][15] = 9'b111111111;
assign micromatrizz[90][16] = 9'b111111111;
assign micromatrizz[90][17] = 9'b111111111;
assign micromatrizz[90][18] = 9'b111111111;
assign micromatrizz[90][19] = 9'b111111111;
assign micromatrizz[90][20] = 9'b111111111;
assign micromatrizz[90][21] = 9'b111111111;
assign micromatrizz[90][22] = 9'b111111111;
assign micromatrizz[90][23] = 9'b111111111;
assign micromatrizz[90][24] = 9'b111111111;
assign micromatrizz[90][25] = 9'b111111111;
assign micromatrizz[90][26] = 9'b111111111;
assign micromatrizz[90][27] = 9'b111111111;
assign micromatrizz[90][28] = 9'b111111111;
assign micromatrizz[90][29] = 9'b111111111;
assign micromatrizz[90][30] = 9'b111111111;
assign micromatrizz[90][31] = 9'b111111111;
assign micromatrizz[90][32] = 9'b111111111;
assign micromatrizz[90][33] = 9'b111111111;
assign micromatrizz[90][34] = 9'b111111111;
assign micromatrizz[90][35] = 9'b111111111;
assign micromatrizz[90][36] = 9'b111111111;
assign micromatrizz[90][37] = 9'b111111111;
assign micromatrizz[90][38] = 9'b111111111;
assign micromatrizz[90][39] = 9'b111111111;
assign micromatrizz[90][40] = 9'b111111111;
assign micromatrizz[90][41] = 9'b111111111;
assign micromatrizz[90][42] = 9'b111111111;
assign micromatrizz[90][43] = 9'b111111111;
assign micromatrizz[90][44] = 9'b111111111;
assign micromatrizz[90][45] = 9'b111111111;
assign micromatrizz[90][46] = 9'b111111111;
assign micromatrizz[90][47] = 9'b111111111;
assign micromatrizz[90][48] = 9'b111111111;
assign micromatrizz[90][49] = 9'b111111111;
assign micromatrizz[90][50] = 9'b111111111;
assign micromatrizz[90][51] = 9'b111111111;
assign micromatrizz[90][52] = 9'b111111111;
assign micromatrizz[90][53] = 9'b111111111;
assign micromatrizz[90][54] = 9'b111111111;
assign micromatrizz[90][55] = 9'b111111111;
assign micromatrizz[90][56] = 9'b111111111;
assign micromatrizz[90][57] = 9'b111111111;
assign micromatrizz[90][58] = 9'b111111111;
assign micromatrizz[90][59] = 9'b111111111;
assign micromatrizz[90][60] = 9'b111111111;
assign micromatrizz[90][61] = 9'b111111111;
assign micromatrizz[90][62] = 9'b111111111;
assign micromatrizz[90][63] = 9'b111111111;
assign micromatrizz[90][64] = 9'b111111111;
assign micromatrizz[90][65] = 9'b111111111;
assign micromatrizz[90][66] = 9'b111111111;
assign micromatrizz[90][67] = 9'b111111111;
assign micromatrizz[90][68] = 9'b111111111;
assign micromatrizz[90][69] = 9'b111111111;
assign micromatrizz[90][70] = 9'b111111111;
assign micromatrizz[90][71] = 9'b111111111;
assign micromatrizz[90][72] = 9'b111111111;
assign micromatrizz[90][73] = 9'b111111111;
assign micromatrizz[90][74] = 9'b111111111;
assign micromatrizz[90][75] = 9'b111111111;
assign micromatrizz[90][76] = 9'b111111111;
assign micromatrizz[90][77] = 9'b111111111;
assign micromatrizz[90][78] = 9'b111111111;
assign micromatrizz[90][79] = 9'b111111111;
assign micromatrizz[90][80] = 9'b111111111;
assign micromatrizz[90][81] = 9'b111111111;
assign micromatrizz[90][82] = 9'b111111111;
assign micromatrizz[90][83] = 9'b111111111;
assign micromatrizz[90][84] = 9'b111111111;
assign micromatrizz[90][85] = 9'b111111111;
assign micromatrizz[90][86] = 9'b111111111;
assign micromatrizz[90][87] = 9'b111111111;
assign micromatrizz[90][88] = 9'b111111111;
assign micromatrizz[90][89] = 9'b111111111;
assign micromatrizz[90][90] = 9'b111111111;
assign micromatrizz[90][91] = 9'b111111111;
assign micromatrizz[90][92] = 9'b111111111;
assign micromatrizz[90][93] = 9'b111111111;
assign micromatrizz[90][94] = 9'b111111111;
assign micromatrizz[90][95] = 9'b111111111;
assign micromatrizz[90][96] = 9'b111111111;
assign micromatrizz[90][97] = 9'b111111111;
assign micromatrizz[90][98] = 9'b111111111;
assign micromatrizz[90][99] = 9'b111111111;
assign micromatrizz[90][100] = 9'b111111111;
assign micromatrizz[90][101] = 9'b111111111;
assign micromatrizz[90][102] = 9'b111111111;
assign micromatrizz[90][103] = 9'b111111111;
assign micromatrizz[90][104] = 9'b111111111;
assign micromatrizz[90][105] = 9'b111111111;
assign micromatrizz[90][106] = 9'b111111111;
assign micromatrizz[90][107] = 9'b111111111;
assign micromatrizz[90][108] = 9'b111111111;
assign micromatrizz[90][109] = 9'b111111111;
assign micromatrizz[90][110] = 9'b111111111;
assign micromatrizz[90][111] = 9'b111111111;
assign micromatrizz[90][112] = 9'b111111111;
assign micromatrizz[90][113] = 9'b111111111;
assign micromatrizz[90][114] = 9'b111111111;
assign micromatrizz[90][115] = 9'b111111111;
assign micromatrizz[90][116] = 9'b111111111;
assign micromatrizz[90][117] = 9'b111111111;
assign micromatrizz[90][118] = 9'b111111111;
assign micromatrizz[90][119] = 9'b111111111;
assign micromatrizz[90][120] = 9'b111111111;
assign micromatrizz[90][121] = 9'b111111111;
assign micromatrizz[90][122] = 9'b111111111;
assign micromatrizz[90][123] = 9'b111111111;
assign micromatrizz[90][124] = 9'b111111111;
assign micromatrizz[90][125] = 9'b111111111;
assign micromatrizz[90][126] = 9'b111111111;
assign micromatrizz[90][127] = 9'b111111111;
assign micromatrizz[90][128] = 9'b111111111;
assign micromatrizz[90][129] = 9'b111111111;
assign micromatrizz[90][130] = 9'b111111111;
assign micromatrizz[90][131] = 9'b111111111;
assign micromatrizz[90][132] = 9'b111111111;
assign micromatrizz[90][133] = 9'b111111111;
assign micromatrizz[90][134] = 9'b111111111;
assign micromatrizz[90][135] = 9'b111111111;
assign micromatrizz[90][136] = 9'b111111111;
assign micromatrizz[90][137] = 9'b111111111;
assign micromatrizz[90][138] = 9'b111111111;
assign micromatrizz[90][139] = 9'b111111111;
assign micromatrizz[90][140] = 9'b111111111;
assign micromatrizz[90][141] = 9'b111111111;
assign micromatrizz[90][142] = 9'b111111111;
assign micromatrizz[90][143] = 9'b111111111;
assign micromatrizz[90][144] = 9'b111111111;
assign micromatrizz[90][145] = 9'b111111111;
assign micromatrizz[90][146] = 9'b111111111;
assign micromatrizz[90][147] = 9'b111111111;
assign micromatrizz[90][148] = 9'b111111111;
assign micromatrizz[90][149] = 9'b111111111;
assign micromatrizz[90][150] = 9'b111111111;
assign micromatrizz[90][151] = 9'b111111111;
assign micromatrizz[90][152] = 9'b111111111;
assign micromatrizz[90][153] = 9'b111111111;
assign micromatrizz[90][154] = 9'b111111111;
assign micromatrizz[90][155] = 9'b111111111;
assign micromatrizz[90][156] = 9'b111111111;
assign micromatrizz[90][157] = 9'b111111111;
assign micromatrizz[90][158] = 9'b111111111;
assign micromatrizz[90][159] = 9'b111111111;
assign micromatrizz[90][160] = 9'b111111111;
assign micromatrizz[90][161] = 9'b111111111;
assign micromatrizz[90][162] = 9'b111111111;
assign micromatrizz[90][163] = 9'b111111111;
assign micromatrizz[90][164] = 9'b111111111;
assign micromatrizz[90][165] = 9'b111111111;
assign micromatrizz[90][166] = 9'b111111111;
assign micromatrizz[90][167] = 9'b111111111;
assign micromatrizz[90][168] = 9'b111111111;
assign micromatrizz[90][169] = 9'b111111111;
assign micromatrizz[90][170] = 9'b111111111;
assign micromatrizz[90][171] = 9'b111111111;
assign micromatrizz[90][172] = 9'b111111111;
assign micromatrizz[90][173] = 9'b111111111;
assign micromatrizz[90][174] = 9'b111111111;
assign micromatrizz[90][175] = 9'b111111111;
assign micromatrizz[90][176] = 9'b111111111;
assign micromatrizz[90][177] = 9'b111111111;
assign micromatrizz[90][178] = 9'b111111111;
assign micromatrizz[90][179] = 9'b111111111;
assign micromatrizz[90][180] = 9'b111111111;
assign micromatrizz[90][181] = 9'b111111111;
assign micromatrizz[90][182] = 9'b111111111;
assign micromatrizz[90][183] = 9'b111111111;
assign micromatrizz[90][184] = 9'b111111111;
assign micromatrizz[90][185] = 9'b111111111;
assign micromatrizz[90][186] = 9'b111111111;
assign micromatrizz[90][187] = 9'b111111111;
assign micromatrizz[90][188] = 9'b111111111;
assign micromatrizz[90][189] = 9'b111111111;
assign micromatrizz[90][190] = 9'b111111111;
assign micromatrizz[90][191] = 9'b111111111;
assign micromatrizz[90][192] = 9'b111111111;
assign micromatrizz[90][193] = 9'b111111111;
assign micromatrizz[90][194] = 9'b111111111;
assign micromatrizz[90][195] = 9'b111111111;
assign micromatrizz[90][196] = 9'b111111111;
assign micromatrizz[90][197] = 9'b111111111;
assign micromatrizz[90][198] = 9'b111111111;
assign micromatrizz[90][199] = 9'b111111111;
assign micromatrizz[90][200] = 9'b111111111;
assign micromatrizz[90][201] = 9'b111111111;
assign micromatrizz[90][202] = 9'b111111111;
assign micromatrizz[90][203] = 9'b111111111;
assign micromatrizz[90][204] = 9'b111111111;
assign micromatrizz[90][205] = 9'b111111111;
assign micromatrizz[90][206] = 9'b111111111;
assign micromatrizz[90][207] = 9'b111111111;
assign micromatrizz[90][208] = 9'b111111111;
assign micromatrizz[90][209] = 9'b111111111;
assign micromatrizz[90][210] = 9'b111111111;
assign micromatrizz[90][211] = 9'b111111111;
assign micromatrizz[90][212] = 9'b111111111;
assign micromatrizz[90][213] = 9'b111111111;
assign micromatrizz[90][214] = 9'b111111111;
assign micromatrizz[90][215] = 9'b111111111;
assign micromatrizz[90][216] = 9'b111111111;
assign micromatrizz[90][217] = 9'b111111111;
assign micromatrizz[90][218] = 9'b111111111;
assign micromatrizz[90][219] = 9'b111111111;
assign micromatrizz[90][220] = 9'b111111111;
assign micromatrizz[90][221] = 9'b111111111;
assign micromatrizz[90][222] = 9'b111111111;
assign micromatrizz[90][223] = 9'b111111111;
assign micromatrizz[90][224] = 9'b111111111;
assign micromatrizz[90][225] = 9'b111111111;
assign micromatrizz[90][226] = 9'b111111111;
assign micromatrizz[90][227] = 9'b111111111;
assign micromatrizz[90][228] = 9'b111111111;
assign micromatrizz[90][229] = 9'b111111111;
assign micromatrizz[90][230] = 9'b111111111;
assign micromatrizz[90][231] = 9'b111111111;
assign micromatrizz[90][232] = 9'b111111111;
assign micromatrizz[90][233] = 9'b111111111;
assign micromatrizz[90][234] = 9'b111111111;
assign micromatrizz[90][235] = 9'b111111111;
assign micromatrizz[90][236] = 9'b111111111;
assign micromatrizz[90][237] = 9'b111111111;
assign micromatrizz[90][238] = 9'b111111111;
assign micromatrizz[90][239] = 9'b111111111;
assign micromatrizz[90][240] = 9'b111111111;
assign micromatrizz[90][241] = 9'b111111111;
assign micromatrizz[90][242] = 9'b111111111;
assign micromatrizz[90][243] = 9'b111111111;
assign micromatrizz[90][244] = 9'b111111111;
assign micromatrizz[90][245] = 9'b111111111;
assign micromatrizz[90][246] = 9'b111111111;
assign micromatrizz[90][247] = 9'b111111111;
assign micromatrizz[90][248] = 9'b111111111;
assign micromatrizz[90][249] = 9'b111111111;
assign micromatrizz[90][250] = 9'b111111111;
assign micromatrizz[90][251] = 9'b111111111;
assign micromatrizz[90][252] = 9'b111111111;
assign micromatrizz[90][253] = 9'b111111111;
assign micromatrizz[90][254] = 9'b111111111;
assign micromatrizz[90][255] = 9'b111111111;
assign micromatrizz[90][256] = 9'b111111111;
assign micromatrizz[90][257] = 9'b111111111;
assign micromatrizz[90][258] = 9'b111111111;
assign micromatrizz[90][259] = 9'b111111111;
assign micromatrizz[90][260] = 9'b111111111;
assign micromatrizz[90][261] = 9'b111111111;
assign micromatrizz[90][262] = 9'b111111111;
assign micromatrizz[90][263] = 9'b111111111;
assign micromatrizz[90][264] = 9'b111111111;
assign micromatrizz[90][265] = 9'b111111111;
assign micromatrizz[90][266] = 9'b111111111;
assign micromatrizz[90][267] = 9'b111111111;
assign micromatrizz[90][268] = 9'b111111111;
assign micromatrizz[90][269] = 9'b111111111;
assign micromatrizz[90][270] = 9'b111111111;
assign micromatrizz[90][271] = 9'b111111111;
assign micromatrizz[90][272] = 9'b111111111;
assign micromatrizz[90][273] = 9'b111111111;
assign micromatrizz[90][274] = 9'b111111111;
assign micromatrizz[90][275] = 9'b111111111;
assign micromatrizz[90][276] = 9'b111111111;
assign micromatrizz[90][277] = 9'b111111111;
assign micromatrizz[90][278] = 9'b111111111;
assign micromatrizz[90][279] = 9'b111111111;
assign micromatrizz[90][280] = 9'b111111111;
assign micromatrizz[90][281] = 9'b111111111;
assign micromatrizz[90][282] = 9'b111111111;
assign micromatrizz[90][283] = 9'b111111111;
assign micromatrizz[90][284] = 9'b111111111;
assign micromatrizz[90][285] = 9'b111111111;
assign micromatrizz[90][286] = 9'b111111111;
assign micromatrizz[90][287] = 9'b111111111;
assign micromatrizz[90][288] = 9'b111111111;
assign micromatrizz[90][289] = 9'b111111111;
assign micromatrizz[90][290] = 9'b111111111;
assign micromatrizz[90][291] = 9'b111111111;
assign micromatrizz[90][292] = 9'b111111111;
assign micromatrizz[90][293] = 9'b111111111;
assign micromatrizz[90][294] = 9'b111111111;
assign micromatrizz[90][295] = 9'b111111111;
assign micromatrizz[90][296] = 9'b111111111;
assign micromatrizz[90][297] = 9'b111111111;
assign micromatrizz[90][298] = 9'b111111111;
assign micromatrizz[90][299] = 9'b111111111;
assign micromatrizz[90][300] = 9'b111111111;
assign micromatrizz[90][301] = 9'b111111111;
assign micromatrizz[90][302] = 9'b111111111;
assign micromatrizz[90][303] = 9'b111111111;
assign micromatrizz[90][304] = 9'b111111111;
assign micromatrizz[90][305] = 9'b111111111;
assign micromatrizz[90][306] = 9'b111111111;
assign micromatrizz[90][307] = 9'b111111111;
assign micromatrizz[90][308] = 9'b111111111;
assign micromatrizz[90][309] = 9'b111111111;
assign micromatrizz[90][310] = 9'b111111111;
assign micromatrizz[90][311] = 9'b111111111;
assign micromatrizz[90][312] = 9'b111111111;
assign micromatrizz[90][313] = 9'b111111111;
assign micromatrizz[90][314] = 9'b111111111;
assign micromatrizz[90][315] = 9'b111111111;
assign micromatrizz[90][316] = 9'b111111111;
assign micromatrizz[90][317] = 9'b111111111;
assign micromatrizz[90][318] = 9'b111111111;
assign micromatrizz[90][319] = 9'b111111111;
assign micromatrizz[90][320] = 9'b111111111;
assign micromatrizz[90][321] = 9'b111111111;
assign micromatrizz[90][322] = 9'b111111111;
assign micromatrizz[90][323] = 9'b111111111;
assign micromatrizz[90][324] = 9'b111111111;
assign micromatrizz[90][325] = 9'b111111111;
assign micromatrizz[90][326] = 9'b111111111;
assign micromatrizz[90][327] = 9'b111111111;
assign micromatrizz[90][328] = 9'b111111111;
assign micromatrizz[90][329] = 9'b111111111;
assign micromatrizz[90][330] = 9'b111111111;
assign micromatrizz[90][331] = 9'b111111111;
assign micromatrizz[90][332] = 9'b111111111;
assign micromatrizz[90][333] = 9'b111111111;
assign micromatrizz[90][334] = 9'b111111111;
assign micromatrizz[90][335] = 9'b111111111;
assign micromatrizz[90][336] = 9'b111111111;
assign micromatrizz[90][337] = 9'b111111111;
assign micromatrizz[90][338] = 9'b111111111;
assign micromatrizz[90][339] = 9'b111111111;
assign micromatrizz[90][340] = 9'b111111111;
assign micromatrizz[90][341] = 9'b111111111;
assign micromatrizz[90][342] = 9'b111111111;
assign micromatrizz[90][343] = 9'b111111111;
assign micromatrizz[90][344] = 9'b111111111;
assign micromatrizz[90][345] = 9'b111111111;
assign micromatrizz[90][346] = 9'b111111111;
assign micromatrizz[90][347] = 9'b111111111;
assign micromatrizz[90][348] = 9'b111111111;
assign micromatrizz[90][349] = 9'b111111111;
assign micromatrizz[90][350] = 9'b111111111;
assign micromatrizz[90][351] = 9'b111111111;
assign micromatrizz[90][352] = 9'b111111111;
assign micromatrizz[90][353] = 9'b111111111;
assign micromatrizz[90][354] = 9'b111111111;
assign micromatrizz[90][355] = 9'b111111111;
assign micromatrizz[90][356] = 9'b111111111;
assign micromatrizz[90][357] = 9'b111111111;
assign micromatrizz[90][358] = 9'b111111111;
assign micromatrizz[90][359] = 9'b111111111;
assign micromatrizz[90][360] = 9'b111111111;
assign micromatrizz[90][361] = 9'b111111111;
assign micromatrizz[90][362] = 9'b111111111;
assign micromatrizz[90][363] = 9'b111111111;
assign micromatrizz[90][364] = 9'b111111111;
assign micromatrizz[90][365] = 9'b111111111;
assign micromatrizz[90][366] = 9'b111111111;
assign micromatrizz[90][367] = 9'b111111111;
assign micromatrizz[90][368] = 9'b111111111;
assign micromatrizz[90][369] = 9'b111111111;
assign micromatrizz[90][370] = 9'b111111111;
assign micromatrizz[90][371] = 9'b111111111;
assign micromatrizz[90][372] = 9'b111111111;
assign micromatrizz[90][373] = 9'b111111111;
assign micromatrizz[90][374] = 9'b111111111;
assign micromatrizz[90][375] = 9'b111111111;
assign micromatrizz[90][376] = 9'b111111111;
assign micromatrizz[90][377] = 9'b111111111;
assign micromatrizz[90][378] = 9'b111111111;
assign micromatrizz[90][379] = 9'b111111111;
assign micromatrizz[90][380] = 9'b111111111;
assign micromatrizz[90][381] = 9'b111111111;
assign micromatrizz[90][382] = 9'b111111111;
assign micromatrizz[90][383] = 9'b111111111;
assign micromatrizz[90][384] = 9'b111111111;
assign micromatrizz[90][385] = 9'b111111111;
assign micromatrizz[90][386] = 9'b111111111;
assign micromatrizz[90][387] = 9'b111111111;
assign micromatrizz[90][388] = 9'b111111111;
assign micromatrizz[90][389] = 9'b111111111;
assign micromatrizz[90][390] = 9'b111111111;
assign micromatrizz[90][391] = 9'b111111111;
assign micromatrizz[90][392] = 9'b111111111;
assign micromatrizz[90][393] = 9'b111111111;
assign micromatrizz[90][394] = 9'b111111111;
assign micromatrizz[90][395] = 9'b111111111;
assign micromatrizz[90][396] = 9'b111111111;
assign micromatrizz[90][397] = 9'b111111111;
assign micromatrizz[90][398] = 9'b111111111;
assign micromatrizz[90][399] = 9'b111111111;
assign micromatrizz[90][400] = 9'b111111111;
assign micromatrizz[90][401] = 9'b111111111;
assign micromatrizz[90][402] = 9'b111111111;
assign micromatrizz[90][403] = 9'b111111111;
assign micromatrizz[90][404] = 9'b111111111;
assign micromatrizz[90][405] = 9'b111111111;
assign micromatrizz[90][406] = 9'b111111111;
assign micromatrizz[90][407] = 9'b111111111;
assign micromatrizz[90][408] = 9'b111111111;
assign micromatrizz[90][409] = 9'b111111111;
assign micromatrizz[90][410] = 9'b111111111;
assign micromatrizz[90][411] = 9'b111111111;
assign micromatrizz[90][412] = 9'b111111111;
assign micromatrizz[90][413] = 9'b111111111;
assign micromatrizz[90][414] = 9'b111111111;
assign micromatrizz[90][415] = 9'b111111111;
assign micromatrizz[90][416] = 9'b111111111;
assign micromatrizz[90][417] = 9'b111111111;
assign micromatrizz[90][418] = 9'b111111111;
assign micromatrizz[90][419] = 9'b111111111;
assign micromatrizz[90][420] = 9'b111111111;
assign micromatrizz[90][421] = 9'b111111111;
assign micromatrizz[90][422] = 9'b111111111;
assign micromatrizz[90][423] = 9'b111111111;
assign micromatrizz[90][424] = 9'b111111111;
assign micromatrizz[90][425] = 9'b111111111;
assign micromatrizz[90][426] = 9'b111111111;
assign micromatrizz[90][427] = 9'b111111111;
assign micromatrizz[90][428] = 9'b111111111;
assign micromatrizz[90][429] = 9'b111111111;
assign micromatrizz[90][430] = 9'b111111111;
assign micromatrizz[90][431] = 9'b111111111;
assign micromatrizz[90][432] = 9'b111111111;
assign micromatrizz[90][433] = 9'b111111111;
assign micromatrizz[90][434] = 9'b111111111;
assign micromatrizz[90][435] = 9'b111111111;
assign micromatrizz[90][436] = 9'b111111111;
assign micromatrizz[90][437] = 9'b111111111;
assign micromatrizz[90][438] = 9'b111111111;
assign micromatrizz[90][439] = 9'b111111111;
assign micromatrizz[90][440] = 9'b111111111;
assign micromatrizz[90][441] = 9'b111111111;
assign micromatrizz[90][442] = 9'b111111111;
assign micromatrizz[90][443] = 9'b111111111;
assign micromatrizz[90][444] = 9'b111111111;
assign micromatrizz[90][445] = 9'b111111111;
assign micromatrizz[90][446] = 9'b111111111;
assign micromatrizz[90][447] = 9'b111111111;
assign micromatrizz[90][448] = 9'b111111111;
assign micromatrizz[90][449] = 9'b111111111;
assign micromatrizz[90][450] = 9'b111111111;
assign micromatrizz[90][451] = 9'b111111111;
assign micromatrizz[90][452] = 9'b111111111;
assign micromatrizz[90][453] = 9'b111111111;
assign micromatrizz[90][454] = 9'b111111111;
assign micromatrizz[90][455] = 9'b111111111;
assign micromatrizz[90][456] = 9'b111111111;
assign micromatrizz[90][457] = 9'b111111111;
assign micromatrizz[90][458] = 9'b111111111;
assign micromatrizz[90][459] = 9'b111111111;
assign micromatrizz[90][460] = 9'b111111111;
assign micromatrizz[90][461] = 9'b111111111;
assign micromatrizz[90][462] = 9'b111111111;
assign micromatrizz[90][463] = 9'b111111111;
assign micromatrizz[90][464] = 9'b111111111;
assign micromatrizz[90][465] = 9'b111111111;
assign micromatrizz[90][466] = 9'b111111111;
assign micromatrizz[90][467] = 9'b111111111;
assign micromatrizz[90][468] = 9'b111111111;
assign micromatrizz[90][469] = 9'b111111111;
assign micromatrizz[90][470] = 9'b111111111;
assign micromatrizz[90][471] = 9'b111111111;
assign micromatrizz[90][472] = 9'b111111111;
assign micromatrizz[90][473] = 9'b111111111;
assign micromatrizz[90][474] = 9'b111111111;
assign micromatrizz[90][475] = 9'b111111111;
assign micromatrizz[90][476] = 9'b111111111;
assign micromatrizz[90][477] = 9'b111111111;
assign micromatrizz[90][478] = 9'b111111111;
assign micromatrizz[90][479] = 9'b111111111;
assign micromatrizz[90][480] = 9'b111111111;
assign micromatrizz[90][481] = 9'b111111111;
assign micromatrizz[90][482] = 9'b111111111;
assign micromatrizz[90][483] = 9'b111111111;
assign micromatrizz[90][484] = 9'b111111111;
assign micromatrizz[90][485] = 9'b111111111;
assign micromatrizz[90][486] = 9'b111111111;
assign micromatrizz[90][487] = 9'b111111111;
assign micromatrizz[90][488] = 9'b111111111;
assign micromatrizz[90][489] = 9'b111111111;
assign micromatrizz[90][490] = 9'b111111111;
assign micromatrizz[90][491] = 9'b111111111;
assign micromatrizz[90][492] = 9'b111111111;
assign micromatrizz[90][493] = 9'b111111111;
assign micromatrizz[90][494] = 9'b111111111;
assign micromatrizz[90][495] = 9'b111111111;
assign micromatrizz[90][496] = 9'b111111111;
assign micromatrizz[90][497] = 9'b111111111;
assign micromatrizz[90][498] = 9'b111111111;
assign micromatrizz[90][499] = 9'b111111111;
assign micromatrizz[90][500] = 9'b111111111;
assign micromatrizz[90][501] = 9'b111111111;
assign micromatrizz[90][502] = 9'b111111111;
assign micromatrizz[90][503] = 9'b111111111;
assign micromatrizz[90][504] = 9'b111111111;
assign micromatrizz[90][505] = 9'b111111111;
assign micromatrizz[90][506] = 9'b111111111;
assign micromatrizz[90][507] = 9'b111111111;
assign micromatrizz[90][508] = 9'b111111111;
assign micromatrizz[90][509] = 9'b111111111;
assign micromatrizz[90][510] = 9'b111111111;
assign micromatrizz[90][511] = 9'b111111111;
assign micromatrizz[90][512] = 9'b111111111;
assign micromatrizz[90][513] = 9'b111111111;
assign micromatrizz[90][514] = 9'b111111111;
assign micromatrizz[90][515] = 9'b111111111;
assign micromatrizz[90][516] = 9'b111111111;
assign micromatrizz[90][517] = 9'b111111111;
assign micromatrizz[90][518] = 9'b111111111;
assign micromatrizz[90][519] = 9'b111111111;
assign micromatrizz[90][520] = 9'b111111111;
assign micromatrizz[90][521] = 9'b111111111;
assign micromatrizz[90][522] = 9'b111111111;
assign micromatrizz[90][523] = 9'b111111111;
assign micromatrizz[90][524] = 9'b111111111;
assign micromatrizz[90][525] = 9'b111111111;
assign micromatrizz[90][526] = 9'b111111111;
assign micromatrizz[90][527] = 9'b111111111;
assign micromatrizz[90][528] = 9'b111111111;
assign micromatrizz[90][529] = 9'b111111111;
assign micromatrizz[90][530] = 9'b111111111;
assign micromatrizz[90][531] = 9'b111111111;
assign micromatrizz[90][532] = 9'b111111111;
assign micromatrizz[90][533] = 9'b111111111;
assign micromatrizz[90][534] = 9'b111111111;
assign micromatrizz[90][535] = 9'b111111111;
assign micromatrizz[90][536] = 9'b111111111;
assign micromatrizz[90][537] = 9'b111111111;
assign micromatrizz[90][538] = 9'b111111111;
assign micromatrizz[90][539] = 9'b111111111;
assign micromatrizz[90][540] = 9'b111111111;
assign micromatrizz[90][541] = 9'b111111111;
assign micromatrizz[90][542] = 9'b111111111;
assign micromatrizz[90][543] = 9'b111111111;
assign micromatrizz[90][544] = 9'b111111111;
assign micromatrizz[90][545] = 9'b111111111;
assign micromatrizz[90][546] = 9'b111111111;
assign micromatrizz[90][547] = 9'b111111111;
assign micromatrizz[90][548] = 9'b111111111;
assign micromatrizz[90][549] = 9'b111111111;
assign micromatrizz[90][550] = 9'b111111111;
assign micromatrizz[90][551] = 9'b111111111;
assign micromatrizz[90][552] = 9'b111111111;
assign micromatrizz[90][553] = 9'b111111111;
assign micromatrizz[90][554] = 9'b111111111;
assign micromatrizz[90][555] = 9'b111111111;
assign micromatrizz[90][556] = 9'b111111111;
assign micromatrizz[90][557] = 9'b111111111;
assign micromatrizz[90][558] = 9'b111111111;
assign micromatrizz[90][559] = 9'b111111111;
assign micromatrizz[90][560] = 9'b111111111;
assign micromatrizz[90][561] = 9'b111111111;
assign micromatrizz[90][562] = 9'b111111111;
assign micromatrizz[90][563] = 9'b111111111;
assign micromatrizz[90][564] = 9'b111111111;
assign micromatrizz[90][565] = 9'b111111111;
assign micromatrizz[90][566] = 9'b111111111;
assign micromatrizz[90][567] = 9'b111111111;
assign micromatrizz[90][568] = 9'b111111111;
assign micromatrizz[90][569] = 9'b111111111;
assign micromatrizz[90][570] = 9'b111111111;
assign micromatrizz[90][571] = 9'b111111111;
assign micromatrizz[90][572] = 9'b111111111;
assign micromatrizz[90][573] = 9'b111111111;
assign micromatrizz[90][574] = 9'b111111111;
assign micromatrizz[90][575] = 9'b111111111;
assign micromatrizz[90][576] = 9'b111111111;
assign micromatrizz[90][577] = 9'b111111111;
assign micromatrizz[90][578] = 9'b111111111;
assign micromatrizz[90][579] = 9'b111111111;
assign micromatrizz[90][580] = 9'b111111111;
assign micromatrizz[90][581] = 9'b111111111;
assign micromatrizz[90][582] = 9'b111111111;
assign micromatrizz[90][583] = 9'b111111111;
assign micromatrizz[90][584] = 9'b111111111;
assign micromatrizz[90][585] = 9'b111111111;
assign micromatrizz[90][586] = 9'b111111111;
assign micromatrizz[90][587] = 9'b111111111;
assign micromatrizz[90][588] = 9'b111111111;
assign micromatrizz[90][589] = 9'b111111111;
assign micromatrizz[90][590] = 9'b111111111;
assign micromatrizz[90][591] = 9'b111111111;
assign micromatrizz[90][592] = 9'b111111111;
assign micromatrizz[90][593] = 9'b111111111;
assign micromatrizz[90][594] = 9'b111111111;
assign micromatrizz[90][595] = 9'b111111111;
assign micromatrizz[90][596] = 9'b111111111;
assign micromatrizz[90][597] = 9'b111111111;
assign micromatrizz[90][598] = 9'b111111111;
assign micromatrizz[90][599] = 9'b111111111;
assign micromatrizz[90][600] = 9'b111111111;
assign micromatrizz[90][601] = 9'b111111111;
assign micromatrizz[90][602] = 9'b111111111;
assign micromatrizz[90][603] = 9'b111111111;
assign micromatrizz[90][604] = 9'b111111111;
assign micromatrizz[90][605] = 9'b111111111;
assign micromatrizz[90][606] = 9'b111111111;
assign micromatrizz[90][607] = 9'b111111111;
assign micromatrizz[90][608] = 9'b111111111;
assign micromatrizz[90][609] = 9'b111111111;
assign micromatrizz[90][610] = 9'b111111111;
assign micromatrizz[90][611] = 9'b111111111;
assign micromatrizz[90][612] = 9'b111111111;
assign micromatrizz[90][613] = 9'b111111111;
assign micromatrizz[90][614] = 9'b111111111;
assign micromatrizz[90][615] = 9'b111111111;
assign micromatrizz[90][616] = 9'b111111111;
assign micromatrizz[90][617] = 9'b111111111;
assign micromatrizz[90][618] = 9'b111111111;
assign micromatrizz[90][619] = 9'b111111111;
assign micromatrizz[90][620] = 9'b111111111;
assign micromatrizz[90][621] = 9'b111111111;
assign micromatrizz[90][622] = 9'b111111111;
assign micromatrizz[90][623] = 9'b111111111;
assign micromatrizz[90][624] = 9'b111111111;
assign micromatrizz[90][625] = 9'b111111111;
assign micromatrizz[90][626] = 9'b111111111;
assign micromatrizz[90][627] = 9'b111111111;
assign micromatrizz[90][628] = 9'b111111111;
assign micromatrizz[90][629] = 9'b111111111;
assign micromatrizz[90][630] = 9'b111111111;
assign micromatrizz[90][631] = 9'b111111111;
assign micromatrizz[90][632] = 9'b111111111;
assign micromatrizz[90][633] = 9'b111111111;
assign micromatrizz[90][634] = 9'b111111111;
assign micromatrizz[90][635] = 9'b111111111;
assign micromatrizz[90][636] = 9'b111111111;
assign micromatrizz[90][637] = 9'b111111111;
assign micromatrizz[90][638] = 9'b111111111;
assign micromatrizz[90][639] = 9'b111111111;
assign micromatrizz[91][0] = 9'b111111111;
assign micromatrizz[91][1] = 9'b111111111;
assign micromatrizz[91][2] = 9'b111111111;
assign micromatrizz[91][3] = 9'b111111111;
assign micromatrizz[91][4] = 9'b111111111;
assign micromatrizz[91][5] = 9'b111111111;
assign micromatrizz[91][6] = 9'b111111111;
assign micromatrizz[91][7] = 9'b111111111;
assign micromatrizz[91][8] = 9'b111111111;
assign micromatrizz[91][9] = 9'b111111111;
assign micromatrizz[91][10] = 9'b111111111;
assign micromatrizz[91][11] = 9'b111111111;
assign micromatrizz[91][12] = 9'b111111111;
assign micromatrizz[91][13] = 9'b111111111;
assign micromatrizz[91][14] = 9'b111111111;
assign micromatrizz[91][15] = 9'b111111111;
assign micromatrizz[91][16] = 9'b111111111;
assign micromatrizz[91][17] = 9'b111111111;
assign micromatrizz[91][18] = 9'b111111111;
assign micromatrizz[91][19] = 9'b111111111;
assign micromatrizz[91][20] = 9'b111111111;
assign micromatrizz[91][21] = 9'b111111111;
assign micromatrizz[91][22] = 9'b111111111;
assign micromatrizz[91][23] = 9'b111111111;
assign micromatrizz[91][24] = 9'b111111111;
assign micromatrizz[91][25] = 9'b111111111;
assign micromatrizz[91][26] = 9'b111111111;
assign micromatrizz[91][27] = 9'b111111111;
assign micromatrizz[91][28] = 9'b111111111;
assign micromatrizz[91][29] = 9'b111111111;
assign micromatrizz[91][30] = 9'b111111111;
assign micromatrizz[91][31] = 9'b111111111;
assign micromatrizz[91][32] = 9'b111111111;
assign micromatrizz[91][33] = 9'b111111111;
assign micromatrizz[91][34] = 9'b111111111;
assign micromatrizz[91][35] = 9'b111111111;
assign micromatrizz[91][36] = 9'b111111111;
assign micromatrizz[91][37] = 9'b111111111;
assign micromatrizz[91][38] = 9'b111111111;
assign micromatrizz[91][39] = 9'b111111111;
assign micromatrizz[91][40] = 9'b111111111;
assign micromatrizz[91][41] = 9'b111111111;
assign micromatrizz[91][42] = 9'b111111111;
assign micromatrizz[91][43] = 9'b111111111;
assign micromatrizz[91][44] = 9'b111111111;
assign micromatrizz[91][45] = 9'b111111111;
assign micromatrizz[91][46] = 9'b111111111;
assign micromatrizz[91][47] = 9'b111111111;
assign micromatrizz[91][48] = 9'b111111111;
assign micromatrizz[91][49] = 9'b111111111;
assign micromatrizz[91][50] = 9'b111111111;
assign micromatrizz[91][51] = 9'b111111111;
assign micromatrizz[91][52] = 9'b111111111;
assign micromatrizz[91][53] = 9'b111111111;
assign micromatrizz[91][54] = 9'b111111111;
assign micromatrizz[91][55] = 9'b111111111;
assign micromatrizz[91][56] = 9'b111111111;
assign micromatrizz[91][57] = 9'b111111111;
assign micromatrizz[91][58] = 9'b111111111;
assign micromatrizz[91][59] = 9'b111111111;
assign micromatrizz[91][60] = 9'b111111111;
assign micromatrizz[91][61] = 9'b111111111;
assign micromatrizz[91][62] = 9'b111111111;
assign micromatrizz[91][63] = 9'b111111111;
assign micromatrizz[91][64] = 9'b111111111;
assign micromatrizz[91][65] = 9'b111111111;
assign micromatrizz[91][66] = 9'b111111111;
assign micromatrizz[91][67] = 9'b111111111;
assign micromatrizz[91][68] = 9'b111111111;
assign micromatrizz[91][69] = 9'b111111111;
assign micromatrizz[91][70] = 9'b111111111;
assign micromatrizz[91][71] = 9'b111111111;
assign micromatrizz[91][72] = 9'b111111111;
assign micromatrizz[91][73] = 9'b111111111;
assign micromatrizz[91][74] = 9'b111111111;
assign micromatrizz[91][75] = 9'b111111111;
assign micromatrizz[91][76] = 9'b111111111;
assign micromatrizz[91][77] = 9'b111111111;
assign micromatrizz[91][78] = 9'b111111111;
assign micromatrizz[91][79] = 9'b111111111;
assign micromatrizz[91][80] = 9'b111111111;
assign micromatrizz[91][81] = 9'b111111111;
assign micromatrizz[91][82] = 9'b111111111;
assign micromatrizz[91][83] = 9'b111111111;
assign micromatrizz[91][84] = 9'b111111111;
assign micromatrizz[91][85] = 9'b111111111;
assign micromatrizz[91][86] = 9'b111111111;
assign micromatrizz[91][87] = 9'b111111111;
assign micromatrizz[91][88] = 9'b111111111;
assign micromatrizz[91][89] = 9'b111111111;
assign micromatrizz[91][90] = 9'b111111111;
assign micromatrizz[91][91] = 9'b111111111;
assign micromatrizz[91][92] = 9'b111111111;
assign micromatrizz[91][93] = 9'b111111111;
assign micromatrizz[91][94] = 9'b111111111;
assign micromatrizz[91][95] = 9'b111111111;
assign micromatrizz[91][96] = 9'b111111111;
assign micromatrizz[91][97] = 9'b111111111;
assign micromatrizz[91][98] = 9'b111111111;
assign micromatrizz[91][99] = 9'b111111111;
assign micromatrizz[91][100] = 9'b111111111;
assign micromatrizz[91][101] = 9'b111111111;
assign micromatrizz[91][102] = 9'b111111111;
assign micromatrizz[91][103] = 9'b111111111;
assign micromatrizz[91][104] = 9'b111111111;
assign micromatrizz[91][105] = 9'b111111111;
assign micromatrizz[91][106] = 9'b111111111;
assign micromatrizz[91][107] = 9'b111111111;
assign micromatrizz[91][108] = 9'b111111111;
assign micromatrizz[91][109] = 9'b111111111;
assign micromatrizz[91][110] = 9'b111111111;
assign micromatrizz[91][111] = 9'b111111111;
assign micromatrizz[91][112] = 9'b111111111;
assign micromatrizz[91][113] = 9'b111111111;
assign micromatrizz[91][114] = 9'b111111111;
assign micromatrizz[91][115] = 9'b111111111;
assign micromatrizz[91][116] = 9'b111111111;
assign micromatrizz[91][117] = 9'b111111111;
assign micromatrizz[91][118] = 9'b111111111;
assign micromatrizz[91][119] = 9'b111111111;
assign micromatrizz[91][120] = 9'b111111111;
assign micromatrizz[91][121] = 9'b111111111;
assign micromatrizz[91][122] = 9'b111111111;
assign micromatrizz[91][123] = 9'b111111111;
assign micromatrizz[91][124] = 9'b111111111;
assign micromatrizz[91][125] = 9'b111111111;
assign micromatrizz[91][126] = 9'b111111111;
assign micromatrizz[91][127] = 9'b111111111;
assign micromatrizz[91][128] = 9'b111111111;
assign micromatrizz[91][129] = 9'b111111111;
assign micromatrizz[91][130] = 9'b111111111;
assign micromatrizz[91][131] = 9'b111111111;
assign micromatrizz[91][132] = 9'b111111111;
assign micromatrizz[91][133] = 9'b111111111;
assign micromatrizz[91][134] = 9'b111111111;
assign micromatrizz[91][135] = 9'b111111111;
assign micromatrizz[91][136] = 9'b111111111;
assign micromatrizz[91][137] = 9'b111111111;
assign micromatrizz[91][138] = 9'b111111111;
assign micromatrizz[91][139] = 9'b111111111;
assign micromatrizz[91][140] = 9'b111111111;
assign micromatrizz[91][141] = 9'b111111111;
assign micromatrizz[91][142] = 9'b111111111;
assign micromatrizz[91][143] = 9'b111111111;
assign micromatrizz[91][144] = 9'b111111111;
assign micromatrizz[91][145] = 9'b111111111;
assign micromatrizz[91][146] = 9'b111111111;
assign micromatrizz[91][147] = 9'b111111111;
assign micromatrizz[91][148] = 9'b111111111;
assign micromatrizz[91][149] = 9'b111111111;
assign micromatrizz[91][150] = 9'b111111111;
assign micromatrizz[91][151] = 9'b111111111;
assign micromatrizz[91][152] = 9'b111111111;
assign micromatrizz[91][153] = 9'b111111111;
assign micromatrizz[91][154] = 9'b111111111;
assign micromatrizz[91][155] = 9'b111111111;
assign micromatrizz[91][156] = 9'b111111111;
assign micromatrizz[91][157] = 9'b111111111;
assign micromatrizz[91][158] = 9'b111111111;
assign micromatrizz[91][159] = 9'b111111111;
assign micromatrizz[91][160] = 9'b111111111;
assign micromatrizz[91][161] = 9'b111111111;
assign micromatrizz[91][162] = 9'b111111111;
assign micromatrizz[91][163] = 9'b111111111;
assign micromatrizz[91][164] = 9'b111111111;
assign micromatrizz[91][165] = 9'b111111111;
assign micromatrizz[91][166] = 9'b111111111;
assign micromatrizz[91][167] = 9'b111111111;
assign micromatrizz[91][168] = 9'b111111111;
assign micromatrizz[91][169] = 9'b111111111;
assign micromatrizz[91][170] = 9'b111111111;
assign micromatrizz[91][171] = 9'b111111111;
assign micromatrizz[91][172] = 9'b111111111;
assign micromatrizz[91][173] = 9'b111111111;
assign micromatrizz[91][174] = 9'b111111111;
assign micromatrizz[91][175] = 9'b111111111;
assign micromatrizz[91][176] = 9'b111111111;
assign micromatrizz[91][177] = 9'b111111111;
assign micromatrizz[91][178] = 9'b111111111;
assign micromatrizz[91][179] = 9'b111111111;
assign micromatrizz[91][180] = 9'b111111111;
assign micromatrizz[91][181] = 9'b111111111;
assign micromatrizz[91][182] = 9'b111111111;
assign micromatrizz[91][183] = 9'b111111111;
assign micromatrizz[91][184] = 9'b111111111;
assign micromatrizz[91][185] = 9'b111111111;
assign micromatrizz[91][186] = 9'b111111111;
assign micromatrizz[91][187] = 9'b111111111;
assign micromatrizz[91][188] = 9'b111111111;
assign micromatrizz[91][189] = 9'b111111111;
assign micromatrizz[91][190] = 9'b111111111;
assign micromatrizz[91][191] = 9'b111111111;
assign micromatrizz[91][192] = 9'b111111111;
assign micromatrizz[91][193] = 9'b111111111;
assign micromatrizz[91][194] = 9'b111111111;
assign micromatrizz[91][195] = 9'b111111111;
assign micromatrizz[91][196] = 9'b111111111;
assign micromatrizz[91][197] = 9'b111111111;
assign micromatrizz[91][198] = 9'b111111111;
assign micromatrizz[91][199] = 9'b111111111;
assign micromatrizz[91][200] = 9'b111111111;
assign micromatrizz[91][201] = 9'b111111111;
assign micromatrizz[91][202] = 9'b111111111;
assign micromatrizz[91][203] = 9'b111111111;
assign micromatrizz[91][204] = 9'b111111111;
assign micromatrizz[91][205] = 9'b111111111;
assign micromatrizz[91][206] = 9'b111111111;
assign micromatrizz[91][207] = 9'b111111111;
assign micromatrizz[91][208] = 9'b111111111;
assign micromatrizz[91][209] = 9'b111111111;
assign micromatrizz[91][210] = 9'b111111111;
assign micromatrizz[91][211] = 9'b111111111;
assign micromatrizz[91][212] = 9'b111111111;
assign micromatrizz[91][213] = 9'b111111111;
assign micromatrizz[91][214] = 9'b111111111;
assign micromatrizz[91][215] = 9'b111111111;
assign micromatrizz[91][216] = 9'b111111111;
assign micromatrizz[91][217] = 9'b111111111;
assign micromatrizz[91][218] = 9'b111111111;
assign micromatrizz[91][219] = 9'b111111111;
assign micromatrizz[91][220] = 9'b111111111;
assign micromatrizz[91][221] = 9'b111111111;
assign micromatrizz[91][222] = 9'b111111111;
assign micromatrizz[91][223] = 9'b111111111;
assign micromatrizz[91][224] = 9'b111111111;
assign micromatrizz[91][225] = 9'b111111111;
assign micromatrizz[91][226] = 9'b111111111;
assign micromatrizz[91][227] = 9'b111111111;
assign micromatrizz[91][228] = 9'b111111111;
assign micromatrizz[91][229] = 9'b111111111;
assign micromatrizz[91][230] = 9'b111111111;
assign micromatrizz[91][231] = 9'b111111111;
assign micromatrizz[91][232] = 9'b111111111;
assign micromatrizz[91][233] = 9'b111111111;
assign micromatrizz[91][234] = 9'b111111111;
assign micromatrizz[91][235] = 9'b111111111;
assign micromatrizz[91][236] = 9'b111111111;
assign micromatrizz[91][237] = 9'b111111111;
assign micromatrizz[91][238] = 9'b111111111;
assign micromatrizz[91][239] = 9'b111111111;
assign micromatrizz[91][240] = 9'b111111111;
assign micromatrizz[91][241] = 9'b111111111;
assign micromatrizz[91][242] = 9'b111111111;
assign micromatrizz[91][243] = 9'b111111111;
assign micromatrizz[91][244] = 9'b111111111;
assign micromatrizz[91][245] = 9'b111111111;
assign micromatrizz[91][246] = 9'b111111111;
assign micromatrizz[91][247] = 9'b111111111;
assign micromatrizz[91][248] = 9'b111111111;
assign micromatrizz[91][249] = 9'b111111111;
assign micromatrizz[91][250] = 9'b111111111;
assign micromatrizz[91][251] = 9'b111111111;
assign micromatrizz[91][252] = 9'b111111111;
assign micromatrizz[91][253] = 9'b111111111;
assign micromatrizz[91][254] = 9'b111111111;
assign micromatrizz[91][255] = 9'b111111111;
assign micromatrizz[91][256] = 9'b111111111;
assign micromatrizz[91][257] = 9'b111111111;
assign micromatrizz[91][258] = 9'b111111111;
assign micromatrizz[91][259] = 9'b111111111;
assign micromatrizz[91][260] = 9'b111111111;
assign micromatrizz[91][261] = 9'b111111111;
assign micromatrizz[91][262] = 9'b111111111;
assign micromatrizz[91][263] = 9'b111111111;
assign micromatrizz[91][264] = 9'b111111111;
assign micromatrizz[91][265] = 9'b111111111;
assign micromatrizz[91][266] = 9'b111111111;
assign micromatrizz[91][267] = 9'b111111111;
assign micromatrizz[91][268] = 9'b111111111;
assign micromatrizz[91][269] = 9'b111111111;
assign micromatrizz[91][270] = 9'b111111111;
assign micromatrizz[91][271] = 9'b111111111;
assign micromatrizz[91][272] = 9'b111111111;
assign micromatrizz[91][273] = 9'b111111111;
assign micromatrizz[91][274] = 9'b111111111;
assign micromatrizz[91][275] = 9'b111111111;
assign micromatrizz[91][276] = 9'b111111111;
assign micromatrizz[91][277] = 9'b111111111;
assign micromatrizz[91][278] = 9'b111111111;
assign micromatrizz[91][279] = 9'b111111111;
assign micromatrizz[91][280] = 9'b111111111;
assign micromatrizz[91][281] = 9'b111111111;
assign micromatrizz[91][282] = 9'b111111111;
assign micromatrizz[91][283] = 9'b111111111;
assign micromatrizz[91][284] = 9'b111111111;
assign micromatrizz[91][285] = 9'b111111111;
assign micromatrizz[91][286] = 9'b111111111;
assign micromatrizz[91][287] = 9'b111111111;
assign micromatrizz[91][288] = 9'b111111111;
assign micromatrizz[91][289] = 9'b111111111;
assign micromatrizz[91][290] = 9'b111111111;
assign micromatrizz[91][291] = 9'b111111111;
assign micromatrizz[91][292] = 9'b111111111;
assign micromatrizz[91][293] = 9'b111111111;
assign micromatrizz[91][294] = 9'b111111111;
assign micromatrizz[91][295] = 9'b111111111;
assign micromatrizz[91][296] = 9'b111111111;
assign micromatrizz[91][297] = 9'b111111111;
assign micromatrizz[91][298] = 9'b111111111;
assign micromatrizz[91][299] = 9'b111111111;
assign micromatrizz[91][300] = 9'b111111111;
assign micromatrizz[91][301] = 9'b111111111;
assign micromatrizz[91][302] = 9'b111111111;
assign micromatrizz[91][303] = 9'b111111111;
assign micromatrizz[91][304] = 9'b111111111;
assign micromatrizz[91][305] = 9'b111111111;
assign micromatrizz[91][306] = 9'b111111111;
assign micromatrizz[91][307] = 9'b111111111;
assign micromatrizz[91][308] = 9'b111111111;
assign micromatrizz[91][309] = 9'b111111111;
assign micromatrizz[91][310] = 9'b111111111;
assign micromatrizz[91][311] = 9'b111111111;
assign micromatrizz[91][312] = 9'b111111111;
assign micromatrizz[91][313] = 9'b111111111;
assign micromatrizz[91][314] = 9'b111111111;
assign micromatrizz[91][315] = 9'b111111111;
assign micromatrizz[91][316] = 9'b111111111;
assign micromatrizz[91][317] = 9'b111111111;
assign micromatrizz[91][318] = 9'b111111111;
assign micromatrizz[91][319] = 9'b111111111;
assign micromatrizz[91][320] = 9'b111111111;
assign micromatrizz[91][321] = 9'b111111111;
assign micromatrizz[91][322] = 9'b111111111;
assign micromatrizz[91][323] = 9'b111111111;
assign micromatrizz[91][324] = 9'b111111111;
assign micromatrizz[91][325] = 9'b111111111;
assign micromatrizz[91][326] = 9'b111111111;
assign micromatrizz[91][327] = 9'b111111111;
assign micromatrizz[91][328] = 9'b111111111;
assign micromatrizz[91][329] = 9'b111111111;
assign micromatrizz[91][330] = 9'b111111111;
assign micromatrizz[91][331] = 9'b111111111;
assign micromatrizz[91][332] = 9'b111111111;
assign micromatrizz[91][333] = 9'b111111111;
assign micromatrizz[91][334] = 9'b111111111;
assign micromatrizz[91][335] = 9'b111111111;
assign micromatrizz[91][336] = 9'b111111111;
assign micromatrizz[91][337] = 9'b111111111;
assign micromatrizz[91][338] = 9'b111111111;
assign micromatrizz[91][339] = 9'b111111111;
assign micromatrizz[91][340] = 9'b111111111;
assign micromatrizz[91][341] = 9'b111111111;
assign micromatrizz[91][342] = 9'b111111111;
assign micromatrizz[91][343] = 9'b111111111;
assign micromatrizz[91][344] = 9'b111111111;
assign micromatrizz[91][345] = 9'b111111111;
assign micromatrizz[91][346] = 9'b111111111;
assign micromatrizz[91][347] = 9'b111111111;
assign micromatrizz[91][348] = 9'b111111111;
assign micromatrizz[91][349] = 9'b111111111;
assign micromatrizz[91][350] = 9'b111111111;
assign micromatrizz[91][351] = 9'b111111111;
assign micromatrizz[91][352] = 9'b111111111;
assign micromatrizz[91][353] = 9'b111111111;
assign micromatrizz[91][354] = 9'b111111111;
assign micromatrizz[91][355] = 9'b111111111;
assign micromatrizz[91][356] = 9'b111111111;
assign micromatrizz[91][357] = 9'b111111111;
assign micromatrizz[91][358] = 9'b111111111;
assign micromatrizz[91][359] = 9'b111111111;
assign micromatrizz[91][360] = 9'b111111111;
assign micromatrizz[91][361] = 9'b111111111;
assign micromatrizz[91][362] = 9'b111111111;
assign micromatrizz[91][363] = 9'b111111111;
assign micromatrizz[91][364] = 9'b111111111;
assign micromatrizz[91][365] = 9'b111111111;
assign micromatrizz[91][366] = 9'b111111111;
assign micromatrizz[91][367] = 9'b111111111;
assign micromatrizz[91][368] = 9'b111111111;
assign micromatrizz[91][369] = 9'b111111111;
assign micromatrizz[91][370] = 9'b111111111;
assign micromatrizz[91][371] = 9'b111111111;
assign micromatrizz[91][372] = 9'b111111111;
assign micromatrizz[91][373] = 9'b111111111;
assign micromatrizz[91][374] = 9'b111111111;
assign micromatrizz[91][375] = 9'b111111111;
assign micromatrizz[91][376] = 9'b111111111;
assign micromatrizz[91][377] = 9'b111111111;
assign micromatrizz[91][378] = 9'b111111111;
assign micromatrizz[91][379] = 9'b111111111;
assign micromatrizz[91][380] = 9'b111111111;
assign micromatrizz[91][381] = 9'b111111111;
assign micromatrizz[91][382] = 9'b111111111;
assign micromatrizz[91][383] = 9'b111111111;
assign micromatrizz[91][384] = 9'b111111111;
assign micromatrizz[91][385] = 9'b111111111;
assign micromatrizz[91][386] = 9'b111111111;
assign micromatrizz[91][387] = 9'b111111111;
assign micromatrizz[91][388] = 9'b111111111;
assign micromatrizz[91][389] = 9'b111111111;
assign micromatrizz[91][390] = 9'b111111111;
assign micromatrizz[91][391] = 9'b111111111;
assign micromatrizz[91][392] = 9'b111111111;
assign micromatrizz[91][393] = 9'b111111111;
assign micromatrizz[91][394] = 9'b111111111;
assign micromatrizz[91][395] = 9'b111111111;
assign micromatrizz[91][396] = 9'b111111111;
assign micromatrizz[91][397] = 9'b111111111;
assign micromatrizz[91][398] = 9'b111111111;
assign micromatrizz[91][399] = 9'b111111111;
assign micromatrizz[91][400] = 9'b111111111;
assign micromatrizz[91][401] = 9'b111111111;
assign micromatrizz[91][402] = 9'b111111111;
assign micromatrizz[91][403] = 9'b111111111;
assign micromatrizz[91][404] = 9'b111111111;
assign micromatrizz[91][405] = 9'b111111111;
assign micromatrizz[91][406] = 9'b111111111;
assign micromatrizz[91][407] = 9'b111111111;
assign micromatrizz[91][408] = 9'b111111111;
assign micromatrizz[91][409] = 9'b111111111;
assign micromatrizz[91][410] = 9'b111111111;
assign micromatrizz[91][411] = 9'b111111111;
assign micromatrizz[91][412] = 9'b111111111;
assign micromatrizz[91][413] = 9'b111111111;
assign micromatrizz[91][414] = 9'b111111111;
assign micromatrizz[91][415] = 9'b111111111;
assign micromatrizz[91][416] = 9'b111111111;
assign micromatrizz[91][417] = 9'b111111111;
assign micromatrizz[91][418] = 9'b111111111;
assign micromatrizz[91][419] = 9'b111111111;
assign micromatrizz[91][420] = 9'b111111111;
assign micromatrizz[91][421] = 9'b111111111;
assign micromatrizz[91][422] = 9'b111111111;
assign micromatrizz[91][423] = 9'b111111111;
assign micromatrizz[91][424] = 9'b111111111;
assign micromatrizz[91][425] = 9'b111111111;
assign micromatrizz[91][426] = 9'b111111111;
assign micromatrizz[91][427] = 9'b111111111;
assign micromatrizz[91][428] = 9'b111111111;
assign micromatrizz[91][429] = 9'b111111111;
assign micromatrizz[91][430] = 9'b111111111;
assign micromatrizz[91][431] = 9'b111111111;
assign micromatrizz[91][432] = 9'b111111111;
assign micromatrizz[91][433] = 9'b111111111;
assign micromatrizz[91][434] = 9'b111111111;
assign micromatrizz[91][435] = 9'b111111111;
assign micromatrizz[91][436] = 9'b111111111;
assign micromatrizz[91][437] = 9'b111111111;
assign micromatrizz[91][438] = 9'b111111111;
assign micromatrizz[91][439] = 9'b111111111;
assign micromatrizz[91][440] = 9'b111111111;
assign micromatrizz[91][441] = 9'b111111111;
assign micromatrizz[91][442] = 9'b111111111;
assign micromatrizz[91][443] = 9'b111111111;
assign micromatrizz[91][444] = 9'b111111111;
assign micromatrizz[91][445] = 9'b111111111;
assign micromatrizz[91][446] = 9'b111111111;
assign micromatrizz[91][447] = 9'b111111111;
assign micromatrizz[91][448] = 9'b111111111;
assign micromatrizz[91][449] = 9'b111111111;
assign micromatrizz[91][450] = 9'b111111111;
assign micromatrizz[91][451] = 9'b111111111;
assign micromatrizz[91][452] = 9'b111111111;
assign micromatrizz[91][453] = 9'b111111111;
assign micromatrizz[91][454] = 9'b111111111;
assign micromatrizz[91][455] = 9'b111111111;
assign micromatrizz[91][456] = 9'b111111111;
assign micromatrizz[91][457] = 9'b111111111;
assign micromatrizz[91][458] = 9'b111111111;
assign micromatrizz[91][459] = 9'b111111111;
assign micromatrizz[91][460] = 9'b111111111;
assign micromatrizz[91][461] = 9'b111111111;
assign micromatrizz[91][462] = 9'b111111111;
assign micromatrizz[91][463] = 9'b111111111;
assign micromatrizz[91][464] = 9'b111111111;
assign micromatrizz[91][465] = 9'b111111111;
assign micromatrizz[91][466] = 9'b111111111;
assign micromatrizz[91][467] = 9'b111111111;
assign micromatrizz[91][468] = 9'b111111111;
assign micromatrizz[91][469] = 9'b111111111;
assign micromatrizz[91][470] = 9'b111111111;
assign micromatrizz[91][471] = 9'b111111111;
assign micromatrizz[91][472] = 9'b111111111;
assign micromatrizz[91][473] = 9'b111111111;
assign micromatrizz[91][474] = 9'b111111111;
assign micromatrizz[91][475] = 9'b111111111;
assign micromatrizz[91][476] = 9'b111111111;
assign micromatrizz[91][477] = 9'b111111111;
assign micromatrizz[91][478] = 9'b111111111;
assign micromatrizz[91][479] = 9'b111111111;
assign micromatrizz[91][480] = 9'b111111111;
assign micromatrizz[91][481] = 9'b111111111;
assign micromatrizz[91][482] = 9'b111111111;
assign micromatrizz[91][483] = 9'b111111111;
assign micromatrizz[91][484] = 9'b111111111;
assign micromatrizz[91][485] = 9'b111111111;
assign micromatrizz[91][486] = 9'b111111111;
assign micromatrizz[91][487] = 9'b111111111;
assign micromatrizz[91][488] = 9'b111111111;
assign micromatrizz[91][489] = 9'b111111111;
assign micromatrizz[91][490] = 9'b111111111;
assign micromatrizz[91][491] = 9'b111111111;
assign micromatrizz[91][492] = 9'b111111111;
assign micromatrizz[91][493] = 9'b111111111;
assign micromatrizz[91][494] = 9'b111111111;
assign micromatrizz[91][495] = 9'b111111111;
assign micromatrizz[91][496] = 9'b111111111;
assign micromatrizz[91][497] = 9'b111111111;
assign micromatrizz[91][498] = 9'b111111111;
assign micromatrizz[91][499] = 9'b111111111;
assign micromatrizz[91][500] = 9'b111111111;
assign micromatrizz[91][501] = 9'b111111111;
assign micromatrizz[91][502] = 9'b111111111;
assign micromatrizz[91][503] = 9'b111111111;
assign micromatrizz[91][504] = 9'b111111111;
assign micromatrizz[91][505] = 9'b111111111;
assign micromatrizz[91][506] = 9'b111111111;
assign micromatrizz[91][507] = 9'b111111111;
assign micromatrizz[91][508] = 9'b111111111;
assign micromatrizz[91][509] = 9'b111111111;
assign micromatrizz[91][510] = 9'b111111111;
assign micromatrizz[91][511] = 9'b111111111;
assign micromatrizz[91][512] = 9'b111111111;
assign micromatrizz[91][513] = 9'b111111111;
assign micromatrizz[91][514] = 9'b111111111;
assign micromatrizz[91][515] = 9'b111111111;
assign micromatrizz[91][516] = 9'b111111111;
assign micromatrizz[91][517] = 9'b111111111;
assign micromatrizz[91][518] = 9'b111111111;
assign micromatrizz[91][519] = 9'b111111111;
assign micromatrizz[91][520] = 9'b111111111;
assign micromatrizz[91][521] = 9'b111111111;
assign micromatrizz[91][522] = 9'b111111111;
assign micromatrizz[91][523] = 9'b111111111;
assign micromatrizz[91][524] = 9'b111111111;
assign micromatrizz[91][525] = 9'b111111111;
assign micromatrizz[91][526] = 9'b111111111;
assign micromatrizz[91][527] = 9'b111111111;
assign micromatrizz[91][528] = 9'b111111111;
assign micromatrizz[91][529] = 9'b111111111;
assign micromatrizz[91][530] = 9'b111111111;
assign micromatrizz[91][531] = 9'b111111111;
assign micromatrizz[91][532] = 9'b111111111;
assign micromatrizz[91][533] = 9'b111111111;
assign micromatrizz[91][534] = 9'b111111111;
assign micromatrizz[91][535] = 9'b111111111;
assign micromatrizz[91][536] = 9'b111111111;
assign micromatrizz[91][537] = 9'b111111111;
assign micromatrizz[91][538] = 9'b111111111;
assign micromatrizz[91][539] = 9'b111111111;
assign micromatrizz[91][540] = 9'b111111111;
assign micromatrizz[91][541] = 9'b111111111;
assign micromatrizz[91][542] = 9'b111111111;
assign micromatrizz[91][543] = 9'b111111111;
assign micromatrizz[91][544] = 9'b111111111;
assign micromatrizz[91][545] = 9'b111111111;
assign micromatrizz[91][546] = 9'b111111111;
assign micromatrizz[91][547] = 9'b111111111;
assign micromatrizz[91][548] = 9'b111111111;
assign micromatrizz[91][549] = 9'b111111111;
assign micromatrizz[91][550] = 9'b111111111;
assign micromatrizz[91][551] = 9'b111111111;
assign micromatrizz[91][552] = 9'b111111111;
assign micromatrizz[91][553] = 9'b111111111;
assign micromatrizz[91][554] = 9'b111111111;
assign micromatrizz[91][555] = 9'b111111111;
assign micromatrizz[91][556] = 9'b111111111;
assign micromatrizz[91][557] = 9'b111111111;
assign micromatrizz[91][558] = 9'b111111111;
assign micromatrizz[91][559] = 9'b111111111;
assign micromatrizz[91][560] = 9'b111111111;
assign micromatrizz[91][561] = 9'b111111111;
assign micromatrizz[91][562] = 9'b111111111;
assign micromatrizz[91][563] = 9'b111111111;
assign micromatrizz[91][564] = 9'b111111111;
assign micromatrizz[91][565] = 9'b111111111;
assign micromatrizz[91][566] = 9'b111111111;
assign micromatrizz[91][567] = 9'b111111111;
assign micromatrizz[91][568] = 9'b111111111;
assign micromatrizz[91][569] = 9'b111111111;
assign micromatrizz[91][570] = 9'b111111111;
assign micromatrizz[91][571] = 9'b111111111;
assign micromatrizz[91][572] = 9'b111111111;
assign micromatrizz[91][573] = 9'b111111111;
assign micromatrizz[91][574] = 9'b111111111;
assign micromatrizz[91][575] = 9'b111111111;
assign micromatrizz[91][576] = 9'b111111111;
assign micromatrizz[91][577] = 9'b111111111;
assign micromatrizz[91][578] = 9'b111111111;
assign micromatrizz[91][579] = 9'b111111111;
assign micromatrizz[91][580] = 9'b111111111;
assign micromatrizz[91][581] = 9'b111111111;
assign micromatrizz[91][582] = 9'b111111111;
assign micromatrizz[91][583] = 9'b111111111;
assign micromatrizz[91][584] = 9'b111111111;
assign micromatrizz[91][585] = 9'b111111111;
assign micromatrizz[91][586] = 9'b111111111;
assign micromatrizz[91][587] = 9'b111111111;
assign micromatrizz[91][588] = 9'b111111111;
assign micromatrizz[91][589] = 9'b111111111;
assign micromatrizz[91][590] = 9'b111111111;
assign micromatrizz[91][591] = 9'b111111111;
assign micromatrizz[91][592] = 9'b111111111;
assign micromatrizz[91][593] = 9'b111111111;
assign micromatrizz[91][594] = 9'b111111111;
assign micromatrizz[91][595] = 9'b111111111;
assign micromatrizz[91][596] = 9'b111111111;
assign micromatrizz[91][597] = 9'b111111111;
assign micromatrizz[91][598] = 9'b111111111;
assign micromatrizz[91][599] = 9'b111111111;
assign micromatrizz[91][600] = 9'b111111111;
assign micromatrizz[91][601] = 9'b111111111;
assign micromatrizz[91][602] = 9'b111111111;
assign micromatrizz[91][603] = 9'b111111111;
assign micromatrizz[91][604] = 9'b111111111;
assign micromatrizz[91][605] = 9'b111111111;
assign micromatrizz[91][606] = 9'b111111111;
assign micromatrizz[91][607] = 9'b111111111;
assign micromatrizz[91][608] = 9'b111111111;
assign micromatrizz[91][609] = 9'b111111111;
assign micromatrizz[91][610] = 9'b111111111;
assign micromatrizz[91][611] = 9'b111111111;
assign micromatrizz[91][612] = 9'b111111111;
assign micromatrizz[91][613] = 9'b111111111;
assign micromatrizz[91][614] = 9'b111111111;
assign micromatrizz[91][615] = 9'b111111111;
assign micromatrizz[91][616] = 9'b111111111;
assign micromatrizz[91][617] = 9'b111111111;
assign micromatrizz[91][618] = 9'b111111111;
assign micromatrizz[91][619] = 9'b111111111;
assign micromatrizz[91][620] = 9'b111111111;
assign micromatrizz[91][621] = 9'b111111111;
assign micromatrizz[91][622] = 9'b111111111;
assign micromatrizz[91][623] = 9'b111111111;
assign micromatrizz[91][624] = 9'b111111111;
assign micromatrizz[91][625] = 9'b111111111;
assign micromatrizz[91][626] = 9'b111111111;
assign micromatrizz[91][627] = 9'b111111111;
assign micromatrizz[91][628] = 9'b111111111;
assign micromatrizz[91][629] = 9'b111111111;
assign micromatrizz[91][630] = 9'b111111111;
assign micromatrizz[91][631] = 9'b111111111;
assign micromatrizz[91][632] = 9'b111111111;
assign micromatrizz[91][633] = 9'b111111111;
assign micromatrizz[91][634] = 9'b111111111;
assign micromatrizz[91][635] = 9'b111111111;
assign micromatrizz[91][636] = 9'b111111111;
assign micromatrizz[91][637] = 9'b111111111;
assign micromatrizz[91][638] = 9'b111111111;
assign micromatrizz[91][639] = 9'b111111111;
assign micromatrizz[92][0] = 9'b111111111;
assign micromatrizz[92][1] = 9'b111111111;
assign micromatrizz[92][2] = 9'b111111111;
assign micromatrizz[92][3] = 9'b111111111;
assign micromatrizz[92][4] = 9'b111111111;
assign micromatrizz[92][5] = 9'b111111111;
assign micromatrizz[92][6] = 9'b111111111;
assign micromatrizz[92][7] = 9'b111111111;
assign micromatrizz[92][8] = 9'b111111111;
assign micromatrizz[92][9] = 9'b111111111;
assign micromatrizz[92][10] = 9'b111111111;
assign micromatrizz[92][11] = 9'b111111111;
assign micromatrizz[92][12] = 9'b111111111;
assign micromatrizz[92][13] = 9'b111111111;
assign micromatrizz[92][14] = 9'b111111111;
assign micromatrizz[92][15] = 9'b111111111;
assign micromatrizz[92][16] = 9'b111111111;
assign micromatrizz[92][17] = 9'b111111111;
assign micromatrizz[92][18] = 9'b111111111;
assign micromatrizz[92][19] = 9'b111111111;
assign micromatrizz[92][20] = 9'b111111111;
assign micromatrizz[92][21] = 9'b111111111;
assign micromatrizz[92][22] = 9'b111111111;
assign micromatrizz[92][23] = 9'b111111111;
assign micromatrizz[92][24] = 9'b111111111;
assign micromatrizz[92][25] = 9'b111111111;
assign micromatrizz[92][26] = 9'b111111111;
assign micromatrizz[92][27] = 9'b111111111;
assign micromatrizz[92][28] = 9'b111111111;
assign micromatrizz[92][29] = 9'b111111111;
assign micromatrizz[92][30] = 9'b111111111;
assign micromatrizz[92][31] = 9'b111111111;
assign micromatrizz[92][32] = 9'b111111111;
assign micromatrizz[92][33] = 9'b111111111;
assign micromatrizz[92][34] = 9'b111111111;
assign micromatrizz[92][35] = 9'b111111111;
assign micromatrizz[92][36] = 9'b111111111;
assign micromatrizz[92][37] = 9'b111111111;
assign micromatrizz[92][38] = 9'b111111111;
assign micromatrizz[92][39] = 9'b111111111;
assign micromatrizz[92][40] = 9'b111111111;
assign micromatrizz[92][41] = 9'b111111111;
assign micromatrizz[92][42] = 9'b111111111;
assign micromatrizz[92][43] = 9'b111111111;
assign micromatrizz[92][44] = 9'b111111111;
assign micromatrizz[92][45] = 9'b111111111;
assign micromatrizz[92][46] = 9'b111111111;
assign micromatrizz[92][47] = 9'b111111111;
assign micromatrizz[92][48] = 9'b111111111;
assign micromatrizz[92][49] = 9'b111111111;
assign micromatrizz[92][50] = 9'b111111111;
assign micromatrizz[92][51] = 9'b111111111;
assign micromatrizz[92][52] = 9'b111111111;
assign micromatrizz[92][53] = 9'b111111111;
assign micromatrizz[92][54] = 9'b111111111;
assign micromatrizz[92][55] = 9'b111111111;
assign micromatrizz[92][56] = 9'b111111111;
assign micromatrizz[92][57] = 9'b111111111;
assign micromatrizz[92][58] = 9'b111111111;
assign micromatrizz[92][59] = 9'b111111111;
assign micromatrizz[92][60] = 9'b111111111;
assign micromatrizz[92][61] = 9'b111111111;
assign micromatrizz[92][62] = 9'b111111111;
assign micromatrizz[92][63] = 9'b111111111;
assign micromatrizz[92][64] = 9'b111111111;
assign micromatrizz[92][65] = 9'b111111111;
assign micromatrizz[92][66] = 9'b111111111;
assign micromatrizz[92][67] = 9'b111111111;
assign micromatrizz[92][68] = 9'b111111111;
assign micromatrizz[92][69] = 9'b111111111;
assign micromatrizz[92][70] = 9'b111111111;
assign micromatrizz[92][71] = 9'b111111111;
assign micromatrizz[92][72] = 9'b111111111;
assign micromatrizz[92][73] = 9'b111111111;
assign micromatrizz[92][74] = 9'b111111111;
assign micromatrizz[92][75] = 9'b111111111;
assign micromatrizz[92][76] = 9'b111111111;
assign micromatrizz[92][77] = 9'b111111111;
assign micromatrizz[92][78] = 9'b111111111;
assign micromatrizz[92][79] = 9'b111111111;
assign micromatrizz[92][80] = 9'b111111111;
assign micromatrizz[92][81] = 9'b111111111;
assign micromatrizz[92][82] = 9'b111111111;
assign micromatrizz[92][83] = 9'b111111111;
assign micromatrizz[92][84] = 9'b111111111;
assign micromatrizz[92][85] = 9'b111111111;
assign micromatrizz[92][86] = 9'b111111111;
assign micromatrizz[92][87] = 9'b111111111;
assign micromatrizz[92][88] = 9'b111111111;
assign micromatrizz[92][89] = 9'b111111111;
assign micromatrizz[92][90] = 9'b111111111;
assign micromatrizz[92][91] = 9'b111111111;
assign micromatrizz[92][92] = 9'b111111111;
assign micromatrizz[92][93] = 9'b111111111;
assign micromatrizz[92][94] = 9'b111111111;
assign micromatrizz[92][95] = 9'b111111111;
assign micromatrizz[92][96] = 9'b111111111;
assign micromatrizz[92][97] = 9'b111111111;
assign micromatrizz[92][98] = 9'b111111111;
assign micromatrizz[92][99] = 9'b111111111;
assign micromatrizz[92][100] = 9'b111111111;
assign micromatrizz[92][101] = 9'b111111111;
assign micromatrizz[92][102] = 9'b111111111;
assign micromatrizz[92][103] = 9'b111111111;
assign micromatrizz[92][104] = 9'b111111111;
assign micromatrizz[92][105] = 9'b111111111;
assign micromatrizz[92][106] = 9'b111111111;
assign micromatrizz[92][107] = 9'b111111111;
assign micromatrizz[92][108] = 9'b111111111;
assign micromatrizz[92][109] = 9'b111111111;
assign micromatrizz[92][110] = 9'b111111111;
assign micromatrizz[92][111] = 9'b111111111;
assign micromatrizz[92][112] = 9'b111111111;
assign micromatrizz[92][113] = 9'b111111111;
assign micromatrizz[92][114] = 9'b111111111;
assign micromatrizz[92][115] = 9'b111111111;
assign micromatrizz[92][116] = 9'b111111111;
assign micromatrizz[92][117] = 9'b111111111;
assign micromatrizz[92][118] = 9'b111111111;
assign micromatrizz[92][119] = 9'b111111111;
assign micromatrizz[92][120] = 9'b111111111;
assign micromatrizz[92][121] = 9'b111111111;
assign micromatrizz[92][122] = 9'b111111111;
assign micromatrizz[92][123] = 9'b111111111;
assign micromatrizz[92][124] = 9'b111111111;
assign micromatrizz[92][125] = 9'b111111111;
assign micromatrizz[92][126] = 9'b111111111;
assign micromatrizz[92][127] = 9'b111111111;
assign micromatrizz[92][128] = 9'b111111111;
assign micromatrizz[92][129] = 9'b111111111;
assign micromatrizz[92][130] = 9'b111111111;
assign micromatrizz[92][131] = 9'b111111111;
assign micromatrizz[92][132] = 9'b111111111;
assign micromatrizz[92][133] = 9'b111111111;
assign micromatrizz[92][134] = 9'b111111111;
assign micromatrizz[92][135] = 9'b111111111;
assign micromatrizz[92][136] = 9'b111111111;
assign micromatrizz[92][137] = 9'b111111111;
assign micromatrizz[92][138] = 9'b111111111;
assign micromatrizz[92][139] = 9'b111111111;
assign micromatrizz[92][140] = 9'b111111111;
assign micromatrizz[92][141] = 9'b111111111;
assign micromatrizz[92][142] = 9'b111111111;
assign micromatrizz[92][143] = 9'b111111111;
assign micromatrizz[92][144] = 9'b111111111;
assign micromatrizz[92][145] = 9'b111111111;
assign micromatrizz[92][146] = 9'b111111111;
assign micromatrizz[92][147] = 9'b111111111;
assign micromatrizz[92][148] = 9'b111111111;
assign micromatrizz[92][149] = 9'b111111111;
assign micromatrizz[92][150] = 9'b111111111;
assign micromatrizz[92][151] = 9'b111111111;
assign micromatrizz[92][152] = 9'b111111111;
assign micromatrizz[92][153] = 9'b111111111;
assign micromatrizz[92][154] = 9'b111111111;
assign micromatrizz[92][155] = 9'b111111111;
assign micromatrizz[92][156] = 9'b111111111;
assign micromatrizz[92][157] = 9'b111111111;
assign micromatrizz[92][158] = 9'b111111111;
assign micromatrizz[92][159] = 9'b111111111;
assign micromatrizz[92][160] = 9'b111111111;
assign micromatrizz[92][161] = 9'b111111111;
assign micromatrizz[92][162] = 9'b111111111;
assign micromatrizz[92][163] = 9'b111111111;
assign micromatrizz[92][164] = 9'b111111111;
assign micromatrizz[92][165] = 9'b111111111;
assign micromatrizz[92][166] = 9'b111111111;
assign micromatrizz[92][167] = 9'b111111111;
assign micromatrizz[92][168] = 9'b111111111;
assign micromatrizz[92][169] = 9'b111111111;
assign micromatrizz[92][170] = 9'b111111111;
assign micromatrizz[92][171] = 9'b111111111;
assign micromatrizz[92][172] = 9'b111111111;
assign micromatrizz[92][173] = 9'b111111111;
assign micromatrizz[92][174] = 9'b111111111;
assign micromatrizz[92][175] = 9'b111111111;
assign micromatrizz[92][176] = 9'b111111111;
assign micromatrizz[92][177] = 9'b111111111;
assign micromatrizz[92][178] = 9'b111111111;
assign micromatrizz[92][179] = 9'b111111111;
assign micromatrizz[92][180] = 9'b111111111;
assign micromatrizz[92][181] = 9'b111111111;
assign micromatrizz[92][182] = 9'b111111111;
assign micromatrizz[92][183] = 9'b111111111;
assign micromatrizz[92][184] = 9'b111111111;
assign micromatrizz[92][185] = 9'b111111111;
assign micromatrizz[92][186] = 9'b111111111;
assign micromatrizz[92][187] = 9'b111111111;
assign micromatrizz[92][188] = 9'b111111111;
assign micromatrizz[92][189] = 9'b111111111;
assign micromatrizz[92][190] = 9'b111111111;
assign micromatrizz[92][191] = 9'b111111111;
assign micromatrizz[92][192] = 9'b111111111;
assign micromatrizz[92][193] = 9'b111111111;
assign micromatrizz[92][194] = 9'b111111111;
assign micromatrizz[92][195] = 9'b111111111;
assign micromatrizz[92][196] = 9'b111111111;
assign micromatrizz[92][197] = 9'b111111111;
assign micromatrizz[92][198] = 9'b111111111;
assign micromatrizz[92][199] = 9'b111111111;
assign micromatrizz[92][200] = 9'b111111111;
assign micromatrizz[92][201] = 9'b111111111;
assign micromatrizz[92][202] = 9'b111111111;
assign micromatrizz[92][203] = 9'b111111111;
assign micromatrizz[92][204] = 9'b111111111;
assign micromatrizz[92][205] = 9'b111111111;
assign micromatrizz[92][206] = 9'b111111111;
assign micromatrizz[92][207] = 9'b111111111;
assign micromatrizz[92][208] = 9'b111111111;
assign micromatrizz[92][209] = 9'b111111111;
assign micromatrizz[92][210] = 9'b111111111;
assign micromatrizz[92][211] = 9'b111111111;
assign micromatrizz[92][212] = 9'b111111111;
assign micromatrizz[92][213] = 9'b111111111;
assign micromatrizz[92][214] = 9'b111111111;
assign micromatrizz[92][215] = 9'b111111111;
assign micromatrizz[92][216] = 9'b111111111;
assign micromatrizz[92][217] = 9'b111111111;
assign micromatrizz[92][218] = 9'b111111111;
assign micromatrizz[92][219] = 9'b111111111;
assign micromatrizz[92][220] = 9'b111111111;
assign micromatrizz[92][221] = 9'b111111111;
assign micromatrizz[92][222] = 9'b111111111;
assign micromatrizz[92][223] = 9'b111111111;
assign micromatrizz[92][224] = 9'b111111111;
assign micromatrizz[92][225] = 9'b111111111;
assign micromatrizz[92][226] = 9'b111111111;
assign micromatrizz[92][227] = 9'b111111111;
assign micromatrizz[92][228] = 9'b111111111;
assign micromatrizz[92][229] = 9'b111111111;
assign micromatrizz[92][230] = 9'b111111111;
assign micromatrizz[92][231] = 9'b111111111;
assign micromatrizz[92][232] = 9'b111111111;
assign micromatrizz[92][233] = 9'b111111111;
assign micromatrizz[92][234] = 9'b111111111;
assign micromatrizz[92][235] = 9'b111111111;
assign micromatrizz[92][236] = 9'b111111111;
assign micromatrizz[92][237] = 9'b111111111;
assign micromatrizz[92][238] = 9'b111111111;
assign micromatrizz[92][239] = 9'b111111111;
assign micromatrizz[92][240] = 9'b111111111;
assign micromatrizz[92][241] = 9'b111111111;
assign micromatrizz[92][242] = 9'b111111111;
assign micromatrizz[92][243] = 9'b111111111;
assign micromatrizz[92][244] = 9'b111111111;
assign micromatrizz[92][245] = 9'b111111111;
assign micromatrizz[92][246] = 9'b111111111;
assign micromatrizz[92][247] = 9'b111111111;
assign micromatrizz[92][248] = 9'b111111111;
assign micromatrizz[92][249] = 9'b111111111;
assign micromatrizz[92][250] = 9'b111111111;
assign micromatrizz[92][251] = 9'b111111111;
assign micromatrizz[92][252] = 9'b111111111;
assign micromatrizz[92][253] = 9'b111111111;
assign micromatrizz[92][254] = 9'b111111111;
assign micromatrizz[92][255] = 9'b111111111;
assign micromatrizz[92][256] = 9'b111111111;
assign micromatrizz[92][257] = 9'b111111111;
assign micromatrizz[92][258] = 9'b111111111;
assign micromatrizz[92][259] = 9'b111111111;
assign micromatrizz[92][260] = 9'b111111111;
assign micromatrizz[92][261] = 9'b111111111;
assign micromatrizz[92][262] = 9'b111111111;
assign micromatrizz[92][263] = 9'b111111111;
assign micromatrizz[92][264] = 9'b111111111;
assign micromatrizz[92][265] = 9'b111111111;
assign micromatrizz[92][266] = 9'b111111111;
assign micromatrizz[92][267] = 9'b111111111;
assign micromatrizz[92][268] = 9'b111111111;
assign micromatrizz[92][269] = 9'b111111111;
assign micromatrizz[92][270] = 9'b111111111;
assign micromatrizz[92][271] = 9'b111111111;
assign micromatrizz[92][272] = 9'b111111111;
assign micromatrizz[92][273] = 9'b111111111;
assign micromatrizz[92][274] = 9'b111111111;
assign micromatrizz[92][275] = 9'b111111111;
assign micromatrizz[92][276] = 9'b111111111;
assign micromatrizz[92][277] = 9'b111111111;
assign micromatrizz[92][278] = 9'b111111111;
assign micromatrizz[92][279] = 9'b111111111;
assign micromatrizz[92][280] = 9'b111111111;
assign micromatrizz[92][281] = 9'b111111111;
assign micromatrizz[92][282] = 9'b111111111;
assign micromatrizz[92][283] = 9'b111111111;
assign micromatrizz[92][284] = 9'b111111111;
assign micromatrizz[92][285] = 9'b111111111;
assign micromatrizz[92][286] = 9'b111111111;
assign micromatrizz[92][287] = 9'b111111111;
assign micromatrizz[92][288] = 9'b111111111;
assign micromatrizz[92][289] = 9'b111111111;
assign micromatrizz[92][290] = 9'b111111111;
assign micromatrizz[92][291] = 9'b111111111;
assign micromatrizz[92][292] = 9'b111111111;
assign micromatrizz[92][293] = 9'b111111111;
assign micromatrizz[92][294] = 9'b111111111;
assign micromatrizz[92][295] = 9'b111111111;
assign micromatrizz[92][296] = 9'b111111111;
assign micromatrizz[92][297] = 9'b111111111;
assign micromatrizz[92][298] = 9'b111111111;
assign micromatrizz[92][299] = 9'b111111111;
assign micromatrizz[92][300] = 9'b111111111;
assign micromatrizz[92][301] = 9'b111111111;
assign micromatrizz[92][302] = 9'b111111111;
assign micromatrizz[92][303] = 9'b111111111;
assign micromatrizz[92][304] = 9'b111111111;
assign micromatrizz[92][305] = 9'b111111111;
assign micromatrizz[92][306] = 9'b111111111;
assign micromatrizz[92][307] = 9'b111111111;
assign micromatrizz[92][308] = 9'b111111111;
assign micromatrizz[92][309] = 9'b111111111;
assign micromatrizz[92][310] = 9'b111111111;
assign micromatrizz[92][311] = 9'b111111111;
assign micromatrizz[92][312] = 9'b111111111;
assign micromatrizz[92][313] = 9'b111111111;
assign micromatrizz[92][314] = 9'b111111111;
assign micromatrizz[92][315] = 9'b111111111;
assign micromatrizz[92][316] = 9'b111111111;
assign micromatrizz[92][317] = 9'b111111111;
assign micromatrizz[92][318] = 9'b111111111;
assign micromatrizz[92][319] = 9'b111111111;
assign micromatrizz[92][320] = 9'b111111111;
assign micromatrizz[92][321] = 9'b111111111;
assign micromatrizz[92][322] = 9'b111111111;
assign micromatrizz[92][323] = 9'b111111111;
assign micromatrizz[92][324] = 9'b111111111;
assign micromatrizz[92][325] = 9'b111111111;
assign micromatrizz[92][326] = 9'b111111111;
assign micromatrizz[92][327] = 9'b111111111;
assign micromatrizz[92][328] = 9'b111111111;
assign micromatrizz[92][329] = 9'b111111111;
assign micromatrizz[92][330] = 9'b111111111;
assign micromatrizz[92][331] = 9'b111111111;
assign micromatrizz[92][332] = 9'b111111111;
assign micromatrizz[92][333] = 9'b111111111;
assign micromatrizz[92][334] = 9'b111111111;
assign micromatrizz[92][335] = 9'b111111111;
assign micromatrizz[92][336] = 9'b111111111;
assign micromatrizz[92][337] = 9'b111111111;
assign micromatrizz[92][338] = 9'b111111111;
assign micromatrizz[92][339] = 9'b111111111;
assign micromatrizz[92][340] = 9'b111111111;
assign micromatrizz[92][341] = 9'b111111111;
assign micromatrizz[92][342] = 9'b111111111;
assign micromatrizz[92][343] = 9'b111111111;
assign micromatrizz[92][344] = 9'b111111111;
assign micromatrizz[92][345] = 9'b111111111;
assign micromatrizz[92][346] = 9'b111111111;
assign micromatrizz[92][347] = 9'b111111111;
assign micromatrizz[92][348] = 9'b111111111;
assign micromatrizz[92][349] = 9'b111111111;
assign micromatrizz[92][350] = 9'b111111111;
assign micromatrizz[92][351] = 9'b111111111;
assign micromatrizz[92][352] = 9'b111111111;
assign micromatrizz[92][353] = 9'b111111111;
assign micromatrizz[92][354] = 9'b111111111;
assign micromatrizz[92][355] = 9'b111111111;
assign micromatrizz[92][356] = 9'b111111111;
assign micromatrizz[92][357] = 9'b111111111;
assign micromatrizz[92][358] = 9'b111111111;
assign micromatrizz[92][359] = 9'b111111111;
assign micromatrizz[92][360] = 9'b111111111;
assign micromatrizz[92][361] = 9'b111111111;
assign micromatrizz[92][362] = 9'b111111111;
assign micromatrizz[92][363] = 9'b111111111;
assign micromatrizz[92][364] = 9'b111111111;
assign micromatrizz[92][365] = 9'b111111111;
assign micromatrizz[92][366] = 9'b111111111;
assign micromatrizz[92][367] = 9'b111111111;
assign micromatrizz[92][368] = 9'b111111111;
assign micromatrizz[92][369] = 9'b111111111;
assign micromatrizz[92][370] = 9'b111111111;
assign micromatrizz[92][371] = 9'b111111111;
assign micromatrizz[92][372] = 9'b111111111;
assign micromatrizz[92][373] = 9'b111111111;
assign micromatrizz[92][374] = 9'b111111111;
assign micromatrizz[92][375] = 9'b111111111;
assign micromatrizz[92][376] = 9'b111111111;
assign micromatrizz[92][377] = 9'b111111111;
assign micromatrizz[92][378] = 9'b111111111;
assign micromatrizz[92][379] = 9'b111111111;
assign micromatrizz[92][380] = 9'b111111111;
assign micromatrizz[92][381] = 9'b111111111;
assign micromatrizz[92][382] = 9'b111111111;
assign micromatrizz[92][383] = 9'b111111111;
assign micromatrizz[92][384] = 9'b111111111;
assign micromatrizz[92][385] = 9'b111111111;
assign micromatrizz[92][386] = 9'b111111111;
assign micromatrizz[92][387] = 9'b111111111;
assign micromatrizz[92][388] = 9'b111111111;
assign micromatrizz[92][389] = 9'b111111111;
assign micromatrizz[92][390] = 9'b111111111;
assign micromatrizz[92][391] = 9'b111111111;
assign micromatrizz[92][392] = 9'b111111111;
assign micromatrizz[92][393] = 9'b111111111;
assign micromatrizz[92][394] = 9'b111111111;
assign micromatrizz[92][395] = 9'b111111111;
assign micromatrizz[92][396] = 9'b111111111;
assign micromatrizz[92][397] = 9'b111111111;
assign micromatrizz[92][398] = 9'b111111111;
assign micromatrizz[92][399] = 9'b111111111;
assign micromatrizz[92][400] = 9'b111111111;
assign micromatrizz[92][401] = 9'b111111111;
assign micromatrizz[92][402] = 9'b111111111;
assign micromatrizz[92][403] = 9'b111111111;
assign micromatrizz[92][404] = 9'b111111111;
assign micromatrizz[92][405] = 9'b111111111;
assign micromatrizz[92][406] = 9'b111111111;
assign micromatrizz[92][407] = 9'b111111111;
assign micromatrizz[92][408] = 9'b111111111;
assign micromatrizz[92][409] = 9'b111111111;
assign micromatrizz[92][410] = 9'b111111111;
assign micromatrizz[92][411] = 9'b111111111;
assign micromatrizz[92][412] = 9'b111111111;
assign micromatrizz[92][413] = 9'b111111111;
assign micromatrizz[92][414] = 9'b111111111;
assign micromatrizz[92][415] = 9'b111111111;
assign micromatrizz[92][416] = 9'b111111111;
assign micromatrizz[92][417] = 9'b111111111;
assign micromatrizz[92][418] = 9'b111111111;
assign micromatrizz[92][419] = 9'b111111111;
assign micromatrizz[92][420] = 9'b111111111;
assign micromatrizz[92][421] = 9'b111111111;
assign micromatrizz[92][422] = 9'b111111111;
assign micromatrizz[92][423] = 9'b111111111;
assign micromatrizz[92][424] = 9'b111111111;
assign micromatrizz[92][425] = 9'b111111111;
assign micromatrizz[92][426] = 9'b111111111;
assign micromatrizz[92][427] = 9'b111111111;
assign micromatrizz[92][428] = 9'b111111111;
assign micromatrizz[92][429] = 9'b111111111;
assign micromatrizz[92][430] = 9'b111111111;
assign micromatrizz[92][431] = 9'b111111111;
assign micromatrizz[92][432] = 9'b111111111;
assign micromatrizz[92][433] = 9'b111111111;
assign micromatrizz[92][434] = 9'b111111111;
assign micromatrizz[92][435] = 9'b111111111;
assign micromatrizz[92][436] = 9'b111111111;
assign micromatrizz[92][437] = 9'b111111111;
assign micromatrizz[92][438] = 9'b111111111;
assign micromatrizz[92][439] = 9'b111111111;
assign micromatrizz[92][440] = 9'b111111111;
assign micromatrizz[92][441] = 9'b111111111;
assign micromatrizz[92][442] = 9'b111111111;
assign micromatrizz[92][443] = 9'b111111111;
assign micromatrizz[92][444] = 9'b111111111;
assign micromatrizz[92][445] = 9'b111111111;
assign micromatrizz[92][446] = 9'b111111111;
assign micromatrizz[92][447] = 9'b111111111;
assign micromatrizz[92][448] = 9'b111111111;
assign micromatrizz[92][449] = 9'b111111111;
assign micromatrizz[92][450] = 9'b111111111;
assign micromatrizz[92][451] = 9'b111111111;
assign micromatrizz[92][452] = 9'b111111111;
assign micromatrizz[92][453] = 9'b111111111;
assign micromatrizz[92][454] = 9'b111111111;
assign micromatrizz[92][455] = 9'b111111111;
assign micromatrizz[92][456] = 9'b111111111;
assign micromatrizz[92][457] = 9'b111111111;
assign micromatrizz[92][458] = 9'b111111111;
assign micromatrizz[92][459] = 9'b111111111;
assign micromatrizz[92][460] = 9'b111111111;
assign micromatrizz[92][461] = 9'b111111111;
assign micromatrizz[92][462] = 9'b111111111;
assign micromatrizz[92][463] = 9'b111111111;
assign micromatrizz[92][464] = 9'b111111111;
assign micromatrizz[92][465] = 9'b111111111;
assign micromatrizz[92][466] = 9'b111111111;
assign micromatrizz[92][467] = 9'b111111111;
assign micromatrizz[92][468] = 9'b111111111;
assign micromatrizz[92][469] = 9'b111111111;
assign micromatrizz[92][470] = 9'b111111111;
assign micromatrizz[92][471] = 9'b111111111;
assign micromatrizz[92][472] = 9'b111111111;
assign micromatrizz[92][473] = 9'b111111111;
assign micromatrizz[92][474] = 9'b111111111;
assign micromatrizz[92][475] = 9'b111111111;
assign micromatrizz[92][476] = 9'b111111111;
assign micromatrizz[92][477] = 9'b111111111;
assign micromatrizz[92][478] = 9'b111111111;
assign micromatrizz[92][479] = 9'b111111111;
assign micromatrizz[92][480] = 9'b111111111;
assign micromatrizz[92][481] = 9'b111111111;
assign micromatrizz[92][482] = 9'b111111111;
assign micromatrizz[92][483] = 9'b111111111;
assign micromatrizz[92][484] = 9'b111111111;
assign micromatrizz[92][485] = 9'b111111111;
assign micromatrizz[92][486] = 9'b111111111;
assign micromatrizz[92][487] = 9'b111111111;
assign micromatrizz[92][488] = 9'b111111111;
assign micromatrizz[92][489] = 9'b111111111;
assign micromatrizz[92][490] = 9'b111111111;
assign micromatrizz[92][491] = 9'b111111111;
assign micromatrizz[92][492] = 9'b111111111;
assign micromatrizz[92][493] = 9'b111111111;
assign micromatrizz[92][494] = 9'b111111111;
assign micromatrizz[92][495] = 9'b111111111;
assign micromatrizz[92][496] = 9'b111111111;
assign micromatrizz[92][497] = 9'b111111111;
assign micromatrizz[92][498] = 9'b111111111;
assign micromatrizz[92][499] = 9'b111111111;
assign micromatrizz[92][500] = 9'b111111111;
assign micromatrizz[92][501] = 9'b111111111;
assign micromatrizz[92][502] = 9'b111111111;
assign micromatrizz[92][503] = 9'b111111111;
assign micromatrizz[92][504] = 9'b111111111;
assign micromatrizz[92][505] = 9'b111111111;
assign micromatrizz[92][506] = 9'b111111111;
assign micromatrizz[92][507] = 9'b111111111;
assign micromatrizz[92][508] = 9'b111111111;
assign micromatrizz[92][509] = 9'b111111111;
assign micromatrizz[92][510] = 9'b111111111;
assign micromatrizz[92][511] = 9'b111111111;
assign micromatrizz[92][512] = 9'b111111111;
assign micromatrizz[92][513] = 9'b111111111;
assign micromatrizz[92][514] = 9'b111111111;
assign micromatrizz[92][515] = 9'b111111111;
assign micromatrizz[92][516] = 9'b111111111;
assign micromatrizz[92][517] = 9'b111111111;
assign micromatrizz[92][518] = 9'b111111111;
assign micromatrizz[92][519] = 9'b111111111;
assign micromatrizz[92][520] = 9'b111111111;
assign micromatrizz[92][521] = 9'b111111111;
assign micromatrizz[92][522] = 9'b111111111;
assign micromatrizz[92][523] = 9'b111111111;
assign micromatrizz[92][524] = 9'b111111111;
assign micromatrizz[92][525] = 9'b111111111;
assign micromatrizz[92][526] = 9'b111111111;
assign micromatrizz[92][527] = 9'b111111111;
assign micromatrizz[92][528] = 9'b111111111;
assign micromatrizz[92][529] = 9'b111111111;
assign micromatrizz[92][530] = 9'b111111111;
assign micromatrizz[92][531] = 9'b111111111;
assign micromatrizz[92][532] = 9'b111111111;
assign micromatrizz[92][533] = 9'b111111111;
assign micromatrizz[92][534] = 9'b111111111;
assign micromatrizz[92][535] = 9'b111111111;
assign micromatrizz[92][536] = 9'b111111111;
assign micromatrizz[92][537] = 9'b111111111;
assign micromatrizz[92][538] = 9'b111111111;
assign micromatrizz[92][539] = 9'b111111111;
assign micromatrizz[92][540] = 9'b111111111;
assign micromatrizz[92][541] = 9'b111111111;
assign micromatrizz[92][542] = 9'b111111111;
assign micromatrizz[92][543] = 9'b111111111;
assign micromatrizz[92][544] = 9'b111111111;
assign micromatrizz[92][545] = 9'b111111111;
assign micromatrizz[92][546] = 9'b111111111;
assign micromatrizz[92][547] = 9'b111111111;
assign micromatrizz[92][548] = 9'b111111111;
assign micromatrizz[92][549] = 9'b111111111;
assign micromatrizz[92][550] = 9'b111111111;
assign micromatrizz[92][551] = 9'b111111111;
assign micromatrizz[92][552] = 9'b111111111;
assign micromatrizz[92][553] = 9'b111111111;
assign micromatrizz[92][554] = 9'b111111111;
assign micromatrizz[92][555] = 9'b111111111;
assign micromatrizz[92][556] = 9'b111111111;
assign micromatrizz[92][557] = 9'b111111111;
assign micromatrizz[92][558] = 9'b111111111;
assign micromatrizz[92][559] = 9'b111111111;
assign micromatrizz[92][560] = 9'b111111111;
assign micromatrizz[92][561] = 9'b111111111;
assign micromatrizz[92][562] = 9'b111111111;
assign micromatrizz[92][563] = 9'b111111111;
assign micromatrizz[92][564] = 9'b111111111;
assign micromatrizz[92][565] = 9'b111111111;
assign micromatrizz[92][566] = 9'b111111111;
assign micromatrizz[92][567] = 9'b111111111;
assign micromatrizz[92][568] = 9'b111111111;
assign micromatrizz[92][569] = 9'b111111111;
assign micromatrizz[92][570] = 9'b111111111;
assign micromatrizz[92][571] = 9'b111111111;
assign micromatrizz[92][572] = 9'b111111111;
assign micromatrizz[92][573] = 9'b111111111;
assign micromatrizz[92][574] = 9'b111111111;
assign micromatrizz[92][575] = 9'b111111111;
assign micromatrizz[92][576] = 9'b111111111;
assign micromatrizz[92][577] = 9'b111111111;
assign micromatrizz[92][578] = 9'b111111111;
assign micromatrizz[92][579] = 9'b111111111;
assign micromatrizz[92][580] = 9'b111111111;
assign micromatrizz[92][581] = 9'b111111111;
assign micromatrizz[92][582] = 9'b111111111;
assign micromatrizz[92][583] = 9'b111111111;
assign micromatrizz[92][584] = 9'b111111111;
assign micromatrizz[92][585] = 9'b111111111;
assign micromatrizz[92][586] = 9'b111111111;
assign micromatrizz[92][587] = 9'b111111111;
assign micromatrizz[92][588] = 9'b111111111;
assign micromatrizz[92][589] = 9'b111111111;
assign micromatrizz[92][590] = 9'b111111111;
assign micromatrizz[92][591] = 9'b111111111;
assign micromatrizz[92][592] = 9'b111111111;
assign micromatrizz[92][593] = 9'b111111111;
assign micromatrizz[92][594] = 9'b111111111;
assign micromatrizz[92][595] = 9'b111111111;
assign micromatrizz[92][596] = 9'b111111111;
assign micromatrizz[92][597] = 9'b111111111;
assign micromatrizz[92][598] = 9'b111111111;
assign micromatrizz[92][599] = 9'b111111111;
assign micromatrizz[92][600] = 9'b111111111;
assign micromatrizz[92][601] = 9'b111111111;
assign micromatrizz[92][602] = 9'b111111111;
assign micromatrizz[92][603] = 9'b111111111;
assign micromatrizz[92][604] = 9'b111111111;
assign micromatrizz[92][605] = 9'b111111111;
assign micromatrizz[92][606] = 9'b111111111;
assign micromatrizz[92][607] = 9'b111111111;
assign micromatrizz[92][608] = 9'b111111111;
assign micromatrizz[92][609] = 9'b111111111;
assign micromatrizz[92][610] = 9'b111111111;
assign micromatrizz[92][611] = 9'b111111111;
assign micromatrizz[92][612] = 9'b111111111;
assign micromatrizz[92][613] = 9'b111111111;
assign micromatrizz[92][614] = 9'b111111111;
assign micromatrizz[92][615] = 9'b111111111;
assign micromatrizz[92][616] = 9'b111111111;
assign micromatrizz[92][617] = 9'b111111111;
assign micromatrizz[92][618] = 9'b111111111;
assign micromatrizz[92][619] = 9'b111111111;
assign micromatrizz[92][620] = 9'b111111111;
assign micromatrizz[92][621] = 9'b111111111;
assign micromatrizz[92][622] = 9'b111111111;
assign micromatrizz[92][623] = 9'b111111111;
assign micromatrizz[92][624] = 9'b111111111;
assign micromatrizz[92][625] = 9'b111111111;
assign micromatrizz[92][626] = 9'b111111111;
assign micromatrizz[92][627] = 9'b111111111;
assign micromatrizz[92][628] = 9'b111111111;
assign micromatrizz[92][629] = 9'b111111111;
assign micromatrizz[92][630] = 9'b111111111;
assign micromatrizz[92][631] = 9'b111111111;
assign micromatrizz[92][632] = 9'b111111111;
assign micromatrizz[92][633] = 9'b111111111;
assign micromatrizz[92][634] = 9'b111111111;
assign micromatrizz[92][635] = 9'b111111111;
assign micromatrizz[92][636] = 9'b111111111;
assign micromatrizz[92][637] = 9'b111111111;
assign micromatrizz[92][638] = 9'b111111111;
assign micromatrizz[92][639] = 9'b111111111;
assign micromatrizz[93][0] = 9'b111111111;
assign micromatrizz[93][1] = 9'b111111111;
assign micromatrizz[93][2] = 9'b111111111;
assign micromatrizz[93][3] = 9'b111111111;
assign micromatrizz[93][4] = 9'b111111111;
assign micromatrizz[93][5] = 9'b111111111;
assign micromatrizz[93][6] = 9'b111111111;
assign micromatrizz[93][7] = 9'b111111111;
assign micromatrizz[93][8] = 9'b111111111;
assign micromatrizz[93][9] = 9'b111111111;
assign micromatrizz[93][10] = 9'b111111111;
assign micromatrizz[93][11] = 9'b111111111;
assign micromatrizz[93][12] = 9'b111111111;
assign micromatrizz[93][13] = 9'b111111111;
assign micromatrizz[93][14] = 9'b111111111;
assign micromatrizz[93][15] = 9'b111111111;
assign micromatrizz[93][16] = 9'b111111111;
assign micromatrizz[93][17] = 9'b111111111;
assign micromatrizz[93][18] = 9'b111111111;
assign micromatrizz[93][19] = 9'b111111111;
assign micromatrizz[93][20] = 9'b111111111;
assign micromatrizz[93][21] = 9'b111111111;
assign micromatrizz[93][22] = 9'b111111111;
assign micromatrizz[93][23] = 9'b111111111;
assign micromatrizz[93][24] = 9'b111111111;
assign micromatrizz[93][25] = 9'b111111111;
assign micromatrizz[93][26] = 9'b111111111;
assign micromatrizz[93][27] = 9'b111111111;
assign micromatrizz[93][28] = 9'b111111111;
assign micromatrizz[93][29] = 9'b111111111;
assign micromatrizz[93][30] = 9'b111111111;
assign micromatrizz[93][31] = 9'b111111111;
assign micromatrizz[93][32] = 9'b111111111;
assign micromatrizz[93][33] = 9'b111111111;
assign micromatrizz[93][34] = 9'b111111111;
assign micromatrizz[93][35] = 9'b111111111;
assign micromatrizz[93][36] = 9'b111111111;
assign micromatrizz[93][37] = 9'b111111111;
assign micromatrizz[93][38] = 9'b111111111;
assign micromatrizz[93][39] = 9'b111111111;
assign micromatrizz[93][40] = 9'b111111111;
assign micromatrizz[93][41] = 9'b111111111;
assign micromatrizz[93][42] = 9'b111111111;
assign micromatrizz[93][43] = 9'b111111111;
assign micromatrizz[93][44] = 9'b111111111;
assign micromatrizz[93][45] = 9'b111111111;
assign micromatrizz[93][46] = 9'b111111111;
assign micromatrizz[93][47] = 9'b111111111;
assign micromatrizz[93][48] = 9'b111111111;
assign micromatrizz[93][49] = 9'b111111111;
assign micromatrizz[93][50] = 9'b111111111;
assign micromatrizz[93][51] = 9'b111111111;
assign micromatrizz[93][52] = 9'b111111111;
assign micromatrizz[93][53] = 9'b111111111;
assign micromatrizz[93][54] = 9'b111111111;
assign micromatrizz[93][55] = 9'b111111111;
assign micromatrizz[93][56] = 9'b111111111;
assign micromatrizz[93][57] = 9'b111111111;
assign micromatrizz[93][58] = 9'b111111111;
assign micromatrizz[93][59] = 9'b111111111;
assign micromatrizz[93][60] = 9'b111111111;
assign micromatrizz[93][61] = 9'b111111111;
assign micromatrizz[93][62] = 9'b111111111;
assign micromatrizz[93][63] = 9'b111111111;
assign micromatrizz[93][64] = 9'b111111111;
assign micromatrizz[93][65] = 9'b111111111;
assign micromatrizz[93][66] = 9'b111111111;
assign micromatrizz[93][67] = 9'b111111111;
assign micromatrizz[93][68] = 9'b111111111;
assign micromatrizz[93][69] = 9'b111111111;
assign micromatrizz[93][70] = 9'b111111111;
assign micromatrizz[93][71] = 9'b111111111;
assign micromatrizz[93][72] = 9'b111111111;
assign micromatrizz[93][73] = 9'b111111111;
assign micromatrizz[93][74] = 9'b111111111;
assign micromatrizz[93][75] = 9'b111111111;
assign micromatrizz[93][76] = 9'b111111111;
assign micromatrizz[93][77] = 9'b111111111;
assign micromatrizz[93][78] = 9'b111111111;
assign micromatrizz[93][79] = 9'b111111111;
assign micromatrizz[93][80] = 9'b111111111;
assign micromatrizz[93][81] = 9'b111111111;
assign micromatrizz[93][82] = 9'b111111111;
assign micromatrizz[93][83] = 9'b111111111;
assign micromatrizz[93][84] = 9'b111111111;
assign micromatrizz[93][85] = 9'b111111111;
assign micromatrizz[93][86] = 9'b111111111;
assign micromatrizz[93][87] = 9'b111111111;
assign micromatrizz[93][88] = 9'b111111111;
assign micromatrizz[93][89] = 9'b111111111;
assign micromatrizz[93][90] = 9'b111111111;
assign micromatrizz[93][91] = 9'b111111111;
assign micromatrizz[93][92] = 9'b111111111;
assign micromatrizz[93][93] = 9'b111111111;
assign micromatrizz[93][94] = 9'b111111111;
assign micromatrizz[93][95] = 9'b111111111;
assign micromatrizz[93][96] = 9'b111111111;
assign micromatrizz[93][97] = 9'b111111111;
assign micromatrizz[93][98] = 9'b111111111;
assign micromatrizz[93][99] = 9'b111111111;
assign micromatrizz[93][100] = 9'b111111111;
assign micromatrizz[93][101] = 9'b111111111;
assign micromatrizz[93][102] = 9'b111111111;
assign micromatrizz[93][103] = 9'b111111111;
assign micromatrizz[93][104] = 9'b111111111;
assign micromatrizz[93][105] = 9'b111111111;
assign micromatrizz[93][106] = 9'b111111111;
assign micromatrizz[93][107] = 9'b111111111;
assign micromatrizz[93][108] = 9'b111111111;
assign micromatrizz[93][109] = 9'b111111111;
assign micromatrizz[93][110] = 9'b111111111;
assign micromatrizz[93][111] = 9'b111111111;
assign micromatrizz[93][112] = 9'b111111111;
assign micromatrizz[93][113] = 9'b111111111;
assign micromatrizz[93][114] = 9'b111111111;
assign micromatrizz[93][115] = 9'b111111111;
assign micromatrizz[93][116] = 9'b111111111;
assign micromatrizz[93][117] = 9'b111111111;
assign micromatrizz[93][118] = 9'b111111111;
assign micromatrizz[93][119] = 9'b111111111;
assign micromatrizz[93][120] = 9'b111111111;
assign micromatrizz[93][121] = 9'b111111111;
assign micromatrizz[93][122] = 9'b111111111;
assign micromatrizz[93][123] = 9'b111111111;
assign micromatrizz[93][124] = 9'b111111111;
assign micromatrizz[93][125] = 9'b111111111;
assign micromatrizz[93][126] = 9'b111111111;
assign micromatrizz[93][127] = 9'b111111111;
assign micromatrizz[93][128] = 9'b111111111;
assign micromatrizz[93][129] = 9'b111111111;
assign micromatrizz[93][130] = 9'b111111111;
assign micromatrizz[93][131] = 9'b111111111;
assign micromatrizz[93][132] = 9'b111111111;
assign micromatrizz[93][133] = 9'b111111111;
assign micromatrizz[93][134] = 9'b111111111;
assign micromatrizz[93][135] = 9'b111111111;
assign micromatrizz[93][136] = 9'b111111111;
assign micromatrizz[93][137] = 9'b111111111;
assign micromatrizz[93][138] = 9'b111111111;
assign micromatrizz[93][139] = 9'b111111111;
assign micromatrizz[93][140] = 9'b111111111;
assign micromatrizz[93][141] = 9'b111111111;
assign micromatrizz[93][142] = 9'b111111111;
assign micromatrizz[93][143] = 9'b111111111;
assign micromatrizz[93][144] = 9'b111111111;
assign micromatrizz[93][145] = 9'b111111111;
assign micromatrizz[93][146] = 9'b111111111;
assign micromatrizz[93][147] = 9'b111111111;
assign micromatrizz[93][148] = 9'b111111111;
assign micromatrizz[93][149] = 9'b111111111;
assign micromatrizz[93][150] = 9'b111111111;
assign micromatrizz[93][151] = 9'b111111111;
assign micromatrizz[93][152] = 9'b111111111;
assign micromatrizz[93][153] = 9'b111111111;
assign micromatrizz[93][154] = 9'b111111111;
assign micromatrizz[93][155] = 9'b111111111;
assign micromatrizz[93][156] = 9'b111111111;
assign micromatrizz[93][157] = 9'b111111111;
assign micromatrizz[93][158] = 9'b111111111;
assign micromatrizz[93][159] = 9'b111111111;
assign micromatrizz[93][160] = 9'b111111111;
assign micromatrizz[93][161] = 9'b111111111;
assign micromatrizz[93][162] = 9'b111111111;
assign micromatrizz[93][163] = 9'b111111111;
assign micromatrizz[93][164] = 9'b111111111;
assign micromatrizz[93][165] = 9'b111111111;
assign micromatrizz[93][166] = 9'b111111111;
assign micromatrizz[93][167] = 9'b111111111;
assign micromatrizz[93][168] = 9'b111111111;
assign micromatrizz[93][169] = 9'b111111111;
assign micromatrizz[93][170] = 9'b111111111;
assign micromatrizz[93][171] = 9'b111111111;
assign micromatrizz[93][172] = 9'b111111111;
assign micromatrizz[93][173] = 9'b111111111;
assign micromatrizz[93][174] = 9'b111111111;
assign micromatrizz[93][175] = 9'b111111111;
assign micromatrizz[93][176] = 9'b111111111;
assign micromatrizz[93][177] = 9'b111111111;
assign micromatrizz[93][178] = 9'b111111111;
assign micromatrizz[93][179] = 9'b111111111;
assign micromatrizz[93][180] = 9'b111111111;
assign micromatrizz[93][181] = 9'b111111111;
assign micromatrizz[93][182] = 9'b111111111;
assign micromatrizz[93][183] = 9'b111111111;
assign micromatrizz[93][184] = 9'b111111111;
assign micromatrizz[93][185] = 9'b111111111;
assign micromatrizz[93][186] = 9'b111111111;
assign micromatrizz[93][187] = 9'b111111111;
assign micromatrizz[93][188] = 9'b111111111;
assign micromatrizz[93][189] = 9'b111111111;
assign micromatrizz[93][190] = 9'b111111111;
assign micromatrizz[93][191] = 9'b111111111;
assign micromatrizz[93][192] = 9'b111111111;
assign micromatrizz[93][193] = 9'b111111111;
assign micromatrizz[93][194] = 9'b111111111;
assign micromatrizz[93][195] = 9'b111111111;
assign micromatrizz[93][196] = 9'b111111111;
assign micromatrizz[93][197] = 9'b111111111;
assign micromatrizz[93][198] = 9'b111111111;
assign micromatrizz[93][199] = 9'b111111111;
assign micromatrizz[93][200] = 9'b111111111;
assign micromatrizz[93][201] = 9'b111111111;
assign micromatrizz[93][202] = 9'b111111111;
assign micromatrizz[93][203] = 9'b111111111;
assign micromatrizz[93][204] = 9'b111111111;
assign micromatrizz[93][205] = 9'b111111111;
assign micromatrizz[93][206] = 9'b111111111;
assign micromatrizz[93][207] = 9'b111111111;
assign micromatrizz[93][208] = 9'b111111111;
assign micromatrizz[93][209] = 9'b111111111;
assign micromatrizz[93][210] = 9'b111111111;
assign micromatrizz[93][211] = 9'b111111111;
assign micromatrizz[93][212] = 9'b111111111;
assign micromatrizz[93][213] = 9'b111111111;
assign micromatrizz[93][214] = 9'b111111111;
assign micromatrizz[93][215] = 9'b111111111;
assign micromatrizz[93][216] = 9'b111111111;
assign micromatrizz[93][217] = 9'b111111111;
assign micromatrizz[93][218] = 9'b111111111;
assign micromatrizz[93][219] = 9'b111111111;
assign micromatrizz[93][220] = 9'b111111111;
assign micromatrizz[93][221] = 9'b111111111;
assign micromatrizz[93][222] = 9'b111111111;
assign micromatrizz[93][223] = 9'b111111111;
assign micromatrizz[93][224] = 9'b111111111;
assign micromatrizz[93][225] = 9'b111111111;
assign micromatrizz[93][226] = 9'b111111111;
assign micromatrizz[93][227] = 9'b111111111;
assign micromatrizz[93][228] = 9'b111111111;
assign micromatrizz[93][229] = 9'b111111111;
assign micromatrizz[93][230] = 9'b111111111;
assign micromatrizz[93][231] = 9'b111111111;
assign micromatrizz[93][232] = 9'b111111111;
assign micromatrizz[93][233] = 9'b111111111;
assign micromatrizz[93][234] = 9'b111111111;
assign micromatrizz[93][235] = 9'b111111111;
assign micromatrizz[93][236] = 9'b111111111;
assign micromatrizz[93][237] = 9'b111111111;
assign micromatrizz[93][238] = 9'b111111111;
assign micromatrizz[93][239] = 9'b111111111;
assign micromatrizz[93][240] = 9'b111111111;
assign micromatrizz[93][241] = 9'b111111111;
assign micromatrizz[93][242] = 9'b111111111;
assign micromatrizz[93][243] = 9'b111111111;
assign micromatrizz[93][244] = 9'b111111111;
assign micromatrizz[93][245] = 9'b111111111;
assign micromatrizz[93][246] = 9'b111111111;
assign micromatrizz[93][247] = 9'b111111111;
assign micromatrizz[93][248] = 9'b111111111;
assign micromatrizz[93][249] = 9'b111111111;
assign micromatrizz[93][250] = 9'b111111111;
assign micromatrizz[93][251] = 9'b111111111;
assign micromatrizz[93][252] = 9'b111111111;
assign micromatrizz[93][253] = 9'b111111111;
assign micromatrizz[93][254] = 9'b111111111;
assign micromatrizz[93][255] = 9'b111111111;
assign micromatrizz[93][256] = 9'b111111111;
assign micromatrizz[93][257] = 9'b111111111;
assign micromatrizz[93][258] = 9'b111111111;
assign micromatrizz[93][259] = 9'b111111111;
assign micromatrizz[93][260] = 9'b111111111;
assign micromatrizz[93][261] = 9'b111111111;
assign micromatrizz[93][262] = 9'b111111111;
assign micromatrizz[93][263] = 9'b111111111;
assign micromatrizz[93][264] = 9'b111111111;
assign micromatrizz[93][265] = 9'b111111111;
assign micromatrizz[93][266] = 9'b111111111;
assign micromatrizz[93][267] = 9'b111111111;
assign micromatrizz[93][268] = 9'b111111111;
assign micromatrizz[93][269] = 9'b111111111;
assign micromatrizz[93][270] = 9'b111111111;
assign micromatrizz[93][271] = 9'b111111111;
assign micromatrizz[93][272] = 9'b111111111;
assign micromatrizz[93][273] = 9'b111111111;
assign micromatrizz[93][274] = 9'b111111111;
assign micromatrizz[93][275] = 9'b111111111;
assign micromatrizz[93][276] = 9'b111111111;
assign micromatrizz[93][277] = 9'b111111111;
assign micromatrizz[93][278] = 9'b111111111;
assign micromatrizz[93][279] = 9'b111111111;
assign micromatrizz[93][280] = 9'b111111111;
assign micromatrizz[93][281] = 9'b111111111;
assign micromatrizz[93][282] = 9'b111111111;
assign micromatrizz[93][283] = 9'b111111111;
assign micromatrizz[93][284] = 9'b111111111;
assign micromatrizz[93][285] = 9'b111111111;
assign micromatrizz[93][286] = 9'b111111111;
assign micromatrizz[93][287] = 9'b111111111;
assign micromatrizz[93][288] = 9'b111111111;
assign micromatrizz[93][289] = 9'b111111111;
assign micromatrizz[93][290] = 9'b111111111;
assign micromatrizz[93][291] = 9'b111111111;
assign micromatrizz[93][292] = 9'b111111111;
assign micromatrizz[93][293] = 9'b111111111;
assign micromatrizz[93][294] = 9'b111111111;
assign micromatrizz[93][295] = 9'b111111111;
assign micromatrizz[93][296] = 9'b111111111;
assign micromatrizz[93][297] = 9'b111111111;
assign micromatrizz[93][298] = 9'b111111111;
assign micromatrizz[93][299] = 9'b111111111;
assign micromatrizz[93][300] = 9'b111111111;
assign micromatrizz[93][301] = 9'b111111111;
assign micromatrizz[93][302] = 9'b111111111;
assign micromatrizz[93][303] = 9'b111111111;
assign micromatrizz[93][304] = 9'b111111111;
assign micromatrizz[93][305] = 9'b111111111;
assign micromatrizz[93][306] = 9'b111111111;
assign micromatrizz[93][307] = 9'b111111111;
assign micromatrizz[93][308] = 9'b111111111;
assign micromatrizz[93][309] = 9'b111111111;
assign micromatrizz[93][310] = 9'b111111111;
assign micromatrizz[93][311] = 9'b111111111;
assign micromatrizz[93][312] = 9'b111111111;
assign micromatrizz[93][313] = 9'b111111111;
assign micromatrizz[93][314] = 9'b111111111;
assign micromatrizz[93][315] = 9'b111111111;
assign micromatrizz[93][316] = 9'b111111111;
assign micromatrizz[93][317] = 9'b111111111;
assign micromatrizz[93][318] = 9'b111111111;
assign micromatrizz[93][319] = 9'b111111111;
assign micromatrizz[93][320] = 9'b111111111;
assign micromatrizz[93][321] = 9'b111111111;
assign micromatrizz[93][322] = 9'b111111111;
assign micromatrizz[93][323] = 9'b111111111;
assign micromatrizz[93][324] = 9'b111111111;
assign micromatrizz[93][325] = 9'b111111111;
assign micromatrizz[93][326] = 9'b111111111;
assign micromatrizz[93][327] = 9'b111111111;
assign micromatrizz[93][328] = 9'b111111111;
assign micromatrizz[93][329] = 9'b111111111;
assign micromatrizz[93][330] = 9'b111111111;
assign micromatrizz[93][331] = 9'b111111111;
assign micromatrizz[93][332] = 9'b111111111;
assign micromatrizz[93][333] = 9'b111111111;
assign micromatrizz[93][334] = 9'b111111111;
assign micromatrizz[93][335] = 9'b111111111;
assign micromatrizz[93][336] = 9'b111111111;
assign micromatrizz[93][337] = 9'b111111111;
assign micromatrizz[93][338] = 9'b111111111;
assign micromatrizz[93][339] = 9'b111111111;
assign micromatrizz[93][340] = 9'b111111111;
assign micromatrizz[93][341] = 9'b111111111;
assign micromatrizz[93][342] = 9'b111111111;
assign micromatrizz[93][343] = 9'b111111111;
assign micromatrizz[93][344] = 9'b111111111;
assign micromatrizz[93][345] = 9'b111111111;
assign micromatrizz[93][346] = 9'b111111111;
assign micromatrizz[93][347] = 9'b111111111;
assign micromatrizz[93][348] = 9'b111111111;
assign micromatrizz[93][349] = 9'b111111111;
assign micromatrizz[93][350] = 9'b111111111;
assign micromatrizz[93][351] = 9'b111111111;
assign micromatrizz[93][352] = 9'b111111111;
assign micromatrizz[93][353] = 9'b111111111;
assign micromatrizz[93][354] = 9'b111111111;
assign micromatrizz[93][355] = 9'b111111111;
assign micromatrizz[93][356] = 9'b111111111;
assign micromatrizz[93][357] = 9'b111111111;
assign micromatrizz[93][358] = 9'b111111111;
assign micromatrizz[93][359] = 9'b111111111;
assign micromatrizz[93][360] = 9'b111111111;
assign micromatrizz[93][361] = 9'b111111111;
assign micromatrizz[93][362] = 9'b111111111;
assign micromatrizz[93][363] = 9'b111111111;
assign micromatrizz[93][364] = 9'b111111111;
assign micromatrizz[93][365] = 9'b111111111;
assign micromatrizz[93][366] = 9'b111111111;
assign micromatrizz[93][367] = 9'b111111111;
assign micromatrizz[93][368] = 9'b111111111;
assign micromatrizz[93][369] = 9'b111111111;
assign micromatrizz[93][370] = 9'b111111111;
assign micromatrizz[93][371] = 9'b111111111;
assign micromatrizz[93][372] = 9'b111111111;
assign micromatrizz[93][373] = 9'b111111111;
assign micromatrizz[93][374] = 9'b111111111;
assign micromatrizz[93][375] = 9'b111111111;
assign micromatrizz[93][376] = 9'b111111111;
assign micromatrizz[93][377] = 9'b111111111;
assign micromatrizz[93][378] = 9'b111111111;
assign micromatrizz[93][379] = 9'b111111111;
assign micromatrizz[93][380] = 9'b111111111;
assign micromatrizz[93][381] = 9'b111111111;
assign micromatrizz[93][382] = 9'b111111111;
assign micromatrizz[93][383] = 9'b111111111;
assign micromatrizz[93][384] = 9'b111111111;
assign micromatrizz[93][385] = 9'b111111111;
assign micromatrizz[93][386] = 9'b111111111;
assign micromatrizz[93][387] = 9'b111111111;
assign micromatrizz[93][388] = 9'b111111111;
assign micromatrizz[93][389] = 9'b111111111;
assign micromatrizz[93][390] = 9'b111111111;
assign micromatrizz[93][391] = 9'b111111111;
assign micromatrizz[93][392] = 9'b111111111;
assign micromatrizz[93][393] = 9'b111111111;
assign micromatrizz[93][394] = 9'b111111111;
assign micromatrizz[93][395] = 9'b111111111;
assign micromatrizz[93][396] = 9'b111111111;
assign micromatrizz[93][397] = 9'b111111111;
assign micromatrizz[93][398] = 9'b111111111;
assign micromatrizz[93][399] = 9'b111111111;
assign micromatrizz[93][400] = 9'b111111111;
assign micromatrizz[93][401] = 9'b111111111;
assign micromatrizz[93][402] = 9'b111111111;
assign micromatrizz[93][403] = 9'b111111111;
assign micromatrizz[93][404] = 9'b111111111;
assign micromatrizz[93][405] = 9'b111111111;
assign micromatrizz[93][406] = 9'b111111111;
assign micromatrizz[93][407] = 9'b111111111;
assign micromatrizz[93][408] = 9'b111111111;
assign micromatrizz[93][409] = 9'b111111111;
assign micromatrizz[93][410] = 9'b111111111;
assign micromatrizz[93][411] = 9'b111111111;
assign micromatrizz[93][412] = 9'b111111111;
assign micromatrizz[93][413] = 9'b111111111;
assign micromatrizz[93][414] = 9'b111111111;
assign micromatrizz[93][415] = 9'b111111111;
assign micromatrizz[93][416] = 9'b111111111;
assign micromatrizz[93][417] = 9'b111111111;
assign micromatrizz[93][418] = 9'b111111111;
assign micromatrizz[93][419] = 9'b111111111;
assign micromatrizz[93][420] = 9'b111111111;
assign micromatrizz[93][421] = 9'b111111111;
assign micromatrizz[93][422] = 9'b111111111;
assign micromatrizz[93][423] = 9'b111111111;
assign micromatrizz[93][424] = 9'b111111111;
assign micromatrizz[93][425] = 9'b111111111;
assign micromatrizz[93][426] = 9'b111111111;
assign micromatrizz[93][427] = 9'b111111111;
assign micromatrizz[93][428] = 9'b111111111;
assign micromatrizz[93][429] = 9'b111111111;
assign micromatrizz[93][430] = 9'b111111111;
assign micromatrizz[93][431] = 9'b111111111;
assign micromatrizz[93][432] = 9'b111111111;
assign micromatrizz[93][433] = 9'b111111111;
assign micromatrizz[93][434] = 9'b111111111;
assign micromatrizz[93][435] = 9'b111111111;
assign micromatrizz[93][436] = 9'b111111111;
assign micromatrizz[93][437] = 9'b111111111;
assign micromatrizz[93][438] = 9'b111111111;
assign micromatrizz[93][439] = 9'b111111111;
assign micromatrizz[93][440] = 9'b111111111;
assign micromatrizz[93][441] = 9'b111111111;
assign micromatrizz[93][442] = 9'b111111111;
assign micromatrizz[93][443] = 9'b111111111;
assign micromatrizz[93][444] = 9'b111111111;
assign micromatrizz[93][445] = 9'b111111111;
assign micromatrizz[93][446] = 9'b111111111;
assign micromatrizz[93][447] = 9'b111111111;
assign micromatrizz[93][448] = 9'b111111111;
assign micromatrizz[93][449] = 9'b111111111;
assign micromatrizz[93][450] = 9'b111111111;
assign micromatrizz[93][451] = 9'b111111111;
assign micromatrizz[93][452] = 9'b111111111;
assign micromatrizz[93][453] = 9'b111111111;
assign micromatrizz[93][454] = 9'b111111111;
assign micromatrizz[93][455] = 9'b111111111;
assign micromatrizz[93][456] = 9'b111111111;
assign micromatrizz[93][457] = 9'b111111111;
assign micromatrizz[93][458] = 9'b111111111;
assign micromatrizz[93][459] = 9'b111111111;
assign micromatrizz[93][460] = 9'b111111111;
assign micromatrizz[93][461] = 9'b111111111;
assign micromatrizz[93][462] = 9'b111111111;
assign micromatrizz[93][463] = 9'b111111111;
assign micromatrizz[93][464] = 9'b111111111;
assign micromatrizz[93][465] = 9'b111111111;
assign micromatrizz[93][466] = 9'b111111111;
assign micromatrizz[93][467] = 9'b111111111;
assign micromatrizz[93][468] = 9'b111111111;
assign micromatrizz[93][469] = 9'b111111111;
assign micromatrizz[93][470] = 9'b111111111;
assign micromatrizz[93][471] = 9'b111111111;
assign micromatrizz[93][472] = 9'b111111111;
assign micromatrizz[93][473] = 9'b111111111;
assign micromatrizz[93][474] = 9'b111111111;
assign micromatrizz[93][475] = 9'b111111111;
assign micromatrizz[93][476] = 9'b111111111;
assign micromatrizz[93][477] = 9'b111111111;
assign micromatrizz[93][478] = 9'b111111111;
assign micromatrizz[93][479] = 9'b111111111;
assign micromatrizz[93][480] = 9'b111111111;
assign micromatrizz[93][481] = 9'b111111111;
assign micromatrizz[93][482] = 9'b111111111;
assign micromatrizz[93][483] = 9'b111111111;
assign micromatrizz[93][484] = 9'b111111111;
assign micromatrizz[93][485] = 9'b111111111;
assign micromatrizz[93][486] = 9'b111111111;
assign micromatrizz[93][487] = 9'b111111111;
assign micromatrizz[93][488] = 9'b111111111;
assign micromatrizz[93][489] = 9'b111111111;
assign micromatrizz[93][490] = 9'b111111111;
assign micromatrizz[93][491] = 9'b111111111;
assign micromatrizz[93][492] = 9'b111111111;
assign micromatrizz[93][493] = 9'b111111111;
assign micromatrizz[93][494] = 9'b111111111;
assign micromatrizz[93][495] = 9'b111111111;
assign micromatrizz[93][496] = 9'b111111111;
assign micromatrizz[93][497] = 9'b111111111;
assign micromatrizz[93][498] = 9'b111111111;
assign micromatrizz[93][499] = 9'b111111111;
assign micromatrizz[93][500] = 9'b111111111;
assign micromatrizz[93][501] = 9'b111111111;
assign micromatrizz[93][502] = 9'b111111111;
assign micromatrizz[93][503] = 9'b111111111;
assign micromatrizz[93][504] = 9'b111111111;
assign micromatrizz[93][505] = 9'b111111111;
assign micromatrizz[93][506] = 9'b111111111;
assign micromatrizz[93][507] = 9'b111111111;
assign micromatrizz[93][508] = 9'b111111111;
assign micromatrizz[93][509] = 9'b111111111;
assign micromatrizz[93][510] = 9'b111111111;
assign micromatrizz[93][511] = 9'b111111111;
assign micromatrizz[93][512] = 9'b111111111;
assign micromatrizz[93][513] = 9'b111111111;
assign micromatrizz[93][514] = 9'b111111111;
assign micromatrizz[93][515] = 9'b111111111;
assign micromatrizz[93][516] = 9'b111111111;
assign micromatrizz[93][517] = 9'b111111111;
assign micromatrizz[93][518] = 9'b111111111;
assign micromatrizz[93][519] = 9'b111111111;
assign micromatrizz[93][520] = 9'b111111111;
assign micromatrizz[93][521] = 9'b111111111;
assign micromatrizz[93][522] = 9'b111111111;
assign micromatrizz[93][523] = 9'b111111111;
assign micromatrizz[93][524] = 9'b111111111;
assign micromatrizz[93][525] = 9'b111111111;
assign micromatrizz[93][526] = 9'b111111111;
assign micromatrizz[93][527] = 9'b111111111;
assign micromatrizz[93][528] = 9'b111111111;
assign micromatrizz[93][529] = 9'b111111111;
assign micromatrizz[93][530] = 9'b111111111;
assign micromatrizz[93][531] = 9'b111111111;
assign micromatrizz[93][532] = 9'b111111111;
assign micromatrizz[93][533] = 9'b111111111;
assign micromatrizz[93][534] = 9'b111111111;
assign micromatrizz[93][535] = 9'b111111111;
assign micromatrizz[93][536] = 9'b111111111;
assign micromatrizz[93][537] = 9'b111111111;
assign micromatrizz[93][538] = 9'b111111111;
assign micromatrizz[93][539] = 9'b111111111;
assign micromatrizz[93][540] = 9'b111111111;
assign micromatrizz[93][541] = 9'b111111111;
assign micromatrizz[93][542] = 9'b111111111;
assign micromatrizz[93][543] = 9'b111111111;
assign micromatrizz[93][544] = 9'b111111111;
assign micromatrizz[93][545] = 9'b111111111;
assign micromatrizz[93][546] = 9'b111111111;
assign micromatrizz[93][547] = 9'b111111111;
assign micromatrizz[93][548] = 9'b111111111;
assign micromatrizz[93][549] = 9'b111111111;
assign micromatrizz[93][550] = 9'b111111111;
assign micromatrizz[93][551] = 9'b111111111;
assign micromatrizz[93][552] = 9'b111111111;
assign micromatrizz[93][553] = 9'b111111111;
assign micromatrizz[93][554] = 9'b111111111;
assign micromatrizz[93][555] = 9'b111111111;
assign micromatrizz[93][556] = 9'b111111111;
assign micromatrizz[93][557] = 9'b111111111;
assign micromatrizz[93][558] = 9'b111111111;
assign micromatrizz[93][559] = 9'b111111111;
assign micromatrizz[93][560] = 9'b111111111;
assign micromatrizz[93][561] = 9'b111111111;
assign micromatrizz[93][562] = 9'b111111111;
assign micromatrizz[93][563] = 9'b111111111;
assign micromatrizz[93][564] = 9'b111111111;
assign micromatrizz[93][565] = 9'b111111111;
assign micromatrizz[93][566] = 9'b111111111;
assign micromatrizz[93][567] = 9'b111111111;
assign micromatrizz[93][568] = 9'b111111111;
assign micromatrizz[93][569] = 9'b111111111;
assign micromatrizz[93][570] = 9'b111111111;
assign micromatrizz[93][571] = 9'b111111111;
assign micromatrizz[93][572] = 9'b111111111;
assign micromatrizz[93][573] = 9'b111111111;
assign micromatrizz[93][574] = 9'b111111111;
assign micromatrizz[93][575] = 9'b111111111;
assign micromatrizz[93][576] = 9'b111111111;
assign micromatrizz[93][577] = 9'b111111111;
assign micromatrizz[93][578] = 9'b111111111;
assign micromatrizz[93][579] = 9'b111111111;
assign micromatrizz[93][580] = 9'b111111111;
assign micromatrizz[93][581] = 9'b111111111;
assign micromatrizz[93][582] = 9'b111111111;
assign micromatrizz[93][583] = 9'b111111111;
assign micromatrizz[93][584] = 9'b111111111;
assign micromatrizz[93][585] = 9'b111111111;
assign micromatrizz[93][586] = 9'b111111111;
assign micromatrizz[93][587] = 9'b111111111;
assign micromatrizz[93][588] = 9'b111111111;
assign micromatrizz[93][589] = 9'b111111111;
assign micromatrizz[93][590] = 9'b111111111;
assign micromatrizz[93][591] = 9'b111111111;
assign micromatrizz[93][592] = 9'b111111111;
assign micromatrizz[93][593] = 9'b111111111;
assign micromatrizz[93][594] = 9'b111111111;
assign micromatrizz[93][595] = 9'b111111111;
assign micromatrizz[93][596] = 9'b111111111;
assign micromatrizz[93][597] = 9'b111111111;
assign micromatrizz[93][598] = 9'b111111111;
assign micromatrizz[93][599] = 9'b111111111;
assign micromatrizz[93][600] = 9'b111111111;
assign micromatrizz[93][601] = 9'b111111111;
assign micromatrizz[93][602] = 9'b111111111;
assign micromatrizz[93][603] = 9'b111111111;
assign micromatrizz[93][604] = 9'b111111111;
assign micromatrizz[93][605] = 9'b111111111;
assign micromatrizz[93][606] = 9'b111111111;
assign micromatrizz[93][607] = 9'b111111111;
assign micromatrizz[93][608] = 9'b111111111;
assign micromatrizz[93][609] = 9'b111111111;
assign micromatrizz[93][610] = 9'b111111111;
assign micromatrizz[93][611] = 9'b111111111;
assign micromatrizz[93][612] = 9'b111111111;
assign micromatrizz[93][613] = 9'b111111111;
assign micromatrizz[93][614] = 9'b111111111;
assign micromatrizz[93][615] = 9'b111111111;
assign micromatrizz[93][616] = 9'b111111111;
assign micromatrizz[93][617] = 9'b111111111;
assign micromatrizz[93][618] = 9'b111111111;
assign micromatrizz[93][619] = 9'b111111111;
assign micromatrizz[93][620] = 9'b111111111;
assign micromatrizz[93][621] = 9'b111111111;
assign micromatrizz[93][622] = 9'b111111111;
assign micromatrizz[93][623] = 9'b111111111;
assign micromatrizz[93][624] = 9'b111111111;
assign micromatrizz[93][625] = 9'b111111111;
assign micromatrizz[93][626] = 9'b111111111;
assign micromatrizz[93][627] = 9'b111111111;
assign micromatrizz[93][628] = 9'b111111111;
assign micromatrizz[93][629] = 9'b111111111;
assign micromatrizz[93][630] = 9'b111111111;
assign micromatrizz[93][631] = 9'b111111111;
assign micromatrizz[93][632] = 9'b111111111;
assign micromatrizz[93][633] = 9'b111111111;
assign micromatrizz[93][634] = 9'b111111111;
assign micromatrizz[93][635] = 9'b111111111;
assign micromatrizz[93][636] = 9'b111111111;
assign micromatrizz[93][637] = 9'b111111111;
assign micromatrizz[93][638] = 9'b111111111;
assign micromatrizz[93][639] = 9'b111111111;
assign micromatrizz[94][0] = 9'b111111111;
assign micromatrizz[94][1] = 9'b111111111;
assign micromatrizz[94][2] = 9'b111111111;
assign micromatrizz[94][3] = 9'b111111111;
assign micromatrizz[94][4] = 9'b111111111;
assign micromatrizz[94][5] = 9'b111111111;
assign micromatrizz[94][6] = 9'b111111111;
assign micromatrizz[94][7] = 9'b111111111;
assign micromatrizz[94][8] = 9'b111111111;
assign micromatrizz[94][9] = 9'b111111111;
assign micromatrizz[94][10] = 9'b111111111;
assign micromatrizz[94][11] = 9'b111111111;
assign micromatrizz[94][12] = 9'b111111111;
assign micromatrizz[94][13] = 9'b111111111;
assign micromatrizz[94][14] = 9'b111111111;
assign micromatrizz[94][15] = 9'b111111111;
assign micromatrizz[94][16] = 9'b111111111;
assign micromatrizz[94][17] = 9'b111111111;
assign micromatrizz[94][18] = 9'b111111111;
assign micromatrizz[94][19] = 9'b111111111;
assign micromatrizz[94][20] = 9'b111111111;
assign micromatrizz[94][21] = 9'b111111111;
assign micromatrizz[94][22] = 9'b111111111;
assign micromatrizz[94][23] = 9'b111111111;
assign micromatrizz[94][24] = 9'b111111111;
assign micromatrizz[94][25] = 9'b111111111;
assign micromatrizz[94][26] = 9'b111111111;
assign micromatrizz[94][27] = 9'b111111111;
assign micromatrizz[94][28] = 9'b111111111;
assign micromatrizz[94][29] = 9'b111111111;
assign micromatrizz[94][30] = 9'b111111111;
assign micromatrizz[94][31] = 9'b111111111;
assign micromatrizz[94][32] = 9'b111111111;
assign micromatrizz[94][33] = 9'b111111111;
assign micromatrizz[94][34] = 9'b111111111;
assign micromatrizz[94][35] = 9'b111111111;
assign micromatrizz[94][36] = 9'b111111111;
assign micromatrizz[94][37] = 9'b111111111;
assign micromatrizz[94][38] = 9'b111111111;
assign micromatrizz[94][39] = 9'b111111111;
assign micromatrizz[94][40] = 9'b111111111;
assign micromatrizz[94][41] = 9'b111111111;
assign micromatrizz[94][42] = 9'b111111111;
assign micromatrizz[94][43] = 9'b111111111;
assign micromatrizz[94][44] = 9'b111111111;
assign micromatrizz[94][45] = 9'b111111111;
assign micromatrizz[94][46] = 9'b111111111;
assign micromatrizz[94][47] = 9'b111111111;
assign micromatrizz[94][48] = 9'b111111111;
assign micromatrizz[94][49] = 9'b111111111;
assign micromatrizz[94][50] = 9'b111111111;
assign micromatrizz[94][51] = 9'b111111111;
assign micromatrizz[94][52] = 9'b111111111;
assign micromatrizz[94][53] = 9'b111111111;
assign micromatrizz[94][54] = 9'b111111111;
assign micromatrizz[94][55] = 9'b111111111;
assign micromatrizz[94][56] = 9'b111111111;
assign micromatrizz[94][57] = 9'b111111111;
assign micromatrizz[94][58] = 9'b111111111;
assign micromatrizz[94][59] = 9'b111111111;
assign micromatrizz[94][60] = 9'b111111111;
assign micromatrizz[94][61] = 9'b111111111;
assign micromatrizz[94][62] = 9'b111111111;
assign micromatrizz[94][63] = 9'b111111111;
assign micromatrizz[94][64] = 9'b111111111;
assign micromatrizz[94][65] = 9'b111111111;
assign micromatrizz[94][66] = 9'b111111111;
assign micromatrizz[94][67] = 9'b111111111;
assign micromatrizz[94][68] = 9'b111111111;
assign micromatrizz[94][69] = 9'b111111111;
assign micromatrizz[94][70] = 9'b111111111;
assign micromatrizz[94][71] = 9'b111111111;
assign micromatrizz[94][72] = 9'b111111111;
assign micromatrizz[94][73] = 9'b111111111;
assign micromatrizz[94][74] = 9'b111111111;
assign micromatrizz[94][75] = 9'b111111111;
assign micromatrizz[94][76] = 9'b111111111;
assign micromatrizz[94][77] = 9'b111111111;
assign micromatrizz[94][78] = 9'b111111111;
assign micromatrizz[94][79] = 9'b111111111;
assign micromatrizz[94][80] = 9'b111111111;
assign micromatrizz[94][81] = 9'b111111111;
assign micromatrizz[94][82] = 9'b111111111;
assign micromatrizz[94][83] = 9'b111111111;
assign micromatrizz[94][84] = 9'b111111111;
assign micromatrizz[94][85] = 9'b111111111;
assign micromatrizz[94][86] = 9'b111111111;
assign micromatrizz[94][87] = 9'b111111111;
assign micromatrizz[94][88] = 9'b111111111;
assign micromatrizz[94][89] = 9'b111111111;
assign micromatrizz[94][90] = 9'b111111111;
assign micromatrizz[94][91] = 9'b111111111;
assign micromatrizz[94][92] = 9'b111111111;
assign micromatrizz[94][93] = 9'b111111111;
assign micromatrizz[94][94] = 9'b111111111;
assign micromatrizz[94][95] = 9'b111111111;
assign micromatrizz[94][96] = 9'b111111111;
assign micromatrizz[94][97] = 9'b111111111;
assign micromatrizz[94][98] = 9'b111111111;
assign micromatrizz[94][99] = 9'b111111111;
assign micromatrizz[94][100] = 9'b111111111;
assign micromatrizz[94][101] = 9'b111111111;
assign micromatrizz[94][102] = 9'b111111111;
assign micromatrizz[94][103] = 9'b111111111;
assign micromatrizz[94][104] = 9'b111111111;
assign micromatrizz[94][105] = 9'b111111111;
assign micromatrizz[94][106] = 9'b111111111;
assign micromatrizz[94][107] = 9'b111111111;
assign micromatrizz[94][108] = 9'b111111111;
assign micromatrizz[94][109] = 9'b111111111;
assign micromatrizz[94][110] = 9'b111111111;
assign micromatrizz[94][111] = 9'b111111111;
assign micromatrizz[94][112] = 9'b111111111;
assign micromatrizz[94][113] = 9'b111111111;
assign micromatrizz[94][114] = 9'b111111111;
assign micromatrizz[94][115] = 9'b111111111;
assign micromatrizz[94][116] = 9'b111111111;
assign micromatrizz[94][117] = 9'b111111111;
assign micromatrizz[94][118] = 9'b111111111;
assign micromatrizz[94][119] = 9'b111111111;
assign micromatrizz[94][120] = 9'b111111111;
assign micromatrizz[94][121] = 9'b111111111;
assign micromatrizz[94][122] = 9'b111111111;
assign micromatrizz[94][123] = 9'b111111111;
assign micromatrizz[94][124] = 9'b111111111;
assign micromatrizz[94][125] = 9'b111111111;
assign micromatrizz[94][126] = 9'b111111111;
assign micromatrizz[94][127] = 9'b111111111;
assign micromatrizz[94][128] = 9'b111111111;
assign micromatrizz[94][129] = 9'b111111111;
assign micromatrizz[94][130] = 9'b111111111;
assign micromatrizz[94][131] = 9'b111111111;
assign micromatrizz[94][132] = 9'b111111111;
assign micromatrizz[94][133] = 9'b111111111;
assign micromatrizz[94][134] = 9'b111111111;
assign micromatrizz[94][135] = 9'b111111111;
assign micromatrizz[94][136] = 9'b111111111;
assign micromatrizz[94][137] = 9'b111111111;
assign micromatrizz[94][138] = 9'b111111111;
assign micromatrizz[94][139] = 9'b111111111;
assign micromatrizz[94][140] = 9'b111111111;
assign micromatrizz[94][141] = 9'b111111111;
assign micromatrizz[94][142] = 9'b111111111;
assign micromatrizz[94][143] = 9'b111111111;
assign micromatrizz[94][144] = 9'b111111111;
assign micromatrizz[94][145] = 9'b111111111;
assign micromatrizz[94][146] = 9'b111111111;
assign micromatrizz[94][147] = 9'b111111111;
assign micromatrizz[94][148] = 9'b111111111;
assign micromatrizz[94][149] = 9'b111111111;
assign micromatrizz[94][150] = 9'b111111111;
assign micromatrizz[94][151] = 9'b111111111;
assign micromatrizz[94][152] = 9'b111111111;
assign micromatrizz[94][153] = 9'b111111111;
assign micromatrizz[94][154] = 9'b111111111;
assign micromatrizz[94][155] = 9'b111111111;
assign micromatrizz[94][156] = 9'b111111111;
assign micromatrizz[94][157] = 9'b111111111;
assign micromatrizz[94][158] = 9'b111111111;
assign micromatrizz[94][159] = 9'b111111111;
assign micromatrizz[94][160] = 9'b111111111;
assign micromatrizz[94][161] = 9'b111111111;
assign micromatrizz[94][162] = 9'b111111111;
assign micromatrizz[94][163] = 9'b111111111;
assign micromatrizz[94][164] = 9'b111111111;
assign micromatrizz[94][165] = 9'b111111111;
assign micromatrizz[94][166] = 9'b111111111;
assign micromatrizz[94][167] = 9'b111111111;
assign micromatrizz[94][168] = 9'b111111111;
assign micromatrizz[94][169] = 9'b111111111;
assign micromatrizz[94][170] = 9'b111111111;
assign micromatrizz[94][171] = 9'b111111111;
assign micromatrizz[94][172] = 9'b111111111;
assign micromatrizz[94][173] = 9'b111111111;
assign micromatrizz[94][174] = 9'b111111111;
assign micromatrizz[94][175] = 9'b111111111;
assign micromatrizz[94][176] = 9'b111111111;
assign micromatrizz[94][177] = 9'b111111111;
assign micromatrizz[94][178] = 9'b111111111;
assign micromatrizz[94][179] = 9'b111111111;
assign micromatrizz[94][180] = 9'b111111111;
assign micromatrizz[94][181] = 9'b111111111;
assign micromatrizz[94][182] = 9'b111111111;
assign micromatrizz[94][183] = 9'b111111111;
assign micromatrizz[94][184] = 9'b111111111;
assign micromatrizz[94][185] = 9'b111111111;
assign micromatrizz[94][186] = 9'b111111111;
assign micromatrizz[94][187] = 9'b111111111;
assign micromatrizz[94][188] = 9'b111111111;
assign micromatrizz[94][189] = 9'b111111111;
assign micromatrizz[94][190] = 9'b111111111;
assign micromatrizz[94][191] = 9'b111111111;
assign micromatrizz[94][192] = 9'b111111111;
assign micromatrizz[94][193] = 9'b111111111;
assign micromatrizz[94][194] = 9'b111111111;
assign micromatrizz[94][195] = 9'b111111111;
assign micromatrizz[94][196] = 9'b111111111;
assign micromatrizz[94][197] = 9'b111111111;
assign micromatrizz[94][198] = 9'b111111111;
assign micromatrizz[94][199] = 9'b111111111;
assign micromatrizz[94][200] = 9'b111111111;
assign micromatrizz[94][201] = 9'b111111111;
assign micromatrizz[94][202] = 9'b111111111;
assign micromatrizz[94][203] = 9'b111111111;
assign micromatrizz[94][204] = 9'b111111111;
assign micromatrizz[94][205] = 9'b111111111;
assign micromatrizz[94][206] = 9'b111111111;
assign micromatrizz[94][207] = 9'b111111111;
assign micromatrizz[94][208] = 9'b111111111;
assign micromatrizz[94][209] = 9'b111111111;
assign micromatrizz[94][210] = 9'b111111111;
assign micromatrizz[94][211] = 9'b111111111;
assign micromatrizz[94][212] = 9'b111111111;
assign micromatrizz[94][213] = 9'b111111111;
assign micromatrizz[94][214] = 9'b111111111;
assign micromatrizz[94][215] = 9'b111111111;
assign micromatrizz[94][216] = 9'b111111111;
assign micromatrizz[94][217] = 9'b111111111;
assign micromatrizz[94][218] = 9'b111111111;
assign micromatrizz[94][219] = 9'b111111111;
assign micromatrizz[94][220] = 9'b111111111;
assign micromatrizz[94][221] = 9'b111111111;
assign micromatrizz[94][222] = 9'b111111111;
assign micromatrizz[94][223] = 9'b111111111;
assign micromatrizz[94][224] = 9'b111111111;
assign micromatrizz[94][225] = 9'b111111111;
assign micromatrizz[94][226] = 9'b111111111;
assign micromatrizz[94][227] = 9'b111111111;
assign micromatrizz[94][228] = 9'b111111111;
assign micromatrizz[94][229] = 9'b111111111;
assign micromatrizz[94][230] = 9'b111111111;
assign micromatrizz[94][231] = 9'b111111111;
assign micromatrizz[94][232] = 9'b111111111;
assign micromatrizz[94][233] = 9'b111111111;
assign micromatrizz[94][234] = 9'b111111111;
assign micromatrizz[94][235] = 9'b111111111;
assign micromatrizz[94][236] = 9'b111111111;
assign micromatrizz[94][237] = 9'b111111111;
assign micromatrizz[94][238] = 9'b111111111;
assign micromatrizz[94][239] = 9'b111111111;
assign micromatrizz[94][240] = 9'b111111111;
assign micromatrizz[94][241] = 9'b111111111;
assign micromatrizz[94][242] = 9'b111111111;
assign micromatrizz[94][243] = 9'b111111111;
assign micromatrizz[94][244] = 9'b111111111;
assign micromatrizz[94][245] = 9'b111111111;
assign micromatrizz[94][246] = 9'b111111111;
assign micromatrizz[94][247] = 9'b111111111;
assign micromatrizz[94][248] = 9'b111111111;
assign micromatrizz[94][249] = 9'b111111111;
assign micromatrizz[94][250] = 9'b111111111;
assign micromatrizz[94][251] = 9'b111111111;
assign micromatrizz[94][252] = 9'b111111111;
assign micromatrizz[94][253] = 9'b111111111;
assign micromatrizz[94][254] = 9'b111111111;
assign micromatrizz[94][255] = 9'b111111111;
assign micromatrizz[94][256] = 9'b111111111;
assign micromatrizz[94][257] = 9'b111111111;
assign micromatrizz[94][258] = 9'b111111111;
assign micromatrizz[94][259] = 9'b111111111;
assign micromatrizz[94][260] = 9'b111111111;
assign micromatrizz[94][261] = 9'b111111111;
assign micromatrizz[94][262] = 9'b111111111;
assign micromatrizz[94][263] = 9'b111111111;
assign micromatrizz[94][264] = 9'b111111111;
assign micromatrizz[94][265] = 9'b111111111;
assign micromatrizz[94][266] = 9'b111111111;
assign micromatrizz[94][267] = 9'b111111111;
assign micromatrizz[94][268] = 9'b111111111;
assign micromatrizz[94][269] = 9'b111111111;
assign micromatrizz[94][270] = 9'b111111111;
assign micromatrizz[94][271] = 9'b111111111;
assign micromatrizz[94][272] = 9'b111111111;
assign micromatrizz[94][273] = 9'b111111111;
assign micromatrizz[94][274] = 9'b111111111;
assign micromatrizz[94][275] = 9'b111111111;
assign micromatrizz[94][276] = 9'b111111111;
assign micromatrizz[94][277] = 9'b111111111;
assign micromatrizz[94][278] = 9'b111111111;
assign micromatrizz[94][279] = 9'b111111111;
assign micromatrizz[94][280] = 9'b111111111;
assign micromatrizz[94][281] = 9'b111111111;
assign micromatrizz[94][282] = 9'b111111111;
assign micromatrizz[94][283] = 9'b111111111;
assign micromatrizz[94][284] = 9'b111111111;
assign micromatrizz[94][285] = 9'b111111111;
assign micromatrizz[94][286] = 9'b111111111;
assign micromatrizz[94][287] = 9'b111111111;
assign micromatrizz[94][288] = 9'b111111111;
assign micromatrizz[94][289] = 9'b111111111;
assign micromatrizz[94][290] = 9'b111111111;
assign micromatrizz[94][291] = 9'b111111111;
assign micromatrizz[94][292] = 9'b111111111;
assign micromatrizz[94][293] = 9'b111111111;
assign micromatrizz[94][294] = 9'b111111111;
assign micromatrizz[94][295] = 9'b111111111;
assign micromatrizz[94][296] = 9'b111111111;
assign micromatrizz[94][297] = 9'b111111111;
assign micromatrizz[94][298] = 9'b111111111;
assign micromatrizz[94][299] = 9'b111111111;
assign micromatrizz[94][300] = 9'b111111111;
assign micromatrizz[94][301] = 9'b111111111;
assign micromatrizz[94][302] = 9'b111111111;
assign micromatrizz[94][303] = 9'b111111111;
assign micromatrizz[94][304] = 9'b111111111;
assign micromatrizz[94][305] = 9'b111111111;
assign micromatrizz[94][306] = 9'b111111111;
assign micromatrizz[94][307] = 9'b111111111;
assign micromatrizz[94][308] = 9'b111111111;
assign micromatrizz[94][309] = 9'b111111111;
assign micromatrizz[94][310] = 9'b111111111;
assign micromatrizz[94][311] = 9'b111111111;
assign micromatrizz[94][312] = 9'b111111111;
assign micromatrizz[94][313] = 9'b111111111;
assign micromatrizz[94][314] = 9'b111111111;
assign micromatrizz[94][315] = 9'b111111111;
assign micromatrizz[94][316] = 9'b111111111;
assign micromatrizz[94][317] = 9'b111111111;
assign micromatrizz[94][318] = 9'b111111111;
assign micromatrizz[94][319] = 9'b111111111;
assign micromatrizz[94][320] = 9'b111111111;
assign micromatrizz[94][321] = 9'b111111111;
assign micromatrizz[94][322] = 9'b111111111;
assign micromatrizz[94][323] = 9'b111111111;
assign micromatrizz[94][324] = 9'b111111111;
assign micromatrizz[94][325] = 9'b111111111;
assign micromatrizz[94][326] = 9'b111111111;
assign micromatrizz[94][327] = 9'b111111111;
assign micromatrizz[94][328] = 9'b111111111;
assign micromatrizz[94][329] = 9'b111111111;
assign micromatrizz[94][330] = 9'b111111111;
assign micromatrizz[94][331] = 9'b111111111;
assign micromatrizz[94][332] = 9'b111111111;
assign micromatrizz[94][333] = 9'b111111111;
assign micromatrizz[94][334] = 9'b111111111;
assign micromatrizz[94][335] = 9'b111111111;
assign micromatrizz[94][336] = 9'b111111111;
assign micromatrizz[94][337] = 9'b111111111;
assign micromatrizz[94][338] = 9'b111111111;
assign micromatrizz[94][339] = 9'b111111111;
assign micromatrizz[94][340] = 9'b111111111;
assign micromatrizz[94][341] = 9'b111111111;
assign micromatrizz[94][342] = 9'b111111111;
assign micromatrizz[94][343] = 9'b111111111;
assign micromatrizz[94][344] = 9'b111111111;
assign micromatrizz[94][345] = 9'b111111111;
assign micromatrizz[94][346] = 9'b111111111;
assign micromatrizz[94][347] = 9'b111111111;
assign micromatrizz[94][348] = 9'b111111111;
assign micromatrizz[94][349] = 9'b111111111;
assign micromatrizz[94][350] = 9'b111111111;
assign micromatrizz[94][351] = 9'b111111111;
assign micromatrizz[94][352] = 9'b111111111;
assign micromatrizz[94][353] = 9'b111111111;
assign micromatrizz[94][354] = 9'b111111111;
assign micromatrizz[94][355] = 9'b111111111;
assign micromatrizz[94][356] = 9'b111111111;
assign micromatrizz[94][357] = 9'b111111111;
assign micromatrizz[94][358] = 9'b111111111;
assign micromatrizz[94][359] = 9'b111111111;
assign micromatrizz[94][360] = 9'b111111111;
assign micromatrizz[94][361] = 9'b111111111;
assign micromatrizz[94][362] = 9'b111111111;
assign micromatrizz[94][363] = 9'b111111111;
assign micromatrizz[94][364] = 9'b111111111;
assign micromatrizz[94][365] = 9'b111111111;
assign micromatrizz[94][366] = 9'b111111111;
assign micromatrizz[94][367] = 9'b111111111;
assign micromatrizz[94][368] = 9'b111111111;
assign micromatrizz[94][369] = 9'b111111111;
assign micromatrizz[94][370] = 9'b111111111;
assign micromatrizz[94][371] = 9'b111111111;
assign micromatrizz[94][372] = 9'b111111111;
assign micromatrizz[94][373] = 9'b111111111;
assign micromatrizz[94][374] = 9'b111111111;
assign micromatrizz[94][375] = 9'b111111111;
assign micromatrizz[94][376] = 9'b111111111;
assign micromatrizz[94][377] = 9'b111111111;
assign micromatrizz[94][378] = 9'b111111111;
assign micromatrizz[94][379] = 9'b111111111;
assign micromatrizz[94][380] = 9'b111111111;
assign micromatrizz[94][381] = 9'b111111111;
assign micromatrizz[94][382] = 9'b111111111;
assign micromatrizz[94][383] = 9'b111111111;
assign micromatrizz[94][384] = 9'b111111111;
assign micromatrizz[94][385] = 9'b111111111;
assign micromatrizz[94][386] = 9'b111111111;
assign micromatrizz[94][387] = 9'b111111111;
assign micromatrizz[94][388] = 9'b111111111;
assign micromatrizz[94][389] = 9'b111111111;
assign micromatrizz[94][390] = 9'b111111111;
assign micromatrizz[94][391] = 9'b111111111;
assign micromatrizz[94][392] = 9'b111111111;
assign micromatrizz[94][393] = 9'b111111111;
assign micromatrizz[94][394] = 9'b111111111;
assign micromatrizz[94][395] = 9'b111111111;
assign micromatrizz[94][396] = 9'b111111111;
assign micromatrizz[94][397] = 9'b111111111;
assign micromatrizz[94][398] = 9'b111111111;
assign micromatrizz[94][399] = 9'b111111111;
assign micromatrizz[94][400] = 9'b111111111;
assign micromatrizz[94][401] = 9'b111111111;
assign micromatrizz[94][402] = 9'b111111111;
assign micromatrizz[94][403] = 9'b111111111;
assign micromatrizz[94][404] = 9'b111111111;
assign micromatrizz[94][405] = 9'b111111111;
assign micromatrizz[94][406] = 9'b111111111;
assign micromatrizz[94][407] = 9'b111111111;
assign micromatrizz[94][408] = 9'b111111111;
assign micromatrizz[94][409] = 9'b111111111;
assign micromatrizz[94][410] = 9'b111111111;
assign micromatrizz[94][411] = 9'b111111111;
assign micromatrizz[94][412] = 9'b111111111;
assign micromatrizz[94][413] = 9'b111111111;
assign micromatrizz[94][414] = 9'b111111111;
assign micromatrizz[94][415] = 9'b111111111;
assign micromatrizz[94][416] = 9'b111111111;
assign micromatrizz[94][417] = 9'b111111111;
assign micromatrizz[94][418] = 9'b111111111;
assign micromatrizz[94][419] = 9'b111111111;
assign micromatrizz[94][420] = 9'b111111111;
assign micromatrizz[94][421] = 9'b111111111;
assign micromatrizz[94][422] = 9'b111111111;
assign micromatrizz[94][423] = 9'b111111111;
assign micromatrizz[94][424] = 9'b111111111;
assign micromatrizz[94][425] = 9'b111111111;
assign micromatrizz[94][426] = 9'b111111111;
assign micromatrizz[94][427] = 9'b111111111;
assign micromatrizz[94][428] = 9'b111111111;
assign micromatrizz[94][429] = 9'b111111111;
assign micromatrizz[94][430] = 9'b111111111;
assign micromatrizz[94][431] = 9'b111111111;
assign micromatrizz[94][432] = 9'b111111111;
assign micromatrizz[94][433] = 9'b111111111;
assign micromatrizz[94][434] = 9'b111111111;
assign micromatrizz[94][435] = 9'b111111111;
assign micromatrizz[94][436] = 9'b111111111;
assign micromatrizz[94][437] = 9'b111111111;
assign micromatrizz[94][438] = 9'b111111111;
assign micromatrizz[94][439] = 9'b111111111;
assign micromatrizz[94][440] = 9'b111111111;
assign micromatrizz[94][441] = 9'b111111111;
assign micromatrizz[94][442] = 9'b111111111;
assign micromatrizz[94][443] = 9'b111111111;
assign micromatrizz[94][444] = 9'b111111111;
assign micromatrizz[94][445] = 9'b111111111;
assign micromatrizz[94][446] = 9'b111111111;
assign micromatrizz[94][447] = 9'b111111111;
assign micromatrizz[94][448] = 9'b111111111;
assign micromatrizz[94][449] = 9'b111111111;
assign micromatrizz[94][450] = 9'b111111111;
assign micromatrizz[94][451] = 9'b111111111;
assign micromatrizz[94][452] = 9'b111111111;
assign micromatrizz[94][453] = 9'b111111111;
assign micromatrizz[94][454] = 9'b111111111;
assign micromatrizz[94][455] = 9'b111111111;
assign micromatrizz[94][456] = 9'b111111111;
assign micromatrizz[94][457] = 9'b111111111;
assign micromatrizz[94][458] = 9'b111111111;
assign micromatrizz[94][459] = 9'b111111111;
assign micromatrizz[94][460] = 9'b111111111;
assign micromatrizz[94][461] = 9'b111111111;
assign micromatrizz[94][462] = 9'b111111111;
assign micromatrizz[94][463] = 9'b111111111;
assign micromatrizz[94][464] = 9'b111111111;
assign micromatrizz[94][465] = 9'b111111111;
assign micromatrizz[94][466] = 9'b111111111;
assign micromatrizz[94][467] = 9'b111111111;
assign micromatrizz[94][468] = 9'b111111111;
assign micromatrizz[94][469] = 9'b111111111;
assign micromatrizz[94][470] = 9'b111111111;
assign micromatrizz[94][471] = 9'b111111111;
assign micromatrizz[94][472] = 9'b111111111;
assign micromatrizz[94][473] = 9'b111111111;
assign micromatrizz[94][474] = 9'b111111111;
assign micromatrizz[94][475] = 9'b111111111;
assign micromatrizz[94][476] = 9'b111111111;
assign micromatrizz[94][477] = 9'b111111111;
assign micromatrizz[94][478] = 9'b111111111;
assign micromatrizz[94][479] = 9'b111111111;
assign micromatrizz[94][480] = 9'b111111111;
assign micromatrizz[94][481] = 9'b111111111;
assign micromatrizz[94][482] = 9'b111111111;
assign micromatrizz[94][483] = 9'b111111111;
assign micromatrizz[94][484] = 9'b111111111;
assign micromatrizz[94][485] = 9'b111111111;
assign micromatrizz[94][486] = 9'b111111111;
assign micromatrizz[94][487] = 9'b111111111;
assign micromatrizz[94][488] = 9'b111111111;
assign micromatrizz[94][489] = 9'b111111111;
assign micromatrizz[94][490] = 9'b111111111;
assign micromatrizz[94][491] = 9'b111111111;
assign micromatrizz[94][492] = 9'b111111111;
assign micromatrizz[94][493] = 9'b111111111;
assign micromatrizz[94][494] = 9'b111111111;
assign micromatrizz[94][495] = 9'b111111111;
assign micromatrizz[94][496] = 9'b111111111;
assign micromatrizz[94][497] = 9'b111111111;
assign micromatrizz[94][498] = 9'b111111111;
assign micromatrizz[94][499] = 9'b111111111;
assign micromatrizz[94][500] = 9'b111111111;
assign micromatrizz[94][501] = 9'b111111111;
assign micromatrizz[94][502] = 9'b111111111;
assign micromatrizz[94][503] = 9'b111111111;
assign micromatrizz[94][504] = 9'b111111111;
assign micromatrizz[94][505] = 9'b111111111;
assign micromatrizz[94][506] = 9'b111111111;
assign micromatrizz[94][507] = 9'b111111111;
assign micromatrizz[94][508] = 9'b111111111;
assign micromatrizz[94][509] = 9'b111111111;
assign micromatrizz[94][510] = 9'b111111111;
assign micromatrizz[94][511] = 9'b111111111;
assign micromatrizz[94][512] = 9'b111111111;
assign micromatrizz[94][513] = 9'b111111111;
assign micromatrizz[94][514] = 9'b111111111;
assign micromatrizz[94][515] = 9'b111111111;
assign micromatrizz[94][516] = 9'b111111111;
assign micromatrizz[94][517] = 9'b111111111;
assign micromatrizz[94][518] = 9'b111111111;
assign micromatrizz[94][519] = 9'b111111111;
assign micromatrizz[94][520] = 9'b111111111;
assign micromatrizz[94][521] = 9'b111111111;
assign micromatrizz[94][522] = 9'b111111111;
assign micromatrizz[94][523] = 9'b111111111;
assign micromatrizz[94][524] = 9'b111111111;
assign micromatrizz[94][525] = 9'b111111111;
assign micromatrizz[94][526] = 9'b111111111;
assign micromatrizz[94][527] = 9'b111111111;
assign micromatrizz[94][528] = 9'b111111111;
assign micromatrizz[94][529] = 9'b111111111;
assign micromatrizz[94][530] = 9'b111111111;
assign micromatrizz[94][531] = 9'b111111111;
assign micromatrizz[94][532] = 9'b111111111;
assign micromatrizz[94][533] = 9'b111111111;
assign micromatrizz[94][534] = 9'b111111111;
assign micromatrizz[94][535] = 9'b111111111;
assign micromatrizz[94][536] = 9'b111111111;
assign micromatrizz[94][537] = 9'b111111111;
assign micromatrizz[94][538] = 9'b111111111;
assign micromatrizz[94][539] = 9'b111111111;
assign micromatrizz[94][540] = 9'b111111111;
assign micromatrizz[94][541] = 9'b111111111;
assign micromatrizz[94][542] = 9'b111111111;
assign micromatrizz[94][543] = 9'b111111111;
assign micromatrizz[94][544] = 9'b111111111;
assign micromatrizz[94][545] = 9'b111111111;
assign micromatrizz[94][546] = 9'b111111111;
assign micromatrizz[94][547] = 9'b111111111;
assign micromatrizz[94][548] = 9'b111111111;
assign micromatrizz[94][549] = 9'b111111111;
assign micromatrizz[94][550] = 9'b111111111;
assign micromatrizz[94][551] = 9'b111111111;
assign micromatrizz[94][552] = 9'b111111111;
assign micromatrizz[94][553] = 9'b111111111;
assign micromatrizz[94][554] = 9'b111111111;
assign micromatrizz[94][555] = 9'b111111111;
assign micromatrizz[94][556] = 9'b111111111;
assign micromatrizz[94][557] = 9'b111111111;
assign micromatrizz[94][558] = 9'b111111111;
assign micromatrizz[94][559] = 9'b111111111;
assign micromatrizz[94][560] = 9'b111111111;
assign micromatrizz[94][561] = 9'b111111111;
assign micromatrizz[94][562] = 9'b111111111;
assign micromatrizz[94][563] = 9'b111111111;
assign micromatrizz[94][564] = 9'b111111111;
assign micromatrizz[94][565] = 9'b111111111;
assign micromatrizz[94][566] = 9'b111111111;
assign micromatrizz[94][567] = 9'b111111111;
assign micromatrizz[94][568] = 9'b111111111;
assign micromatrizz[94][569] = 9'b111111111;
assign micromatrizz[94][570] = 9'b111111111;
assign micromatrizz[94][571] = 9'b111111111;
assign micromatrizz[94][572] = 9'b111111111;
assign micromatrizz[94][573] = 9'b111111111;
assign micromatrizz[94][574] = 9'b111111111;
assign micromatrizz[94][575] = 9'b111111111;
assign micromatrizz[94][576] = 9'b111111111;
assign micromatrizz[94][577] = 9'b111111111;
assign micromatrizz[94][578] = 9'b111111111;
assign micromatrizz[94][579] = 9'b111111111;
assign micromatrizz[94][580] = 9'b111111111;
assign micromatrizz[94][581] = 9'b111111111;
assign micromatrizz[94][582] = 9'b111111111;
assign micromatrizz[94][583] = 9'b111111111;
assign micromatrizz[94][584] = 9'b111111111;
assign micromatrizz[94][585] = 9'b111111111;
assign micromatrizz[94][586] = 9'b111111111;
assign micromatrizz[94][587] = 9'b111111111;
assign micromatrizz[94][588] = 9'b111111111;
assign micromatrizz[94][589] = 9'b111111111;
assign micromatrizz[94][590] = 9'b111111111;
assign micromatrizz[94][591] = 9'b111111111;
assign micromatrizz[94][592] = 9'b111111111;
assign micromatrizz[94][593] = 9'b111111111;
assign micromatrizz[94][594] = 9'b111111111;
assign micromatrizz[94][595] = 9'b111111111;
assign micromatrizz[94][596] = 9'b111111111;
assign micromatrizz[94][597] = 9'b111111111;
assign micromatrizz[94][598] = 9'b111111111;
assign micromatrizz[94][599] = 9'b111111111;
assign micromatrizz[94][600] = 9'b111111111;
assign micromatrizz[94][601] = 9'b111111111;
assign micromatrizz[94][602] = 9'b111111111;
assign micromatrizz[94][603] = 9'b111111111;
assign micromatrizz[94][604] = 9'b111111111;
assign micromatrizz[94][605] = 9'b111111111;
assign micromatrizz[94][606] = 9'b111111111;
assign micromatrizz[94][607] = 9'b111111111;
assign micromatrizz[94][608] = 9'b111111111;
assign micromatrizz[94][609] = 9'b111111111;
assign micromatrizz[94][610] = 9'b111111111;
assign micromatrizz[94][611] = 9'b111111111;
assign micromatrizz[94][612] = 9'b111111111;
assign micromatrizz[94][613] = 9'b111111111;
assign micromatrizz[94][614] = 9'b111111111;
assign micromatrizz[94][615] = 9'b111111111;
assign micromatrizz[94][616] = 9'b111111111;
assign micromatrizz[94][617] = 9'b111111111;
assign micromatrizz[94][618] = 9'b111111111;
assign micromatrizz[94][619] = 9'b111111111;
assign micromatrizz[94][620] = 9'b111111111;
assign micromatrizz[94][621] = 9'b111111111;
assign micromatrizz[94][622] = 9'b111111111;
assign micromatrizz[94][623] = 9'b111111111;
assign micromatrizz[94][624] = 9'b111111111;
assign micromatrizz[94][625] = 9'b111111111;
assign micromatrizz[94][626] = 9'b111111111;
assign micromatrizz[94][627] = 9'b111111111;
assign micromatrizz[94][628] = 9'b111111111;
assign micromatrizz[94][629] = 9'b111111111;
assign micromatrizz[94][630] = 9'b111111111;
assign micromatrizz[94][631] = 9'b111111111;
assign micromatrizz[94][632] = 9'b111111111;
assign micromatrizz[94][633] = 9'b111111111;
assign micromatrizz[94][634] = 9'b111111111;
assign micromatrizz[94][635] = 9'b111111111;
assign micromatrizz[94][636] = 9'b111111111;
assign micromatrizz[94][637] = 9'b111111111;
assign micromatrizz[94][638] = 9'b111111111;
assign micromatrizz[94][639] = 9'b111111111;
assign micromatrizz[95][0] = 9'b111111111;
assign micromatrizz[95][1] = 9'b111111111;
assign micromatrizz[95][2] = 9'b111111111;
assign micromatrizz[95][3] = 9'b111111111;
assign micromatrizz[95][4] = 9'b111111111;
assign micromatrizz[95][5] = 9'b111111111;
assign micromatrizz[95][6] = 9'b111111111;
assign micromatrizz[95][7] = 9'b111111111;
assign micromatrizz[95][8] = 9'b111111111;
assign micromatrizz[95][9] = 9'b111111111;
assign micromatrizz[95][10] = 9'b111111111;
assign micromatrizz[95][11] = 9'b111111111;
assign micromatrizz[95][12] = 9'b111111111;
assign micromatrizz[95][13] = 9'b111111111;
assign micromatrizz[95][14] = 9'b111111111;
assign micromatrizz[95][15] = 9'b111111111;
assign micromatrizz[95][16] = 9'b111111111;
assign micromatrizz[95][17] = 9'b111111111;
assign micromatrizz[95][18] = 9'b111111111;
assign micromatrizz[95][19] = 9'b111111111;
assign micromatrizz[95][20] = 9'b111111111;
assign micromatrizz[95][21] = 9'b111111111;
assign micromatrizz[95][22] = 9'b111111111;
assign micromatrizz[95][23] = 9'b111111111;
assign micromatrizz[95][24] = 9'b111111111;
assign micromatrizz[95][25] = 9'b111111111;
assign micromatrizz[95][26] = 9'b111111111;
assign micromatrizz[95][27] = 9'b111111111;
assign micromatrizz[95][28] = 9'b111111111;
assign micromatrizz[95][29] = 9'b111111111;
assign micromatrizz[95][30] = 9'b111111111;
assign micromatrizz[95][31] = 9'b111111111;
assign micromatrizz[95][32] = 9'b111111111;
assign micromatrizz[95][33] = 9'b111111111;
assign micromatrizz[95][34] = 9'b111111111;
assign micromatrizz[95][35] = 9'b111111111;
assign micromatrizz[95][36] = 9'b111111111;
assign micromatrizz[95][37] = 9'b111111111;
assign micromatrizz[95][38] = 9'b111111111;
assign micromatrizz[95][39] = 9'b111111111;
assign micromatrizz[95][40] = 9'b111111111;
assign micromatrizz[95][41] = 9'b111111111;
assign micromatrizz[95][42] = 9'b111111111;
assign micromatrizz[95][43] = 9'b111111111;
assign micromatrizz[95][44] = 9'b111111111;
assign micromatrizz[95][45] = 9'b111111111;
assign micromatrizz[95][46] = 9'b111111111;
assign micromatrizz[95][47] = 9'b111111111;
assign micromatrizz[95][48] = 9'b111111111;
assign micromatrizz[95][49] = 9'b111111111;
assign micromatrizz[95][50] = 9'b111111111;
assign micromatrizz[95][51] = 9'b111111111;
assign micromatrizz[95][52] = 9'b111111111;
assign micromatrizz[95][53] = 9'b111111111;
assign micromatrizz[95][54] = 9'b111111111;
assign micromatrizz[95][55] = 9'b111111111;
assign micromatrizz[95][56] = 9'b111111111;
assign micromatrizz[95][57] = 9'b111111111;
assign micromatrizz[95][58] = 9'b111111111;
assign micromatrizz[95][59] = 9'b111111111;
assign micromatrizz[95][60] = 9'b111111111;
assign micromatrizz[95][61] = 9'b111111111;
assign micromatrizz[95][62] = 9'b111111111;
assign micromatrizz[95][63] = 9'b111111111;
assign micromatrizz[95][64] = 9'b111111111;
assign micromatrizz[95][65] = 9'b111111111;
assign micromatrizz[95][66] = 9'b111111111;
assign micromatrizz[95][67] = 9'b111111111;
assign micromatrizz[95][68] = 9'b111111111;
assign micromatrizz[95][69] = 9'b111111111;
assign micromatrizz[95][70] = 9'b111111111;
assign micromatrizz[95][71] = 9'b111111111;
assign micromatrizz[95][72] = 9'b111111111;
assign micromatrizz[95][73] = 9'b111111111;
assign micromatrizz[95][74] = 9'b111111111;
assign micromatrizz[95][75] = 9'b111111111;
assign micromatrizz[95][76] = 9'b111111111;
assign micromatrizz[95][77] = 9'b111111111;
assign micromatrizz[95][78] = 9'b111111111;
assign micromatrizz[95][79] = 9'b111111111;
assign micromatrizz[95][80] = 9'b111111111;
assign micromatrizz[95][81] = 9'b111111111;
assign micromatrizz[95][82] = 9'b111111111;
assign micromatrizz[95][83] = 9'b111111111;
assign micromatrizz[95][84] = 9'b111111111;
assign micromatrizz[95][85] = 9'b111111111;
assign micromatrizz[95][86] = 9'b111111111;
assign micromatrizz[95][87] = 9'b111111111;
assign micromatrizz[95][88] = 9'b111111111;
assign micromatrizz[95][89] = 9'b111111111;
assign micromatrizz[95][90] = 9'b111111111;
assign micromatrizz[95][91] = 9'b111111111;
assign micromatrizz[95][92] = 9'b111111111;
assign micromatrizz[95][93] = 9'b111111111;
assign micromatrizz[95][94] = 9'b111111111;
assign micromatrizz[95][95] = 9'b111111111;
assign micromatrizz[95][96] = 9'b111111111;
assign micromatrizz[95][97] = 9'b111111111;
assign micromatrizz[95][98] = 9'b111111111;
assign micromatrizz[95][99] = 9'b111111111;
assign micromatrizz[95][100] = 9'b111111111;
assign micromatrizz[95][101] = 9'b111111111;
assign micromatrizz[95][102] = 9'b111111111;
assign micromatrizz[95][103] = 9'b111111111;
assign micromatrizz[95][104] = 9'b111111111;
assign micromatrizz[95][105] = 9'b111111111;
assign micromatrizz[95][106] = 9'b111111111;
assign micromatrizz[95][107] = 9'b111111111;
assign micromatrizz[95][108] = 9'b111111111;
assign micromatrizz[95][109] = 9'b111111111;
assign micromatrizz[95][110] = 9'b111111111;
assign micromatrizz[95][111] = 9'b111111111;
assign micromatrizz[95][112] = 9'b111111111;
assign micromatrizz[95][113] = 9'b111111111;
assign micromatrizz[95][114] = 9'b111111111;
assign micromatrizz[95][115] = 9'b111111111;
assign micromatrizz[95][116] = 9'b111111111;
assign micromatrizz[95][117] = 9'b111111111;
assign micromatrizz[95][118] = 9'b111111111;
assign micromatrizz[95][119] = 9'b111111111;
assign micromatrizz[95][120] = 9'b111111111;
assign micromatrizz[95][121] = 9'b111111111;
assign micromatrizz[95][122] = 9'b111111111;
assign micromatrizz[95][123] = 9'b111111111;
assign micromatrizz[95][124] = 9'b111111111;
assign micromatrizz[95][125] = 9'b111111111;
assign micromatrizz[95][126] = 9'b111111111;
assign micromatrizz[95][127] = 9'b111111111;
assign micromatrizz[95][128] = 9'b111111111;
assign micromatrizz[95][129] = 9'b111111111;
assign micromatrizz[95][130] = 9'b111111111;
assign micromatrizz[95][131] = 9'b111111111;
assign micromatrizz[95][132] = 9'b111111111;
assign micromatrizz[95][133] = 9'b111111111;
assign micromatrizz[95][134] = 9'b111111111;
assign micromatrizz[95][135] = 9'b111111111;
assign micromatrizz[95][136] = 9'b111111111;
assign micromatrizz[95][137] = 9'b111111111;
assign micromatrizz[95][138] = 9'b111111111;
assign micromatrizz[95][139] = 9'b111111111;
assign micromatrizz[95][140] = 9'b111111111;
assign micromatrizz[95][141] = 9'b111111111;
assign micromatrizz[95][142] = 9'b111111111;
assign micromatrizz[95][143] = 9'b111111111;
assign micromatrizz[95][144] = 9'b111111111;
assign micromatrizz[95][145] = 9'b111111111;
assign micromatrizz[95][146] = 9'b111111111;
assign micromatrizz[95][147] = 9'b111111111;
assign micromatrizz[95][148] = 9'b111111111;
assign micromatrizz[95][149] = 9'b111111111;
assign micromatrizz[95][150] = 9'b111111111;
assign micromatrizz[95][151] = 9'b111111111;
assign micromatrizz[95][152] = 9'b111111111;
assign micromatrizz[95][153] = 9'b111111111;
assign micromatrizz[95][154] = 9'b111111111;
assign micromatrizz[95][155] = 9'b111111111;
assign micromatrizz[95][156] = 9'b111111111;
assign micromatrizz[95][157] = 9'b111111111;
assign micromatrizz[95][158] = 9'b111111111;
assign micromatrizz[95][159] = 9'b111111111;
assign micromatrizz[95][160] = 9'b111111111;
assign micromatrizz[95][161] = 9'b111111111;
assign micromatrizz[95][162] = 9'b111111111;
assign micromatrizz[95][163] = 9'b111111111;
assign micromatrizz[95][164] = 9'b111111111;
assign micromatrizz[95][165] = 9'b111111111;
assign micromatrizz[95][166] = 9'b111111111;
assign micromatrizz[95][167] = 9'b111111111;
assign micromatrizz[95][168] = 9'b111111111;
assign micromatrizz[95][169] = 9'b111111111;
assign micromatrizz[95][170] = 9'b111111111;
assign micromatrizz[95][171] = 9'b111111111;
assign micromatrizz[95][172] = 9'b111111111;
assign micromatrizz[95][173] = 9'b111111111;
assign micromatrizz[95][174] = 9'b111111111;
assign micromatrizz[95][175] = 9'b111111111;
assign micromatrizz[95][176] = 9'b111111111;
assign micromatrizz[95][177] = 9'b111111111;
assign micromatrizz[95][178] = 9'b111111111;
assign micromatrizz[95][179] = 9'b111111111;
assign micromatrizz[95][180] = 9'b111111111;
assign micromatrizz[95][181] = 9'b111111111;
assign micromatrizz[95][182] = 9'b111111111;
assign micromatrizz[95][183] = 9'b111111111;
assign micromatrizz[95][184] = 9'b111111111;
assign micromatrizz[95][185] = 9'b111111111;
assign micromatrizz[95][186] = 9'b111111111;
assign micromatrizz[95][187] = 9'b111111111;
assign micromatrizz[95][188] = 9'b111111111;
assign micromatrizz[95][189] = 9'b111111111;
assign micromatrizz[95][190] = 9'b111111111;
assign micromatrizz[95][191] = 9'b111111111;
assign micromatrizz[95][192] = 9'b111111111;
assign micromatrizz[95][193] = 9'b111111111;
assign micromatrizz[95][194] = 9'b111111111;
assign micromatrizz[95][195] = 9'b111111111;
assign micromatrizz[95][196] = 9'b111111111;
assign micromatrizz[95][197] = 9'b111111111;
assign micromatrizz[95][198] = 9'b111111111;
assign micromatrizz[95][199] = 9'b111111111;
assign micromatrizz[95][200] = 9'b111111111;
assign micromatrizz[95][201] = 9'b111111111;
assign micromatrizz[95][202] = 9'b111111111;
assign micromatrizz[95][203] = 9'b111111111;
assign micromatrizz[95][204] = 9'b111111111;
assign micromatrizz[95][205] = 9'b111111111;
assign micromatrizz[95][206] = 9'b111111111;
assign micromatrizz[95][207] = 9'b111111111;
assign micromatrizz[95][208] = 9'b111111111;
assign micromatrizz[95][209] = 9'b111111111;
assign micromatrizz[95][210] = 9'b111111111;
assign micromatrizz[95][211] = 9'b111111111;
assign micromatrizz[95][212] = 9'b111111111;
assign micromatrizz[95][213] = 9'b111111111;
assign micromatrizz[95][214] = 9'b111111111;
assign micromatrizz[95][215] = 9'b111111111;
assign micromatrizz[95][216] = 9'b111111111;
assign micromatrizz[95][217] = 9'b111111111;
assign micromatrizz[95][218] = 9'b111111111;
assign micromatrizz[95][219] = 9'b111111111;
assign micromatrizz[95][220] = 9'b111111111;
assign micromatrizz[95][221] = 9'b111111111;
assign micromatrizz[95][222] = 9'b111111111;
assign micromatrizz[95][223] = 9'b111111111;
assign micromatrizz[95][224] = 9'b111111111;
assign micromatrizz[95][225] = 9'b111111111;
assign micromatrizz[95][226] = 9'b111111111;
assign micromatrizz[95][227] = 9'b111111111;
assign micromatrizz[95][228] = 9'b111111111;
assign micromatrizz[95][229] = 9'b111111111;
assign micromatrizz[95][230] = 9'b111111111;
assign micromatrizz[95][231] = 9'b111111111;
assign micromatrizz[95][232] = 9'b111111111;
assign micromatrizz[95][233] = 9'b111111111;
assign micromatrizz[95][234] = 9'b111111111;
assign micromatrizz[95][235] = 9'b111111111;
assign micromatrizz[95][236] = 9'b111111111;
assign micromatrizz[95][237] = 9'b111111111;
assign micromatrizz[95][238] = 9'b111111111;
assign micromatrizz[95][239] = 9'b111111111;
assign micromatrizz[95][240] = 9'b111111111;
assign micromatrizz[95][241] = 9'b111111111;
assign micromatrizz[95][242] = 9'b111111111;
assign micromatrizz[95][243] = 9'b111111111;
assign micromatrizz[95][244] = 9'b111111111;
assign micromatrizz[95][245] = 9'b111111111;
assign micromatrizz[95][246] = 9'b111111111;
assign micromatrizz[95][247] = 9'b111111111;
assign micromatrizz[95][248] = 9'b111111111;
assign micromatrizz[95][249] = 9'b111111111;
assign micromatrizz[95][250] = 9'b111111111;
assign micromatrizz[95][251] = 9'b111111111;
assign micromatrizz[95][252] = 9'b111111111;
assign micromatrizz[95][253] = 9'b111111111;
assign micromatrizz[95][254] = 9'b111111111;
assign micromatrizz[95][255] = 9'b111111111;
assign micromatrizz[95][256] = 9'b111111111;
assign micromatrizz[95][257] = 9'b111111111;
assign micromatrizz[95][258] = 9'b111111111;
assign micromatrizz[95][259] = 9'b111111111;
assign micromatrizz[95][260] = 9'b111111111;
assign micromatrizz[95][261] = 9'b111111111;
assign micromatrizz[95][262] = 9'b111111111;
assign micromatrizz[95][263] = 9'b111111111;
assign micromatrizz[95][264] = 9'b111111111;
assign micromatrizz[95][265] = 9'b111111111;
assign micromatrizz[95][266] = 9'b111111111;
assign micromatrizz[95][267] = 9'b111111111;
assign micromatrizz[95][268] = 9'b111111111;
assign micromatrizz[95][269] = 9'b111111111;
assign micromatrizz[95][270] = 9'b111111111;
assign micromatrizz[95][271] = 9'b111111111;
assign micromatrizz[95][272] = 9'b111111111;
assign micromatrizz[95][273] = 9'b111111111;
assign micromatrizz[95][274] = 9'b111111111;
assign micromatrizz[95][275] = 9'b111111111;
assign micromatrizz[95][276] = 9'b111111111;
assign micromatrizz[95][277] = 9'b111111111;
assign micromatrizz[95][278] = 9'b111111111;
assign micromatrizz[95][279] = 9'b111111111;
assign micromatrizz[95][280] = 9'b111111111;
assign micromatrizz[95][281] = 9'b111111111;
assign micromatrizz[95][282] = 9'b111111111;
assign micromatrizz[95][283] = 9'b111111111;
assign micromatrizz[95][284] = 9'b111111111;
assign micromatrizz[95][285] = 9'b111111111;
assign micromatrizz[95][286] = 9'b111111111;
assign micromatrizz[95][287] = 9'b111111111;
assign micromatrizz[95][288] = 9'b111111111;
assign micromatrizz[95][289] = 9'b111111111;
assign micromatrizz[95][290] = 9'b111111111;
assign micromatrizz[95][291] = 9'b111111111;
assign micromatrizz[95][292] = 9'b111111111;
assign micromatrizz[95][293] = 9'b111111111;
assign micromatrizz[95][294] = 9'b111111111;
assign micromatrizz[95][295] = 9'b111111111;
assign micromatrizz[95][296] = 9'b111111111;
assign micromatrizz[95][297] = 9'b111111111;
assign micromatrizz[95][298] = 9'b111111111;
assign micromatrizz[95][299] = 9'b111111111;
assign micromatrizz[95][300] = 9'b111111111;
assign micromatrizz[95][301] = 9'b111111111;
assign micromatrizz[95][302] = 9'b111111111;
assign micromatrizz[95][303] = 9'b111111111;
assign micromatrizz[95][304] = 9'b111111111;
assign micromatrizz[95][305] = 9'b111111111;
assign micromatrizz[95][306] = 9'b111111111;
assign micromatrizz[95][307] = 9'b111111111;
assign micromatrizz[95][308] = 9'b111111111;
assign micromatrizz[95][309] = 9'b111111111;
assign micromatrizz[95][310] = 9'b111111111;
assign micromatrizz[95][311] = 9'b111111111;
assign micromatrizz[95][312] = 9'b111111111;
assign micromatrizz[95][313] = 9'b111111111;
assign micromatrizz[95][314] = 9'b111111111;
assign micromatrizz[95][315] = 9'b111111111;
assign micromatrizz[95][316] = 9'b111111111;
assign micromatrizz[95][317] = 9'b111111111;
assign micromatrizz[95][318] = 9'b111111111;
assign micromatrizz[95][319] = 9'b111111111;
assign micromatrizz[95][320] = 9'b111111111;
assign micromatrizz[95][321] = 9'b111111111;
assign micromatrizz[95][322] = 9'b111111111;
assign micromatrizz[95][323] = 9'b111111111;
assign micromatrizz[95][324] = 9'b111111111;
assign micromatrizz[95][325] = 9'b111111111;
assign micromatrizz[95][326] = 9'b111111111;
assign micromatrizz[95][327] = 9'b111111111;
assign micromatrizz[95][328] = 9'b111111111;
assign micromatrizz[95][329] = 9'b111111111;
assign micromatrizz[95][330] = 9'b111111111;
assign micromatrizz[95][331] = 9'b111111111;
assign micromatrizz[95][332] = 9'b111111111;
assign micromatrizz[95][333] = 9'b111111111;
assign micromatrizz[95][334] = 9'b111111111;
assign micromatrizz[95][335] = 9'b111111111;
assign micromatrizz[95][336] = 9'b111111111;
assign micromatrizz[95][337] = 9'b111111111;
assign micromatrizz[95][338] = 9'b111111111;
assign micromatrizz[95][339] = 9'b111111111;
assign micromatrizz[95][340] = 9'b111111111;
assign micromatrizz[95][341] = 9'b111111111;
assign micromatrizz[95][342] = 9'b111111111;
assign micromatrizz[95][343] = 9'b111111111;
assign micromatrizz[95][344] = 9'b111111111;
assign micromatrizz[95][345] = 9'b111111111;
assign micromatrizz[95][346] = 9'b111111111;
assign micromatrizz[95][347] = 9'b111111111;
assign micromatrizz[95][348] = 9'b111111111;
assign micromatrizz[95][349] = 9'b111111111;
assign micromatrizz[95][350] = 9'b111111111;
assign micromatrizz[95][351] = 9'b111111111;
assign micromatrizz[95][352] = 9'b111111111;
assign micromatrizz[95][353] = 9'b111111111;
assign micromatrizz[95][354] = 9'b111111111;
assign micromatrizz[95][355] = 9'b111111111;
assign micromatrizz[95][356] = 9'b111111111;
assign micromatrizz[95][357] = 9'b111111111;
assign micromatrizz[95][358] = 9'b111111111;
assign micromatrizz[95][359] = 9'b111111111;
assign micromatrizz[95][360] = 9'b111111111;
assign micromatrizz[95][361] = 9'b111111111;
assign micromatrizz[95][362] = 9'b111111111;
assign micromatrizz[95][363] = 9'b111111111;
assign micromatrizz[95][364] = 9'b111111111;
assign micromatrizz[95][365] = 9'b111111111;
assign micromatrizz[95][366] = 9'b111111111;
assign micromatrizz[95][367] = 9'b111111111;
assign micromatrizz[95][368] = 9'b111111111;
assign micromatrizz[95][369] = 9'b111111111;
assign micromatrizz[95][370] = 9'b111111111;
assign micromatrizz[95][371] = 9'b111111111;
assign micromatrizz[95][372] = 9'b111111111;
assign micromatrizz[95][373] = 9'b111111111;
assign micromatrizz[95][374] = 9'b111111111;
assign micromatrizz[95][375] = 9'b111111111;
assign micromatrizz[95][376] = 9'b111111111;
assign micromatrizz[95][377] = 9'b111111111;
assign micromatrizz[95][378] = 9'b111111111;
assign micromatrizz[95][379] = 9'b111111111;
assign micromatrizz[95][380] = 9'b111111111;
assign micromatrizz[95][381] = 9'b111111111;
assign micromatrizz[95][382] = 9'b111111111;
assign micromatrizz[95][383] = 9'b111111111;
assign micromatrizz[95][384] = 9'b111111111;
assign micromatrizz[95][385] = 9'b111111111;
assign micromatrizz[95][386] = 9'b111111111;
assign micromatrizz[95][387] = 9'b111111111;
assign micromatrizz[95][388] = 9'b111111111;
assign micromatrizz[95][389] = 9'b111111111;
assign micromatrizz[95][390] = 9'b111111111;
assign micromatrizz[95][391] = 9'b111111111;
assign micromatrizz[95][392] = 9'b111111111;
assign micromatrizz[95][393] = 9'b111111111;
assign micromatrizz[95][394] = 9'b111111111;
assign micromatrizz[95][395] = 9'b111111111;
assign micromatrizz[95][396] = 9'b111111111;
assign micromatrizz[95][397] = 9'b111111111;
assign micromatrizz[95][398] = 9'b111111111;
assign micromatrizz[95][399] = 9'b111111111;
assign micromatrizz[95][400] = 9'b111111111;
assign micromatrizz[95][401] = 9'b111111111;
assign micromatrizz[95][402] = 9'b111111111;
assign micromatrizz[95][403] = 9'b111111111;
assign micromatrizz[95][404] = 9'b111111111;
assign micromatrizz[95][405] = 9'b111111111;
assign micromatrizz[95][406] = 9'b111111111;
assign micromatrizz[95][407] = 9'b111111111;
assign micromatrizz[95][408] = 9'b111111111;
assign micromatrizz[95][409] = 9'b111111111;
assign micromatrizz[95][410] = 9'b111111111;
assign micromatrizz[95][411] = 9'b111111111;
assign micromatrizz[95][412] = 9'b111111111;
assign micromatrizz[95][413] = 9'b111111111;
assign micromatrizz[95][414] = 9'b111111111;
assign micromatrizz[95][415] = 9'b111111111;
assign micromatrizz[95][416] = 9'b111111111;
assign micromatrizz[95][417] = 9'b111111111;
assign micromatrizz[95][418] = 9'b111111111;
assign micromatrizz[95][419] = 9'b111111111;
assign micromatrizz[95][420] = 9'b111111111;
assign micromatrizz[95][421] = 9'b111111111;
assign micromatrizz[95][422] = 9'b111111111;
assign micromatrizz[95][423] = 9'b111111111;
assign micromatrizz[95][424] = 9'b111111111;
assign micromatrizz[95][425] = 9'b111111111;
assign micromatrizz[95][426] = 9'b111111111;
assign micromatrizz[95][427] = 9'b111111111;
assign micromatrizz[95][428] = 9'b111111111;
assign micromatrizz[95][429] = 9'b111111111;
assign micromatrizz[95][430] = 9'b111111111;
assign micromatrizz[95][431] = 9'b111111111;
assign micromatrizz[95][432] = 9'b111111111;
assign micromatrizz[95][433] = 9'b111111111;
assign micromatrizz[95][434] = 9'b111111111;
assign micromatrizz[95][435] = 9'b111111111;
assign micromatrizz[95][436] = 9'b111111111;
assign micromatrizz[95][437] = 9'b111111111;
assign micromatrizz[95][438] = 9'b111111111;
assign micromatrizz[95][439] = 9'b111111111;
assign micromatrizz[95][440] = 9'b111111111;
assign micromatrizz[95][441] = 9'b111111111;
assign micromatrizz[95][442] = 9'b111111111;
assign micromatrizz[95][443] = 9'b111111111;
assign micromatrizz[95][444] = 9'b111111111;
assign micromatrizz[95][445] = 9'b111111111;
assign micromatrizz[95][446] = 9'b111111111;
assign micromatrizz[95][447] = 9'b111111111;
assign micromatrizz[95][448] = 9'b111111111;
assign micromatrizz[95][449] = 9'b111111111;
assign micromatrizz[95][450] = 9'b111111111;
assign micromatrizz[95][451] = 9'b111111111;
assign micromatrizz[95][452] = 9'b111111111;
assign micromatrizz[95][453] = 9'b111111111;
assign micromatrizz[95][454] = 9'b111111111;
assign micromatrizz[95][455] = 9'b111111111;
assign micromatrizz[95][456] = 9'b111111111;
assign micromatrizz[95][457] = 9'b111111111;
assign micromatrizz[95][458] = 9'b111111111;
assign micromatrizz[95][459] = 9'b111111111;
assign micromatrizz[95][460] = 9'b111111111;
assign micromatrizz[95][461] = 9'b111111111;
assign micromatrizz[95][462] = 9'b111111111;
assign micromatrizz[95][463] = 9'b111111111;
assign micromatrizz[95][464] = 9'b111111111;
assign micromatrizz[95][465] = 9'b111111111;
assign micromatrizz[95][466] = 9'b111111111;
assign micromatrizz[95][467] = 9'b111111111;
assign micromatrizz[95][468] = 9'b111111111;
assign micromatrizz[95][469] = 9'b111111111;
assign micromatrizz[95][470] = 9'b111111111;
assign micromatrizz[95][471] = 9'b111111111;
assign micromatrizz[95][472] = 9'b111111111;
assign micromatrizz[95][473] = 9'b111111111;
assign micromatrizz[95][474] = 9'b111111111;
assign micromatrizz[95][475] = 9'b111111111;
assign micromatrizz[95][476] = 9'b111111111;
assign micromatrizz[95][477] = 9'b111111111;
assign micromatrizz[95][478] = 9'b111111111;
assign micromatrizz[95][479] = 9'b111111111;
assign micromatrizz[95][480] = 9'b111111111;
assign micromatrizz[95][481] = 9'b111111111;
assign micromatrizz[95][482] = 9'b111111111;
assign micromatrizz[95][483] = 9'b111111111;
assign micromatrizz[95][484] = 9'b111111111;
assign micromatrizz[95][485] = 9'b111111111;
assign micromatrizz[95][486] = 9'b111111111;
assign micromatrizz[95][487] = 9'b111111111;
assign micromatrizz[95][488] = 9'b111111111;
assign micromatrizz[95][489] = 9'b111111111;
assign micromatrizz[95][490] = 9'b111111111;
assign micromatrizz[95][491] = 9'b111111111;
assign micromatrizz[95][492] = 9'b111111111;
assign micromatrizz[95][493] = 9'b111111111;
assign micromatrizz[95][494] = 9'b111111111;
assign micromatrizz[95][495] = 9'b111111111;
assign micromatrizz[95][496] = 9'b111111111;
assign micromatrizz[95][497] = 9'b111111111;
assign micromatrizz[95][498] = 9'b111111111;
assign micromatrizz[95][499] = 9'b111111111;
assign micromatrizz[95][500] = 9'b111111111;
assign micromatrizz[95][501] = 9'b111111111;
assign micromatrizz[95][502] = 9'b111111111;
assign micromatrizz[95][503] = 9'b111111111;
assign micromatrizz[95][504] = 9'b111111111;
assign micromatrizz[95][505] = 9'b111111111;
assign micromatrizz[95][506] = 9'b111111111;
assign micromatrizz[95][507] = 9'b111111111;
assign micromatrizz[95][508] = 9'b111111111;
assign micromatrizz[95][509] = 9'b111111111;
assign micromatrizz[95][510] = 9'b111111111;
assign micromatrizz[95][511] = 9'b111111111;
assign micromatrizz[95][512] = 9'b111111111;
assign micromatrizz[95][513] = 9'b111111111;
assign micromatrizz[95][514] = 9'b111111111;
assign micromatrizz[95][515] = 9'b111111111;
assign micromatrizz[95][516] = 9'b111111111;
assign micromatrizz[95][517] = 9'b111111111;
assign micromatrizz[95][518] = 9'b111111111;
assign micromatrizz[95][519] = 9'b111111111;
assign micromatrizz[95][520] = 9'b111111111;
assign micromatrizz[95][521] = 9'b111111111;
assign micromatrizz[95][522] = 9'b111111111;
assign micromatrizz[95][523] = 9'b111111111;
assign micromatrizz[95][524] = 9'b111111111;
assign micromatrizz[95][525] = 9'b111111111;
assign micromatrizz[95][526] = 9'b111111111;
assign micromatrizz[95][527] = 9'b111111111;
assign micromatrizz[95][528] = 9'b111111111;
assign micromatrizz[95][529] = 9'b111111111;
assign micromatrizz[95][530] = 9'b111111111;
assign micromatrizz[95][531] = 9'b111111111;
assign micromatrizz[95][532] = 9'b111111111;
assign micromatrizz[95][533] = 9'b111111111;
assign micromatrizz[95][534] = 9'b111111111;
assign micromatrizz[95][535] = 9'b111111111;
assign micromatrizz[95][536] = 9'b111111111;
assign micromatrizz[95][537] = 9'b111111111;
assign micromatrizz[95][538] = 9'b111111111;
assign micromatrizz[95][539] = 9'b111111111;
assign micromatrizz[95][540] = 9'b111111111;
assign micromatrizz[95][541] = 9'b111111111;
assign micromatrizz[95][542] = 9'b111111111;
assign micromatrizz[95][543] = 9'b111111111;
assign micromatrizz[95][544] = 9'b111111111;
assign micromatrizz[95][545] = 9'b111111111;
assign micromatrizz[95][546] = 9'b111111111;
assign micromatrizz[95][547] = 9'b111111111;
assign micromatrizz[95][548] = 9'b111111111;
assign micromatrizz[95][549] = 9'b111111111;
assign micromatrizz[95][550] = 9'b111111111;
assign micromatrizz[95][551] = 9'b111111111;
assign micromatrizz[95][552] = 9'b111111111;
assign micromatrizz[95][553] = 9'b111111111;
assign micromatrizz[95][554] = 9'b111111111;
assign micromatrizz[95][555] = 9'b111111111;
assign micromatrizz[95][556] = 9'b111111111;
assign micromatrizz[95][557] = 9'b111111111;
assign micromatrizz[95][558] = 9'b111111111;
assign micromatrizz[95][559] = 9'b111111111;
assign micromatrizz[95][560] = 9'b111111111;
assign micromatrizz[95][561] = 9'b111111111;
assign micromatrizz[95][562] = 9'b111111111;
assign micromatrizz[95][563] = 9'b111111111;
assign micromatrizz[95][564] = 9'b111111111;
assign micromatrizz[95][565] = 9'b111111111;
assign micromatrizz[95][566] = 9'b111111111;
assign micromatrizz[95][567] = 9'b111111111;
assign micromatrizz[95][568] = 9'b111111111;
assign micromatrizz[95][569] = 9'b111111111;
assign micromatrizz[95][570] = 9'b111111111;
assign micromatrizz[95][571] = 9'b111111111;
assign micromatrizz[95][572] = 9'b111111111;
assign micromatrizz[95][573] = 9'b111111111;
assign micromatrizz[95][574] = 9'b111111111;
assign micromatrizz[95][575] = 9'b111111111;
assign micromatrizz[95][576] = 9'b111111111;
assign micromatrizz[95][577] = 9'b111111111;
assign micromatrizz[95][578] = 9'b111111111;
assign micromatrizz[95][579] = 9'b111111111;
assign micromatrizz[95][580] = 9'b111111111;
assign micromatrizz[95][581] = 9'b111111111;
assign micromatrizz[95][582] = 9'b111111111;
assign micromatrizz[95][583] = 9'b111111111;
assign micromatrizz[95][584] = 9'b111111111;
assign micromatrizz[95][585] = 9'b111111111;
assign micromatrizz[95][586] = 9'b111111111;
assign micromatrizz[95][587] = 9'b111111111;
assign micromatrizz[95][588] = 9'b111111111;
assign micromatrizz[95][589] = 9'b111111111;
assign micromatrizz[95][590] = 9'b111111111;
assign micromatrizz[95][591] = 9'b111111111;
assign micromatrizz[95][592] = 9'b111111111;
assign micromatrizz[95][593] = 9'b111111111;
assign micromatrizz[95][594] = 9'b111111111;
assign micromatrizz[95][595] = 9'b111111111;
assign micromatrizz[95][596] = 9'b111111111;
assign micromatrizz[95][597] = 9'b111111111;
assign micromatrizz[95][598] = 9'b111111111;
assign micromatrizz[95][599] = 9'b111111111;
assign micromatrizz[95][600] = 9'b111111111;
assign micromatrizz[95][601] = 9'b111111111;
assign micromatrizz[95][602] = 9'b111111111;
assign micromatrizz[95][603] = 9'b111111111;
assign micromatrizz[95][604] = 9'b111111111;
assign micromatrizz[95][605] = 9'b111111111;
assign micromatrizz[95][606] = 9'b111111111;
assign micromatrizz[95][607] = 9'b111111111;
assign micromatrizz[95][608] = 9'b111111111;
assign micromatrizz[95][609] = 9'b111111111;
assign micromatrizz[95][610] = 9'b111111111;
assign micromatrizz[95][611] = 9'b111111111;
assign micromatrizz[95][612] = 9'b111111111;
assign micromatrizz[95][613] = 9'b111111111;
assign micromatrizz[95][614] = 9'b111111111;
assign micromatrizz[95][615] = 9'b111111111;
assign micromatrizz[95][616] = 9'b111111111;
assign micromatrizz[95][617] = 9'b111111111;
assign micromatrizz[95][618] = 9'b111111111;
assign micromatrizz[95][619] = 9'b111111111;
assign micromatrizz[95][620] = 9'b111111111;
assign micromatrizz[95][621] = 9'b111111111;
assign micromatrizz[95][622] = 9'b111111111;
assign micromatrizz[95][623] = 9'b111111111;
assign micromatrizz[95][624] = 9'b111111111;
assign micromatrizz[95][625] = 9'b111111111;
assign micromatrizz[95][626] = 9'b111111111;
assign micromatrizz[95][627] = 9'b111111111;
assign micromatrizz[95][628] = 9'b111111111;
assign micromatrizz[95][629] = 9'b111111111;
assign micromatrizz[95][630] = 9'b111111111;
assign micromatrizz[95][631] = 9'b111111111;
assign micromatrizz[95][632] = 9'b111111111;
assign micromatrizz[95][633] = 9'b111111111;
assign micromatrizz[95][634] = 9'b111111111;
assign micromatrizz[95][635] = 9'b111111111;
assign micromatrizz[95][636] = 9'b111111111;
assign micromatrizz[95][637] = 9'b111111111;
assign micromatrizz[95][638] = 9'b111111111;
assign micromatrizz[95][639] = 9'b111111111;
assign micromatrizz[96][0] = 9'b111111111;
assign micromatrizz[96][1] = 9'b111111111;
assign micromatrizz[96][2] = 9'b111111111;
assign micromatrizz[96][3] = 9'b111111111;
assign micromatrizz[96][4] = 9'b111111111;
assign micromatrizz[96][5] = 9'b111111111;
assign micromatrizz[96][6] = 9'b111111111;
assign micromatrizz[96][7] = 9'b111111111;
assign micromatrizz[96][8] = 9'b111111111;
assign micromatrizz[96][9] = 9'b111111111;
assign micromatrizz[96][10] = 9'b111111111;
assign micromatrizz[96][11] = 9'b111111111;
assign micromatrizz[96][12] = 9'b111111111;
assign micromatrizz[96][13] = 9'b111111111;
assign micromatrizz[96][14] = 9'b111111111;
assign micromatrizz[96][15] = 9'b111111111;
assign micromatrizz[96][16] = 9'b111111111;
assign micromatrizz[96][17] = 9'b111111111;
assign micromatrizz[96][18] = 9'b111111111;
assign micromatrizz[96][19] = 9'b111111111;
assign micromatrizz[96][20] = 9'b111111111;
assign micromatrizz[96][21] = 9'b111111111;
assign micromatrizz[96][22] = 9'b111111111;
assign micromatrizz[96][23] = 9'b111111111;
assign micromatrizz[96][24] = 9'b111111111;
assign micromatrizz[96][25] = 9'b111111111;
assign micromatrizz[96][26] = 9'b111111111;
assign micromatrizz[96][27] = 9'b111111111;
assign micromatrizz[96][28] = 9'b111111111;
assign micromatrizz[96][29] = 9'b111111111;
assign micromatrizz[96][30] = 9'b111111111;
assign micromatrizz[96][31] = 9'b111111111;
assign micromatrizz[96][32] = 9'b111111111;
assign micromatrizz[96][33] = 9'b111111111;
assign micromatrizz[96][34] = 9'b111111111;
assign micromatrizz[96][35] = 9'b111111111;
assign micromatrizz[96][36] = 9'b111111111;
assign micromatrizz[96][37] = 9'b111111111;
assign micromatrizz[96][38] = 9'b111111111;
assign micromatrizz[96][39] = 9'b111111111;
assign micromatrizz[96][40] = 9'b111111111;
assign micromatrizz[96][41] = 9'b111111111;
assign micromatrizz[96][42] = 9'b111111111;
assign micromatrizz[96][43] = 9'b111111111;
assign micromatrizz[96][44] = 9'b111111111;
assign micromatrizz[96][45] = 9'b111111111;
assign micromatrizz[96][46] = 9'b111111111;
assign micromatrizz[96][47] = 9'b111111111;
assign micromatrizz[96][48] = 9'b111111111;
assign micromatrizz[96][49] = 9'b111111111;
assign micromatrizz[96][50] = 9'b111111111;
assign micromatrizz[96][51] = 9'b111111111;
assign micromatrizz[96][52] = 9'b111111111;
assign micromatrizz[96][53] = 9'b111111111;
assign micromatrizz[96][54] = 9'b111111111;
assign micromatrizz[96][55] = 9'b111111111;
assign micromatrizz[96][56] = 9'b111111111;
assign micromatrizz[96][57] = 9'b111111111;
assign micromatrizz[96][58] = 9'b111111111;
assign micromatrizz[96][59] = 9'b111111111;
assign micromatrizz[96][60] = 9'b111111111;
assign micromatrizz[96][61] = 9'b111111111;
assign micromatrizz[96][62] = 9'b111111111;
assign micromatrizz[96][63] = 9'b111111111;
assign micromatrizz[96][64] = 9'b111111111;
assign micromatrizz[96][65] = 9'b111111111;
assign micromatrizz[96][66] = 9'b111111111;
assign micromatrizz[96][67] = 9'b111111111;
assign micromatrizz[96][68] = 9'b111111111;
assign micromatrizz[96][69] = 9'b111111111;
assign micromatrizz[96][70] = 9'b111111111;
assign micromatrizz[96][71] = 9'b111111111;
assign micromatrizz[96][72] = 9'b111111111;
assign micromatrizz[96][73] = 9'b111111111;
assign micromatrizz[96][74] = 9'b111111111;
assign micromatrizz[96][75] = 9'b111111111;
assign micromatrizz[96][76] = 9'b111111111;
assign micromatrizz[96][77] = 9'b111111111;
assign micromatrizz[96][78] = 9'b111111111;
assign micromatrizz[96][79] = 9'b111111111;
assign micromatrizz[96][80] = 9'b111111111;
assign micromatrizz[96][81] = 9'b111111111;
assign micromatrizz[96][82] = 9'b111111111;
assign micromatrizz[96][83] = 9'b111111111;
assign micromatrizz[96][84] = 9'b111111111;
assign micromatrizz[96][85] = 9'b111111111;
assign micromatrizz[96][86] = 9'b111111111;
assign micromatrizz[96][87] = 9'b111111111;
assign micromatrizz[96][88] = 9'b111111111;
assign micromatrizz[96][89] = 9'b111111111;
assign micromatrizz[96][90] = 9'b111111111;
assign micromatrizz[96][91] = 9'b111111111;
assign micromatrizz[96][92] = 9'b111111111;
assign micromatrizz[96][93] = 9'b111111111;
assign micromatrizz[96][94] = 9'b111111111;
assign micromatrizz[96][95] = 9'b111111111;
assign micromatrizz[96][96] = 9'b111111111;
assign micromatrizz[96][97] = 9'b111111111;
assign micromatrizz[96][98] = 9'b111111111;
assign micromatrizz[96][99] = 9'b111111111;
assign micromatrizz[96][100] = 9'b111111111;
assign micromatrizz[96][101] = 9'b111111111;
assign micromatrizz[96][102] = 9'b111111111;
assign micromatrizz[96][103] = 9'b111111111;
assign micromatrizz[96][104] = 9'b111111111;
assign micromatrizz[96][105] = 9'b111111111;
assign micromatrizz[96][106] = 9'b111111111;
assign micromatrizz[96][107] = 9'b111111111;
assign micromatrizz[96][108] = 9'b111111111;
assign micromatrizz[96][109] = 9'b111111111;
assign micromatrizz[96][110] = 9'b111111111;
assign micromatrizz[96][111] = 9'b111111111;
assign micromatrizz[96][112] = 9'b111111111;
assign micromatrizz[96][113] = 9'b111111111;
assign micromatrizz[96][114] = 9'b111111111;
assign micromatrizz[96][115] = 9'b111111111;
assign micromatrizz[96][116] = 9'b111111111;
assign micromatrizz[96][117] = 9'b111111111;
assign micromatrizz[96][118] = 9'b111111111;
assign micromatrizz[96][119] = 9'b111111111;
assign micromatrizz[96][120] = 9'b111111111;
assign micromatrizz[96][121] = 9'b111111111;
assign micromatrizz[96][122] = 9'b111111111;
assign micromatrizz[96][123] = 9'b111111111;
assign micromatrizz[96][124] = 9'b111111111;
assign micromatrizz[96][125] = 9'b111111111;
assign micromatrizz[96][126] = 9'b111111111;
assign micromatrizz[96][127] = 9'b111111111;
assign micromatrizz[96][128] = 9'b111111111;
assign micromatrizz[96][129] = 9'b111111111;
assign micromatrizz[96][130] = 9'b111111111;
assign micromatrizz[96][131] = 9'b111111111;
assign micromatrizz[96][132] = 9'b111111111;
assign micromatrizz[96][133] = 9'b111111111;
assign micromatrizz[96][134] = 9'b111111111;
assign micromatrizz[96][135] = 9'b111111111;
assign micromatrizz[96][136] = 9'b111111111;
assign micromatrizz[96][137] = 9'b111111111;
assign micromatrizz[96][138] = 9'b111111111;
assign micromatrizz[96][139] = 9'b111111111;
assign micromatrizz[96][140] = 9'b111111111;
assign micromatrizz[96][141] = 9'b111111111;
assign micromatrizz[96][142] = 9'b111111111;
assign micromatrizz[96][143] = 9'b111111111;
assign micromatrizz[96][144] = 9'b111111111;
assign micromatrizz[96][145] = 9'b111111111;
assign micromatrizz[96][146] = 9'b111111111;
assign micromatrizz[96][147] = 9'b111111111;
assign micromatrizz[96][148] = 9'b111111111;
assign micromatrizz[96][149] = 9'b111111111;
assign micromatrizz[96][150] = 9'b111111111;
assign micromatrizz[96][151] = 9'b111111111;
assign micromatrizz[96][152] = 9'b111111111;
assign micromatrizz[96][153] = 9'b111111111;
assign micromatrizz[96][154] = 9'b111111111;
assign micromatrizz[96][155] = 9'b111111111;
assign micromatrizz[96][156] = 9'b111111111;
assign micromatrizz[96][157] = 9'b111111111;
assign micromatrizz[96][158] = 9'b111111111;
assign micromatrizz[96][159] = 9'b111111111;
assign micromatrizz[96][160] = 9'b111111111;
assign micromatrizz[96][161] = 9'b111111111;
assign micromatrizz[96][162] = 9'b111111111;
assign micromatrizz[96][163] = 9'b111111111;
assign micromatrizz[96][164] = 9'b111111111;
assign micromatrizz[96][165] = 9'b111111111;
assign micromatrizz[96][166] = 9'b111111111;
assign micromatrizz[96][167] = 9'b111111111;
assign micromatrizz[96][168] = 9'b111111111;
assign micromatrizz[96][169] = 9'b111111111;
assign micromatrizz[96][170] = 9'b111111111;
assign micromatrizz[96][171] = 9'b111111111;
assign micromatrizz[96][172] = 9'b111111111;
assign micromatrizz[96][173] = 9'b111111111;
assign micromatrizz[96][174] = 9'b111111111;
assign micromatrizz[96][175] = 9'b111111111;
assign micromatrizz[96][176] = 9'b111111111;
assign micromatrizz[96][177] = 9'b111111111;
assign micromatrizz[96][178] = 9'b111111111;
assign micromatrizz[96][179] = 9'b111111111;
assign micromatrizz[96][180] = 9'b111111111;
assign micromatrizz[96][181] = 9'b111111111;
assign micromatrizz[96][182] = 9'b111111111;
assign micromatrizz[96][183] = 9'b111111111;
assign micromatrizz[96][184] = 9'b111111111;
assign micromatrizz[96][185] = 9'b111111111;
assign micromatrizz[96][186] = 9'b111111111;
assign micromatrizz[96][187] = 9'b111111111;
assign micromatrizz[96][188] = 9'b111111111;
assign micromatrizz[96][189] = 9'b111111111;
assign micromatrizz[96][190] = 9'b111111111;
assign micromatrizz[96][191] = 9'b111111111;
assign micromatrizz[96][192] = 9'b111111111;
assign micromatrizz[96][193] = 9'b111111111;
assign micromatrizz[96][194] = 9'b111111111;
assign micromatrizz[96][195] = 9'b111111111;
assign micromatrizz[96][196] = 9'b111111111;
assign micromatrizz[96][197] = 9'b111111111;
assign micromatrizz[96][198] = 9'b111111111;
assign micromatrizz[96][199] = 9'b111111111;
assign micromatrizz[96][200] = 9'b111111111;
assign micromatrizz[96][201] = 9'b111111111;
assign micromatrizz[96][202] = 9'b111111111;
assign micromatrizz[96][203] = 9'b111111111;
assign micromatrizz[96][204] = 9'b111111111;
assign micromatrizz[96][205] = 9'b111111111;
assign micromatrizz[96][206] = 9'b111111111;
assign micromatrizz[96][207] = 9'b111111111;
assign micromatrizz[96][208] = 9'b111111111;
assign micromatrizz[96][209] = 9'b111111111;
assign micromatrizz[96][210] = 9'b111111111;
assign micromatrizz[96][211] = 9'b111111111;
assign micromatrizz[96][212] = 9'b111111111;
assign micromatrizz[96][213] = 9'b111111111;
assign micromatrizz[96][214] = 9'b111111111;
assign micromatrizz[96][215] = 9'b111111111;
assign micromatrizz[96][216] = 9'b111111111;
assign micromatrizz[96][217] = 9'b111111111;
assign micromatrizz[96][218] = 9'b111111111;
assign micromatrizz[96][219] = 9'b111111111;
assign micromatrizz[96][220] = 9'b111111111;
assign micromatrizz[96][221] = 9'b111111111;
assign micromatrizz[96][222] = 9'b111111111;
assign micromatrizz[96][223] = 9'b111111111;
assign micromatrizz[96][224] = 9'b111111111;
assign micromatrizz[96][225] = 9'b111111111;
assign micromatrizz[96][226] = 9'b111111111;
assign micromatrizz[96][227] = 9'b111111111;
assign micromatrizz[96][228] = 9'b111111111;
assign micromatrizz[96][229] = 9'b111111111;
assign micromatrizz[96][230] = 9'b111111111;
assign micromatrizz[96][231] = 9'b111111111;
assign micromatrizz[96][232] = 9'b111111111;
assign micromatrizz[96][233] = 9'b111111111;
assign micromatrizz[96][234] = 9'b111111111;
assign micromatrizz[96][235] = 9'b111111111;
assign micromatrizz[96][236] = 9'b111111111;
assign micromatrizz[96][237] = 9'b111111111;
assign micromatrizz[96][238] = 9'b111111111;
assign micromatrizz[96][239] = 9'b111111111;
assign micromatrizz[96][240] = 9'b111111111;
assign micromatrizz[96][241] = 9'b111111111;
assign micromatrizz[96][242] = 9'b111111111;
assign micromatrizz[96][243] = 9'b111111111;
assign micromatrizz[96][244] = 9'b111111111;
assign micromatrizz[96][245] = 9'b111111111;
assign micromatrizz[96][246] = 9'b111111111;
assign micromatrizz[96][247] = 9'b111111111;
assign micromatrizz[96][248] = 9'b111111111;
assign micromatrizz[96][249] = 9'b111111111;
assign micromatrizz[96][250] = 9'b111111111;
assign micromatrizz[96][251] = 9'b111111111;
assign micromatrizz[96][252] = 9'b111111111;
assign micromatrizz[96][253] = 9'b111111111;
assign micromatrizz[96][254] = 9'b111111111;
assign micromatrizz[96][255] = 9'b111111111;
assign micromatrizz[96][256] = 9'b111111111;
assign micromatrizz[96][257] = 9'b111111111;
assign micromatrizz[96][258] = 9'b111111111;
assign micromatrizz[96][259] = 9'b111111111;
assign micromatrizz[96][260] = 9'b111111111;
assign micromatrizz[96][261] = 9'b111111111;
assign micromatrizz[96][262] = 9'b111111111;
assign micromatrizz[96][263] = 9'b111111111;
assign micromatrizz[96][264] = 9'b111111111;
assign micromatrizz[96][265] = 9'b111111111;
assign micromatrizz[96][266] = 9'b111111111;
assign micromatrizz[96][267] = 9'b111111111;
assign micromatrizz[96][268] = 9'b111111111;
assign micromatrizz[96][269] = 9'b111111111;
assign micromatrizz[96][270] = 9'b111111111;
assign micromatrizz[96][271] = 9'b111111111;
assign micromatrizz[96][272] = 9'b111111111;
assign micromatrizz[96][273] = 9'b111111111;
assign micromatrizz[96][274] = 9'b111111111;
assign micromatrizz[96][275] = 9'b111111111;
assign micromatrizz[96][276] = 9'b111111111;
assign micromatrizz[96][277] = 9'b111111111;
assign micromatrizz[96][278] = 9'b111111111;
assign micromatrizz[96][279] = 9'b111111111;
assign micromatrizz[96][280] = 9'b111111111;
assign micromatrizz[96][281] = 9'b111111111;
assign micromatrizz[96][282] = 9'b111111111;
assign micromatrizz[96][283] = 9'b111111111;
assign micromatrizz[96][284] = 9'b111111111;
assign micromatrizz[96][285] = 9'b111111111;
assign micromatrizz[96][286] = 9'b111111111;
assign micromatrizz[96][287] = 9'b111111111;
assign micromatrizz[96][288] = 9'b111111111;
assign micromatrizz[96][289] = 9'b111111111;
assign micromatrizz[96][290] = 9'b111111111;
assign micromatrizz[96][291] = 9'b111111111;
assign micromatrizz[96][292] = 9'b111111111;
assign micromatrizz[96][293] = 9'b111111111;
assign micromatrizz[96][294] = 9'b111111111;
assign micromatrizz[96][295] = 9'b111111111;
assign micromatrizz[96][296] = 9'b111111111;
assign micromatrizz[96][297] = 9'b111111111;
assign micromatrizz[96][298] = 9'b111111111;
assign micromatrizz[96][299] = 9'b111111111;
assign micromatrizz[96][300] = 9'b111111111;
assign micromatrizz[96][301] = 9'b111111111;
assign micromatrizz[96][302] = 9'b111111111;
assign micromatrizz[96][303] = 9'b111111111;
assign micromatrizz[96][304] = 9'b111111111;
assign micromatrizz[96][305] = 9'b111111111;
assign micromatrizz[96][306] = 9'b111111111;
assign micromatrizz[96][307] = 9'b111111111;
assign micromatrizz[96][308] = 9'b111111111;
assign micromatrizz[96][309] = 9'b111111111;
assign micromatrizz[96][310] = 9'b111111111;
assign micromatrizz[96][311] = 9'b111111111;
assign micromatrizz[96][312] = 9'b111111111;
assign micromatrizz[96][313] = 9'b111111111;
assign micromatrizz[96][314] = 9'b111111111;
assign micromatrizz[96][315] = 9'b111111111;
assign micromatrizz[96][316] = 9'b111111111;
assign micromatrizz[96][317] = 9'b111111111;
assign micromatrizz[96][318] = 9'b111111111;
assign micromatrizz[96][319] = 9'b111111111;
assign micromatrizz[96][320] = 9'b111111111;
assign micromatrizz[96][321] = 9'b111111111;
assign micromatrizz[96][322] = 9'b111111111;
assign micromatrizz[96][323] = 9'b111111111;
assign micromatrizz[96][324] = 9'b111111111;
assign micromatrizz[96][325] = 9'b111111111;
assign micromatrizz[96][326] = 9'b111111111;
assign micromatrizz[96][327] = 9'b111111111;
assign micromatrizz[96][328] = 9'b111111111;
assign micromatrizz[96][329] = 9'b111111111;
assign micromatrizz[96][330] = 9'b111111111;
assign micromatrizz[96][331] = 9'b111111111;
assign micromatrizz[96][332] = 9'b111111111;
assign micromatrizz[96][333] = 9'b111111111;
assign micromatrizz[96][334] = 9'b111111111;
assign micromatrizz[96][335] = 9'b111111111;
assign micromatrizz[96][336] = 9'b111111111;
assign micromatrizz[96][337] = 9'b111111111;
assign micromatrizz[96][338] = 9'b111111111;
assign micromatrizz[96][339] = 9'b111111111;
assign micromatrizz[96][340] = 9'b111111111;
assign micromatrizz[96][341] = 9'b111111111;
assign micromatrizz[96][342] = 9'b111111111;
assign micromatrizz[96][343] = 9'b111111111;
assign micromatrizz[96][344] = 9'b111111111;
assign micromatrizz[96][345] = 9'b111111111;
assign micromatrizz[96][346] = 9'b111111111;
assign micromatrizz[96][347] = 9'b111111111;
assign micromatrizz[96][348] = 9'b111111111;
assign micromatrizz[96][349] = 9'b111111111;
assign micromatrizz[96][350] = 9'b111111111;
assign micromatrizz[96][351] = 9'b111111111;
assign micromatrizz[96][352] = 9'b111111111;
assign micromatrizz[96][353] = 9'b111111111;
assign micromatrizz[96][354] = 9'b111111111;
assign micromatrizz[96][355] = 9'b111111111;
assign micromatrizz[96][356] = 9'b111111111;
assign micromatrizz[96][357] = 9'b111111111;
assign micromatrizz[96][358] = 9'b111111111;
assign micromatrizz[96][359] = 9'b111111111;
assign micromatrizz[96][360] = 9'b111111111;
assign micromatrizz[96][361] = 9'b111111111;
assign micromatrizz[96][362] = 9'b111111111;
assign micromatrizz[96][363] = 9'b111111111;
assign micromatrizz[96][364] = 9'b111111111;
assign micromatrizz[96][365] = 9'b111111111;
assign micromatrizz[96][366] = 9'b111111111;
assign micromatrizz[96][367] = 9'b111111111;
assign micromatrizz[96][368] = 9'b111111111;
assign micromatrizz[96][369] = 9'b111111111;
assign micromatrizz[96][370] = 9'b111111111;
assign micromatrizz[96][371] = 9'b111111111;
assign micromatrizz[96][372] = 9'b111111111;
assign micromatrizz[96][373] = 9'b111111111;
assign micromatrizz[96][374] = 9'b111111111;
assign micromatrizz[96][375] = 9'b111111111;
assign micromatrizz[96][376] = 9'b111111111;
assign micromatrizz[96][377] = 9'b111111111;
assign micromatrizz[96][378] = 9'b111111111;
assign micromatrizz[96][379] = 9'b111111111;
assign micromatrizz[96][380] = 9'b111111111;
assign micromatrizz[96][381] = 9'b111111111;
assign micromatrizz[96][382] = 9'b111111111;
assign micromatrizz[96][383] = 9'b111111111;
assign micromatrizz[96][384] = 9'b111111111;
assign micromatrizz[96][385] = 9'b111111111;
assign micromatrizz[96][386] = 9'b111111111;
assign micromatrizz[96][387] = 9'b111111111;
assign micromatrizz[96][388] = 9'b111111111;
assign micromatrizz[96][389] = 9'b111111111;
assign micromatrizz[96][390] = 9'b111111111;
assign micromatrizz[96][391] = 9'b111111111;
assign micromatrizz[96][392] = 9'b111111111;
assign micromatrizz[96][393] = 9'b111111111;
assign micromatrizz[96][394] = 9'b111111111;
assign micromatrizz[96][395] = 9'b111111111;
assign micromatrizz[96][396] = 9'b111111111;
assign micromatrizz[96][397] = 9'b111111111;
assign micromatrizz[96][398] = 9'b111111111;
assign micromatrizz[96][399] = 9'b111111111;
assign micromatrizz[96][400] = 9'b111111111;
assign micromatrizz[96][401] = 9'b111111111;
assign micromatrizz[96][402] = 9'b111111111;
assign micromatrizz[96][403] = 9'b111111111;
assign micromatrizz[96][404] = 9'b111111111;
assign micromatrizz[96][405] = 9'b111111111;
assign micromatrizz[96][406] = 9'b111111111;
assign micromatrizz[96][407] = 9'b111111111;
assign micromatrizz[96][408] = 9'b111111111;
assign micromatrizz[96][409] = 9'b111111111;
assign micromatrizz[96][410] = 9'b111111111;
assign micromatrizz[96][411] = 9'b111111111;
assign micromatrizz[96][412] = 9'b111111111;
assign micromatrizz[96][413] = 9'b111111111;
assign micromatrizz[96][414] = 9'b111111111;
assign micromatrizz[96][415] = 9'b111111111;
assign micromatrizz[96][416] = 9'b111111111;
assign micromatrizz[96][417] = 9'b111111111;
assign micromatrizz[96][418] = 9'b111111111;
assign micromatrizz[96][419] = 9'b111111111;
assign micromatrizz[96][420] = 9'b111111111;
assign micromatrizz[96][421] = 9'b111111111;
assign micromatrizz[96][422] = 9'b111111111;
assign micromatrizz[96][423] = 9'b111111111;
assign micromatrizz[96][424] = 9'b111111111;
assign micromatrizz[96][425] = 9'b111111111;
assign micromatrizz[96][426] = 9'b111111111;
assign micromatrizz[96][427] = 9'b111111111;
assign micromatrizz[96][428] = 9'b111111111;
assign micromatrizz[96][429] = 9'b111111111;
assign micromatrizz[96][430] = 9'b111111111;
assign micromatrizz[96][431] = 9'b111111111;
assign micromatrizz[96][432] = 9'b111111111;
assign micromatrizz[96][433] = 9'b111111111;
assign micromatrizz[96][434] = 9'b111111111;
assign micromatrizz[96][435] = 9'b111111111;
assign micromatrizz[96][436] = 9'b111111111;
assign micromatrizz[96][437] = 9'b111111111;
assign micromatrizz[96][438] = 9'b111111111;
assign micromatrizz[96][439] = 9'b111111111;
assign micromatrizz[96][440] = 9'b111111111;
assign micromatrizz[96][441] = 9'b111111111;
assign micromatrizz[96][442] = 9'b111111111;
assign micromatrizz[96][443] = 9'b111111111;
assign micromatrizz[96][444] = 9'b111111111;
assign micromatrizz[96][445] = 9'b111111111;
assign micromatrizz[96][446] = 9'b111111111;
assign micromatrizz[96][447] = 9'b111111111;
assign micromatrizz[96][448] = 9'b111111111;
assign micromatrizz[96][449] = 9'b111111111;
assign micromatrizz[96][450] = 9'b111111111;
assign micromatrizz[96][451] = 9'b111111111;
assign micromatrizz[96][452] = 9'b111111111;
assign micromatrizz[96][453] = 9'b111111111;
assign micromatrizz[96][454] = 9'b111111111;
assign micromatrizz[96][455] = 9'b111111111;
assign micromatrizz[96][456] = 9'b111111111;
assign micromatrizz[96][457] = 9'b111111111;
assign micromatrizz[96][458] = 9'b111111111;
assign micromatrizz[96][459] = 9'b111111111;
assign micromatrizz[96][460] = 9'b111111111;
assign micromatrizz[96][461] = 9'b111111111;
assign micromatrizz[96][462] = 9'b111111111;
assign micromatrizz[96][463] = 9'b111111111;
assign micromatrizz[96][464] = 9'b111111111;
assign micromatrizz[96][465] = 9'b111111111;
assign micromatrizz[96][466] = 9'b111111111;
assign micromatrizz[96][467] = 9'b111111111;
assign micromatrizz[96][468] = 9'b111111111;
assign micromatrizz[96][469] = 9'b111111111;
assign micromatrizz[96][470] = 9'b111111111;
assign micromatrizz[96][471] = 9'b111111111;
assign micromatrizz[96][472] = 9'b111111111;
assign micromatrizz[96][473] = 9'b111111111;
assign micromatrizz[96][474] = 9'b111111111;
assign micromatrizz[96][475] = 9'b111111111;
assign micromatrizz[96][476] = 9'b111111111;
assign micromatrizz[96][477] = 9'b111111111;
assign micromatrizz[96][478] = 9'b111111111;
assign micromatrizz[96][479] = 9'b111111111;
assign micromatrizz[96][480] = 9'b111111111;
assign micromatrizz[96][481] = 9'b111111111;
assign micromatrizz[96][482] = 9'b111111111;
assign micromatrizz[96][483] = 9'b111111111;
assign micromatrizz[96][484] = 9'b111111111;
assign micromatrizz[96][485] = 9'b111111111;
assign micromatrizz[96][486] = 9'b111111111;
assign micromatrizz[96][487] = 9'b111111111;
assign micromatrizz[96][488] = 9'b111111111;
assign micromatrizz[96][489] = 9'b111111111;
assign micromatrizz[96][490] = 9'b111111111;
assign micromatrizz[96][491] = 9'b111111111;
assign micromatrizz[96][492] = 9'b111111111;
assign micromatrizz[96][493] = 9'b111111111;
assign micromatrizz[96][494] = 9'b111111111;
assign micromatrizz[96][495] = 9'b111111111;
assign micromatrizz[96][496] = 9'b111111111;
assign micromatrizz[96][497] = 9'b111111111;
assign micromatrizz[96][498] = 9'b111111111;
assign micromatrizz[96][499] = 9'b111111111;
assign micromatrizz[96][500] = 9'b111111111;
assign micromatrizz[96][501] = 9'b111111111;
assign micromatrizz[96][502] = 9'b111111111;
assign micromatrizz[96][503] = 9'b111111111;
assign micromatrizz[96][504] = 9'b111111111;
assign micromatrizz[96][505] = 9'b111111111;
assign micromatrizz[96][506] = 9'b111111111;
assign micromatrizz[96][507] = 9'b111111111;
assign micromatrizz[96][508] = 9'b111111111;
assign micromatrizz[96][509] = 9'b111111111;
assign micromatrizz[96][510] = 9'b111111111;
assign micromatrizz[96][511] = 9'b111111111;
assign micromatrizz[96][512] = 9'b111111111;
assign micromatrizz[96][513] = 9'b111111111;
assign micromatrizz[96][514] = 9'b111111111;
assign micromatrizz[96][515] = 9'b111111111;
assign micromatrizz[96][516] = 9'b111111111;
assign micromatrizz[96][517] = 9'b111111111;
assign micromatrizz[96][518] = 9'b111111111;
assign micromatrizz[96][519] = 9'b111111111;
assign micromatrizz[96][520] = 9'b111111111;
assign micromatrizz[96][521] = 9'b111111111;
assign micromatrizz[96][522] = 9'b111111111;
assign micromatrizz[96][523] = 9'b111111111;
assign micromatrizz[96][524] = 9'b111111111;
assign micromatrizz[96][525] = 9'b111111111;
assign micromatrizz[96][526] = 9'b111111111;
assign micromatrizz[96][527] = 9'b111111111;
assign micromatrizz[96][528] = 9'b111111111;
assign micromatrizz[96][529] = 9'b111111111;
assign micromatrizz[96][530] = 9'b111111111;
assign micromatrizz[96][531] = 9'b111111111;
assign micromatrizz[96][532] = 9'b111111111;
assign micromatrizz[96][533] = 9'b111111111;
assign micromatrizz[96][534] = 9'b111111111;
assign micromatrizz[96][535] = 9'b111111111;
assign micromatrizz[96][536] = 9'b111111111;
assign micromatrizz[96][537] = 9'b111111111;
assign micromatrizz[96][538] = 9'b111111111;
assign micromatrizz[96][539] = 9'b111111111;
assign micromatrizz[96][540] = 9'b111111111;
assign micromatrizz[96][541] = 9'b111111111;
assign micromatrizz[96][542] = 9'b111111111;
assign micromatrizz[96][543] = 9'b111111111;
assign micromatrizz[96][544] = 9'b111111111;
assign micromatrizz[96][545] = 9'b111111111;
assign micromatrizz[96][546] = 9'b111111111;
assign micromatrizz[96][547] = 9'b111111111;
assign micromatrizz[96][548] = 9'b111111111;
assign micromatrizz[96][549] = 9'b111111111;
assign micromatrizz[96][550] = 9'b111111111;
assign micromatrizz[96][551] = 9'b111111111;
assign micromatrizz[96][552] = 9'b111111111;
assign micromatrizz[96][553] = 9'b111111111;
assign micromatrizz[96][554] = 9'b111111111;
assign micromatrizz[96][555] = 9'b111111111;
assign micromatrizz[96][556] = 9'b111111111;
assign micromatrizz[96][557] = 9'b111111111;
assign micromatrizz[96][558] = 9'b111111111;
assign micromatrizz[96][559] = 9'b111111111;
assign micromatrizz[96][560] = 9'b111111111;
assign micromatrizz[96][561] = 9'b111111111;
assign micromatrizz[96][562] = 9'b111111111;
assign micromatrizz[96][563] = 9'b111111111;
assign micromatrizz[96][564] = 9'b111111111;
assign micromatrizz[96][565] = 9'b111111111;
assign micromatrizz[96][566] = 9'b111111111;
assign micromatrizz[96][567] = 9'b111111111;
assign micromatrizz[96][568] = 9'b111111111;
assign micromatrizz[96][569] = 9'b111111111;
assign micromatrizz[96][570] = 9'b111111111;
assign micromatrizz[96][571] = 9'b111111111;
assign micromatrizz[96][572] = 9'b111111111;
assign micromatrizz[96][573] = 9'b111111111;
assign micromatrizz[96][574] = 9'b111111111;
assign micromatrizz[96][575] = 9'b111111111;
assign micromatrizz[96][576] = 9'b111111111;
assign micromatrizz[96][577] = 9'b111111111;
assign micromatrizz[96][578] = 9'b111111111;
assign micromatrizz[96][579] = 9'b111111111;
assign micromatrizz[96][580] = 9'b111111111;
assign micromatrizz[96][581] = 9'b111111111;
assign micromatrizz[96][582] = 9'b111111111;
assign micromatrizz[96][583] = 9'b111111111;
assign micromatrizz[96][584] = 9'b111111111;
assign micromatrizz[96][585] = 9'b111111111;
assign micromatrizz[96][586] = 9'b111111111;
assign micromatrizz[96][587] = 9'b111111111;
assign micromatrizz[96][588] = 9'b111111111;
assign micromatrizz[96][589] = 9'b111111111;
assign micromatrizz[96][590] = 9'b111111111;
assign micromatrizz[96][591] = 9'b111111111;
assign micromatrizz[96][592] = 9'b111111111;
assign micromatrizz[96][593] = 9'b111111111;
assign micromatrizz[96][594] = 9'b111111111;
assign micromatrizz[96][595] = 9'b111111111;
assign micromatrizz[96][596] = 9'b111111111;
assign micromatrizz[96][597] = 9'b111111111;
assign micromatrizz[96][598] = 9'b111111111;
assign micromatrizz[96][599] = 9'b111111111;
assign micromatrizz[96][600] = 9'b111111111;
assign micromatrizz[96][601] = 9'b111111111;
assign micromatrizz[96][602] = 9'b111111111;
assign micromatrizz[96][603] = 9'b111111111;
assign micromatrizz[96][604] = 9'b111111111;
assign micromatrizz[96][605] = 9'b111111111;
assign micromatrizz[96][606] = 9'b111111111;
assign micromatrizz[96][607] = 9'b111111111;
assign micromatrizz[96][608] = 9'b111111111;
assign micromatrizz[96][609] = 9'b111111111;
assign micromatrizz[96][610] = 9'b111111111;
assign micromatrizz[96][611] = 9'b111111111;
assign micromatrizz[96][612] = 9'b111111111;
assign micromatrizz[96][613] = 9'b111111111;
assign micromatrizz[96][614] = 9'b111111111;
assign micromatrizz[96][615] = 9'b111111111;
assign micromatrizz[96][616] = 9'b111111111;
assign micromatrizz[96][617] = 9'b111111111;
assign micromatrizz[96][618] = 9'b111111111;
assign micromatrizz[96][619] = 9'b111111111;
assign micromatrizz[96][620] = 9'b111111111;
assign micromatrizz[96][621] = 9'b111111111;
assign micromatrizz[96][622] = 9'b111111111;
assign micromatrizz[96][623] = 9'b111111111;
assign micromatrizz[96][624] = 9'b111111111;
assign micromatrizz[96][625] = 9'b111111111;
assign micromatrizz[96][626] = 9'b111111111;
assign micromatrizz[96][627] = 9'b111111111;
assign micromatrizz[96][628] = 9'b111111111;
assign micromatrizz[96][629] = 9'b111111111;
assign micromatrizz[96][630] = 9'b111111111;
assign micromatrizz[96][631] = 9'b111111111;
assign micromatrizz[96][632] = 9'b111111111;
assign micromatrizz[96][633] = 9'b111111111;
assign micromatrizz[96][634] = 9'b111111111;
assign micromatrizz[96][635] = 9'b111111111;
assign micromatrizz[96][636] = 9'b111111111;
assign micromatrizz[96][637] = 9'b111111111;
assign micromatrizz[96][638] = 9'b111111111;
assign micromatrizz[96][639] = 9'b111111111;
assign micromatrizz[97][0] = 9'b111111111;
assign micromatrizz[97][1] = 9'b111111111;
assign micromatrizz[97][2] = 9'b111111111;
assign micromatrizz[97][3] = 9'b111111111;
assign micromatrizz[97][4] = 9'b111111111;
assign micromatrizz[97][5] = 9'b111111111;
assign micromatrizz[97][6] = 9'b111111111;
assign micromatrizz[97][7] = 9'b111111111;
assign micromatrizz[97][8] = 9'b111111111;
assign micromatrizz[97][9] = 9'b111111111;
assign micromatrizz[97][10] = 9'b111111111;
assign micromatrizz[97][11] = 9'b111111111;
assign micromatrizz[97][12] = 9'b111111111;
assign micromatrizz[97][13] = 9'b111111111;
assign micromatrizz[97][14] = 9'b111111111;
assign micromatrizz[97][15] = 9'b111111111;
assign micromatrizz[97][16] = 9'b111111111;
assign micromatrizz[97][17] = 9'b111111111;
assign micromatrizz[97][18] = 9'b111111111;
assign micromatrizz[97][19] = 9'b111111111;
assign micromatrizz[97][20] = 9'b111111111;
assign micromatrizz[97][21] = 9'b111111111;
assign micromatrizz[97][22] = 9'b111111111;
assign micromatrizz[97][23] = 9'b111111111;
assign micromatrizz[97][24] = 9'b111111111;
assign micromatrizz[97][25] = 9'b111111111;
assign micromatrizz[97][26] = 9'b111111111;
assign micromatrizz[97][27] = 9'b111111111;
assign micromatrizz[97][28] = 9'b111111111;
assign micromatrizz[97][29] = 9'b111111111;
assign micromatrizz[97][30] = 9'b111111111;
assign micromatrizz[97][31] = 9'b111111111;
assign micromatrizz[97][32] = 9'b111111111;
assign micromatrizz[97][33] = 9'b111111111;
assign micromatrizz[97][34] = 9'b111111111;
assign micromatrizz[97][35] = 9'b111111111;
assign micromatrizz[97][36] = 9'b111111111;
assign micromatrizz[97][37] = 9'b111111111;
assign micromatrizz[97][38] = 9'b111111111;
assign micromatrizz[97][39] = 9'b111111111;
assign micromatrizz[97][40] = 9'b111111111;
assign micromatrizz[97][41] = 9'b111111111;
assign micromatrizz[97][42] = 9'b111111111;
assign micromatrizz[97][43] = 9'b111111111;
assign micromatrizz[97][44] = 9'b111111111;
assign micromatrizz[97][45] = 9'b111111111;
assign micromatrizz[97][46] = 9'b111111111;
assign micromatrizz[97][47] = 9'b111111111;
assign micromatrizz[97][48] = 9'b111111111;
assign micromatrizz[97][49] = 9'b111111111;
assign micromatrizz[97][50] = 9'b111111111;
assign micromatrizz[97][51] = 9'b111111111;
assign micromatrizz[97][52] = 9'b111111111;
assign micromatrizz[97][53] = 9'b111111111;
assign micromatrizz[97][54] = 9'b111111111;
assign micromatrizz[97][55] = 9'b111111111;
assign micromatrizz[97][56] = 9'b111111111;
assign micromatrizz[97][57] = 9'b111111111;
assign micromatrizz[97][58] = 9'b111111111;
assign micromatrizz[97][59] = 9'b111111111;
assign micromatrizz[97][60] = 9'b111111111;
assign micromatrizz[97][61] = 9'b111111111;
assign micromatrizz[97][62] = 9'b111111111;
assign micromatrizz[97][63] = 9'b111111111;
assign micromatrizz[97][64] = 9'b111111111;
assign micromatrizz[97][65] = 9'b111111111;
assign micromatrizz[97][66] = 9'b111111111;
assign micromatrizz[97][67] = 9'b111111111;
assign micromatrizz[97][68] = 9'b111111111;
assign micromatrizz[97][69] = 9'b111111111;
assign micromatrizz[97][70] = 9'b111111111;
assign micromatrizz[97][71] = 9'b111111111;
assign micromatrizz[97][72] = 9'b111111111;
assign micromatrizz[97][73] = 9'b111111111;
assign micromatrizz[97][74] = 9'b111111111;
assign micromatrizz[97][75] = 9'b111111111;
assign micromatrizz[97][76] = 9'b111111111;
assign micromatrizz[97][77] = 9'b111111111;
assign micromatrizz[97][78] = 9'b111111111;
assign micromatrizz[97][79] = 9'b111111111;
assign micromatrizz[97][80] = 9'b111111111;
assign micromatrizz[97][81] = 9'b111111111;
assign micromatrizz[97][82] = 9'b111111111;
assign micromatrizz[97][83] = 9'b111111111;
assign micromatrizz[97][84] = 9'b111111111;
assign micromatrizz[97][85] = 9'b111111111;
assign micromatrizz[97][86] = 9'b111111111;
assign micromatrizz[97][87] = 9'b111111111;
assign micromatrizz[97][88] = 9'b111111111;
assign micromatrizz[97][89] = 9'b111111111;
assign micromatrizz[97][90] = 9'b111111111;
assign micromatrizz[97][91] = 9'b111111111;
assign micromatrizz[97][92] = 9'b111111111;
assign micromatrizz[97][93] = 9'b111111111;
assign micromatrizz[97][94] = 9'b111111111;
assign micromatrizz[97][95] = 9'b111111111;
assign micromatrizz[97][96] = 9'b111111111;
assign micromatrizz[97][97] = 9'b111111111;
assign micromatrizz[97][98] = 9'b111111111;
assign micromatrizz[97][99] = 9'b111111111;
assign micromatrizz[97][100] = 9'b111111111;
assign micromatrizz[97][101] = 9'b111111111;
assign micromatrizz[97][102] = 9'b111111111;
assign micromatrizz[97][103] = 9'b111111111;
assign micromatrizz[97][104] = 9'b111111111;
assign micromatrizz[97][105] = 9'b111111111;
assign micromatrizz[97][106] = 9'b111111111;
assign micromatrizz[97][107] = 9'b111111111;
assign micromatrizz[97][108] = 9'b111111111;
assign micromatrizz[97][109] = 9'b111111111;
assign micromatrizz[97][110] = 9'b111111111;
assign micromatrizz[97][111] = 9'b111111111;
assign micromatrizz[97][112] = 9'b111111111;
assign micromatrizz[97][113] = 9'b111111111;
assign micromatrizz[97][114] = 9'b111111111;
assign micromatrizz[97][115] = 9'b111111111;
assign micromatrizz[97][116] = 9'b111111111;
assign micromatrizz[97][117] = 9'b111111111;
assign micromatrizz[97][118] = 9'b111111111;
assign micromatrizz[97][119] = 9'b111111111;
assign micromatrizz[97][120] = 9'b111111111;
assign micromatrizz[97][121] = 9'b111111111;
assign micromatrizz[97][122] = 9'b111111111;
assign micromatrizz[97][123] = 9'b111111111;
assign micromatrizz[97][124] = 9'b111111111;
assign micromatrizz[97][125] = 9'b111111111;
assign micromatrizz[97][126] = 9'b111111111;
assign micromatrizz[97][127] = 9'b111111111;
assign micromatrizz[97][128] = 9'b111111111;
assign micromatrizz[97][129] = 9'b111111111;
assign micromatrizz[97][130] = 9'b111111111;
assign micromatrizz[97][131] = 9'b111111111;
assign micromatrizz[97][132] = 9'b111111111;
assign micromatrizz[97][133] = 9'b111111111;
assign micromatrizz[97][134] = 9'b111111111;
assign micromatrizz[97][135] = 9'b111111111;
assign micromatrizz[97][136] = 9'b111111111;
assign micromatrizz[97][137] = 9'b111111111;
assign micromatrizz[97][138] = 9'b111111111;
assign micromatrizz[97][139] = 9'b111111111;
assign micromatrizz[97][140] = 9'b111111111;
assign micromatrizz[97][141] = 9'b111111111;
assign micromatrizz[97][142] = 9'b111111111;
assign micromatrizz[97][143] = 9'b111111111;
assign micromatrizz[97][144] = 9'b111111111;
assign micromatrizz[97][145] = 9'b111111111;
assign micromatrizz[97][146] = 9'b111111111;
assign micromatrizz[97][147] = 9'b111111111;
assign micromatrizz[97][148] = 9'b111111111;
assign micromatrizz[97][149] = 9'b111111111;
assign micromatrizz[97][150] = 9'b111111111;
assign micromatrizz[97][151] = 9'b111111111;
assign micromatrizz[97][152] = 9'b111111111;
assign micromatrizz[97][153] = 9'b111111111;
assign micromatrizz[97][154] = 9'b111111111;
assign micromatrizz[97][155] = 9'b111111111;
assign micromatrizz[97][156] = 9'b111111111;
assign micromatrizz[97][157] = 9'b111111111;
assign micromatrizz[97][158] = 9'b111111111;
assign micromatrizz[97][159] = 9'b111111111;
assign micromatrizz[97][160] = 9'b111111111;
assign micromatrizz[97][161] = 9'b111111111;
assign micromatrizz[97][162] = 9'b111111111;
assign micromatrizz[97][163] = 9'b111111111;
assign micromatrizz[97][164] = 9'b111111111;
assign micromatrizz[97][165] = 9'b111111111;
assign micromatrizz[97][166] = 9'b111111111;
assign micromatrizz[97][167] = 9'b111111111;
assign micromatrizz[97][168] = 9'b111111111;
assign micromatrizz[97][169] = 9'b111111111;
assign micromatrizz[97][170] = 9'b111111111;
assign micromatrizz[97][171] = 9'b111111111;
assign micromatrizz[97][172] = 9'b111111111;
assign micromatrizz[97][173] = 9'b111111111;
assign micromatrizz[97][174] = 9'b111111111;
assign micromatrizz[97][175] = 9'b111111111;
assign micromatrizz[97][176] = 9'b111111111;
assign micromatrizz[97][177] = 9'b111111111;
assign micromatrizz[97][178] = 9'b111111111;
assign micromatrizz[97][179] = 9'b111111111;
assign micromatrizz[97][180] = 9'b111111111;
assign micromatrizz[97][181] = 9'b111111111;
assign micromatrizz[97][182] = 9'b111111111;
assign micromatrizz[97][183] = 9'b111111111;
assign micromatrizz[97][184] = 9'b111111111;
assign micromatrizz[97][185] = 9'b111111111;
assign micromatrizz[97][186] = 9'b111111111;
assign micromatrizz[97][187] = 9'b111111111;
assign micromatrizz[97][188] = 9'b111111111;
assign micromatrizz[97][189] = 9'b111111111;
assign micromatrizz[97][190] = 9'b111111111;
assign micromatrizz[97][191] = 9'b111111111;
assign micromatrizz[97][192] = 9'b111111111;
assign micromatrizz[97][193] = 9'b111111111;
assign micromatrizz[97][194] = 9'b111111111;
assign micromatrizz[97][195] = 9'b111111111;
assign micromatrizz[97][196] = 9'b111111111;
assign micromatrizz[97][197] = 9'b111111111;
assign micromatrizz[97][198] = 9'b111111111;
assign micromatrizz[97][199] = 9'b111111111;
assign micromatrizz[97][200] = 9'b111111111;
assign micromatrizz[97][201] = 9'b111111111;
assign micromatrizz[97][202] = 9'b111111111;
assign micromatrizz[97][203] = 9'b111111111;
assign micromatrizz[97][204] = 9'b111111111;
assign micromatrizz[97][205] = 9'b111111111;
assign micromatrizz[97][206] = 9'b111111111;
assign micromatrizz[97][207] = 9'b111111111;
assign micromatrizz[97][208] = 9'b111111111;
assign micromatrizz[97][209] = 9'b111111111;
assign micromatrizz[97][210] = 9'b111111111;
assign micromatrizz[97][211] = 9'b111111111;
assign micromatrizz[97][212] = 9'b111111111;
assign micromatrizz[97][213] = 9'b111111111;
assign micromatrizz[97][214] = 9'b111111111;
assign micromatrizz[97][215] = 9'b111111111;
assign micromatrizz[97][216] = 9'b111111111;
assign micromatrizz[97][217] = 9'b111111111;
assign micromatrizz[97][218] = 9'b111111111;
assign micromatrizz[97][219] = 9'b111111111;
assign micromatrizz[97][220] = 9'b111111111;
assign micromatrizz[97][221] = 9'b111111111;
assign micromatrizz[97][222] = 9'b111111111;
assign micromatrizz[97][223] = 9'b111111111;
assign micromatrizz[97][224] = 9'b111111111;
assign micromatrizz[97][225] = 9'b111111111;
assign micromatrizz[97][226] = 9'b111111111;
assign micromatrizz[97][227] = 9'b111111111;
assign micromatrizz[97][228] = 9'b111111111;
assign micromatrizz[97][229] = 9'b111111111;
assign micromatrizz[97][230] = 9'b111111111;
assign micromatrizz[97][231] = 9'b111111111;
assign micromatrizz[97][232] = 9'b111111111;
assign micromatrizz[97][233] = 9'b111111111;
assign micromatrizz[97][234] = 9'b111111111;
assign micromatrizz[97][235] = 9'b111111111;
assign micromatrizz[97][236] = 9'b111111111;
assign micromatrizz[97][237] = 9'b111111111;
assign micromatrizz[97][238] = 9'b111111111;
assign micromatrizz[97][239] = 9'b111111111;
assign micromatrizz[97][240] = 9'b111111111;
assign micromatrizz[97][241] = 9'b111111111;
assign micromatrizz[97][242] = 9'b111111111;
assign micromatrizz[97][243] = 9'b111111111;
assign micromatrizz[97][244] = 9'b111111111;
assign micromatrizz[97][245] = 9'b111111111;
assign micromatrizz[97][246] = 9'b111111111;
assign micromatrizz[97][247] = 9'b111111111;
assign micromatrizz[97][248] = 9'b111111111;
assign micromatrizz[97][249] = 9'b111111111;
assign micromatrizz[97][250] = 9'b111111111;
assign micromatrizz[97][251] = 9'b111111111;
assign micromatrizz[97][252] = 9'b111111111;
assign micromatrizz[97][253] = 9'b111111111;
assign micromatrizz[97][254] = 9'b111111111;
assign micromatrizz[97][255] = 9'b111111111;
assign micromatrizz[97][256] = 9'b111111111;
assign micromatrizz[97][257] = 9'b111111111;
assign micromatrizz[97][258] = 9'b111111111;
assign micromatrizz[97][259] = 9'b111111111;
assign micromatrizz[97][260] = 9'b111111111;
assign micromatrizz[97][261] = 9'b111111111;
assign micromatrizz[97][262] = 9'b111111111;
assign micromatrizz[97][263] = 9'b111111111;
assign micromatrizz[97][264] = 9'b111111111;
assign micromatrizz[97][265] = 9'b111111111;
assign micromatrizz[97][266] = 9'b111111111;
assign micromatrizz[97][267] = 9'b111111111;
assign micromatrizz[97][268] = 9'b111111111;
assign micromatrizz[97][269] = 9'b111111111;
assign micromatrizz[97][270] = 9'b111111111;
assign micromatrizz[97][271] = 9'b111111111;
assign micromatrizz[97][272] = 9'b111111111;
assign micromatrizz[97][273] = 9'b111111111;
assign micromatrizz[97][274] = 9'b111111111;
assign micromatrizz[97][275] = 9'b111111111;
assign micromatrizz[97][276] = 9'b111111111;
assign micromatrizz[97][277] = 9'b111111111;
assign micromatrizz[97][278] = 9'b111111111;
assign micromatrizz[97][279] = 9'b111111111;
assign micromatrizz[97][280] = 9'b111111111;
assign micromatrizz[97][281] = 9'b111111111;
assign micromatrizz[97][282] = 9'b111111111;
assign micromatrizz[97][283] = 9'b111111111;
assign micromatrizz[97][284] = 9'b111111111;
assign micromatrizz[97][285] = 9'b111111111;
assign micromatrizz[97][286] = 9'b111111111;
assign micromatrizz[97][287] = 9'b111111111;
assign micromatrizz[97][288] = 9'b111111111;
assign micromatrizz[97][289] = 9'b111111111;
assign micromatrizz[97][290] = 9'b111111111;
assign micromatrizz[97][291] = 9'b111111111;
assign micromatrizz[97][292] = 9'b111111111;
assign micromatrizz[97][293] = 9'b111111111;
assign micromatrizz[97][294] = 9'b111111111;
assign micromatrizz[97][295] = 9'b111111111;
assign micromatrizz[97][296] = 9'b111111111;
assign micromatrizz[97][297] = 9'b111111111;
assign micromatrizz[97][298] = 9'b111111111;
assign micromatrizz[97][299] = 9'b111111111;
assign micromatrizz[97][300] = 9'b111111111;
assign micromatrizz[97][301] = 9'b111111111;
assign micromatrizz[97][302] = 9'b111111111;
assign micromatrizz[97][303] = 9'b111111111;
assign micromatrizz[97][304] = 9'b111111111;
assign micromatrizz[97][305] = 9'b111111111;
assign micromatrizz[97][306] = 9'b111111111;
assign micromatrizz[97][307] = 9'b111111111;
assign micromatrizz[97][308] = 9'b111111111;
assign micromatrizz[97][309] = 9'b111111111;
assign micromatrizz[97][310] = 9'b111111111;
assign micromatrizz[97][311] = 9'b111111111;
assign micromatrizz[97][312] = 9'b111111111;
assign micromatrizz[97][313] = 9'b111111111;
assign micromatrizz[97][314] = 9'b111111111;
assign micromatrizz[97][315] = 9'b111111111;
assign micromatrizz[97][316] = 9'b111111111;
assign micromatrizz[97][317] = 9'b111111111;
assign micromatrizz[97][318] = 9'b111111111;
assign micromatrizz[97][319] = 9'b111111111;
assign micromatrizz[97][320] = 9'b111111111;
assign micromatrizz[97][321] = 9'b111111111;
assign micromatrizz[97][322] = 9'b111111111;
assign micromatrizz[97][323] = 9'b111111111;
assign micromatrizz[97][324] = 9'b111111111;
assign micromatrizz[97][325] = 9'b111111111;
assign micromatrizz[97][326] = 9'b111111111;
assign micromatrizz[97][327] = 9'b111111111;
assign micromatrizz[97][328] = 9'b111111111;
assign micromatrizz[97][329] = 9'b111111111;
assign micromatrizz[97][330] = 9'b111111111;
assign micromatrizz[97][331] = 9'b111111111;
assign micromatrizz[97][332] = 9'b111111111;
assign micromatrizz[97][333] = 9'b111111111;
assign micromatrizz[97][334] = 9'b111111111;
assign micromatrizz[97][335] = 9'b111111111;
assign micromatrizz[97][336] = 9'b111111111;
assign micromatrizz[97][337] = 9'b111111111;
assign micromatrizz[97][338] = 9'b111111111;
assign micromatrizz[97][339] = 9'b111111111;
assign micromatrizz[97][340] = 9'b111111111;
assign micromatrizz[97][341] = 9'b111111111;
assign micromatrizz[97][342] = 9'b111111111;
assign micromatrizz[97][343] = 9'b111111111;
assign micromatrizz[97][344] = 9'b111111111;
assign micromatrizz[97][345] = 9'b111111111;
assign micromatrizz[97][346] = 9'b111111111;
assign micromatrizz[97][347] = 9'b111111111;
assign micromatrizz[97][348] = 9'b111111111;
assign micromatrizz[97][349] = 9'b111111111;
assign micromatrizz[97][350] = 9'b111111111;
assign micromatrizz[97][351] = 9'b111111111;
assign micromatrizz[97][352] = 9'b111111111;
assign micromatrizz[97][353] = 9'b111111111;
assign micromatrizz[97][354] = 9'b111111111;
assign micromatrizz[97][355] = 9'b111111111;
assign micromatrizz[97][356] = 9'b111111111;
assign micromatrizz[97][357] = 9'b111111111;
assign micromatrizz[97][358] = 9'b111111111;
assign micromatrizz[97][359] = 9'b111111111;
assign micromatrizz[97][360] = 9'b111111111;
assign micromatrizz[97][361] = 9'b111111111;
assign micromatrizz[97][362] = 9'b111111111;
assign micromatrizz[97][363] = 9'b111111111;
assign micromatrizz[97][364] = 9'b111111111;
assign micromatrizz[97][365] = 9'b111111111;
assign micromatrizz[97][366] = 9'b111111111;
assign micromatrizz[97][367] = 9'b111111111;
assign micromatrizz[97][368] = 9'b111111111;
assign micromatrizz[97][369] = 9'b111111111;
assign micromatrizz[97][370] = 9'b111111111;
assign micromatrizz[97][371] = 9'b111111111;
assign micromatrizz[97][372] = 9'b111111111;
assign micromatrizz[97][373] = 9'b111111111;
assign micromatrizz[97][374] = 9'b111111111;
assign micromatrizz[97][375] = 9'b111111111;
assign micromatrizz[97][376] = 9'b111111111;
assign micromatrizz[97][377] = 9'b111111111;
assign micromatrizz[97][378] = 9'b111111111;
assign micromatrizz[97][379] = 9'b111111111;
assign micromatrizz[97][380] = 9'b111111111;
assign micromatrizz[97][381] = 9'b111111111;
assign micromatrizz[97][382] = 9'b111111111;
assign micromatrizz[97][383] = 9'b111111111;
assign micromatrizz[97][384] = 9'b111111111;
assign micromatrizz[97][385] = 9'b111111111;
assign micromatrizz[97][386] = 9'b111111111;
assign micromatrizz[97][387] = 9'b111111111;
assign micromatrizz[97][388] = 9'b111111111;
assign micromatrizz[97][389] = 9'b111111111;
assign micromatrizz[97][390] = 9'b111111111;
assign micromatrizz[97][391] = 9'b111111111;
assign micromatrizz[97][392] = 9'b111111111;
assign micromatrizz[97][393] = 9'b111111111;
assign micromatrizz[97][394] = 9'b111111111;
assign micromatrizz[97][395] = 9'b111111111;
assign micromatrizz[97][396] = 9'b111111111;
assign micromatrizz[97][397] = 9'b111111111;
assign micromatrizz[97][398] = 9'b111111111;
assign micromatrizz[97][399] = 9'b111111111;
assign micromatrizz[97][400] = 9'b111111111;
assign micromatrizz[97][401] = 9'b111111111;
assign micromatrizz[97][402] = 9'b111111111;
assign micromatrizz[97][403] = 9'b111111111;
assign micromatrizz[97][404] = 9'b111111111;
assign micromatrizz[97][405] = 9'b111111111;
assign micromatrizz[97][406] = 9'b111111111;
assign micromatrizz[97][407] = 9'b111111111;
assign micromatrizz[97][408] = 9'b111111111;
assign micromatrizz[97][409] = 9'b111111111;
assign micromatrizz[97][410] = 9'b111111111;
assign micromatrizz[97][411] = 9'b111111111;
assign micromatrizz[97][412] = 9'b111111111;
assign micromatrizz[97][413] = 9'b111111111;
assign micromatrizz[97][414] = 9'b111111111;
assign micromatrizz[97][415] = 9'b111111111;
assign micromatrizz[97][416] = 9'b111111111;
assign micromatrizz[97][417] = 9'b111111111;
assign micromatrizz[97][418] = 9'b111111111;
assign micromatrizz[97][419] = 9'b111111111;
assign micromatrizz[97][420] = 9'b111111111;
assign micromatrizz[97][421] = 9'b111111111;
assign micromatrizz[97][422] = 9'b111111111;
assign micromatrizz[97][423] = 9'b111111111;
assign micromatrizz[97][424] = 9'b111111111;
assign micromatrizz[97][425] = 9'b111111111;
assign micromatrizz[97][426] = 9'b111111111;
assign micromatrizz[97][427] = 9'b111111111;
assign micromatrizz[97][428] = 9'b111111111;
assign micromatrizz[97][429] = 9'b111111111;
assign micromatrizz[97][430] = 9'b111111111;
assign micromatrizz[97][431] = 9'b111111111;
assign micromatrizz[97][432] = 9'b111111111;
assign micromatrizz[97][433] = 9'b111111111;
assign micromatrizz[97][434] = 9'b111111111;
assign micromatrizz[97][435] = 9'b111111111;
assign micromatrizz[97][436] = 9'b111111111;
assign micromatrizz[97][437] = 9'b111111111;
assign micromatrizz[97][438] = 9'b111111111;
assign micromatrizz[97][439] = 9'b111111111;
assign micromatrizz[97][440] = 9'b111111111;
assign micromatrizz[97][441] = 9'b111111111;
assign micromatrizz[97][442] = 9'b111111111;
assign micromatrizz[97][443] = 9'b111111111;
assign micromatrizz[97][444] = 9'b111111111;
assign micromatrizz[97][445] = 9'b111111111;
assign micromatrizz[97][446] = 9'b111111111;
assign micromatrizz[97][447] = 9'b111111111;
assign micromatrizz[97][448] = 9'b111111111;
assign micromatrizz[97][449] = 9'b111111111;
assign micromatrizz[97][450] = 9'b111111111;
assign micromatrizz[97][451] = 9'b111111111;
assign micromatrizz[97][452] = 9'b111111111;
assign micromatrizz[97][453] = 9'b111111111;
assign micromatrizz[97][454] = 9'b111111111;
assign micromatrizz[97][455] = 9'b111111111;
assign micromatrizz[97][456] = 9'b111111111;
assign micromatrizz[97][457] = 9'b111111111;
assign micromatrizz[97][458] = 9'b111111111;
assign micromatrizz[97][459] = 9'b111111111;
assign micromatrizz[97][460] = 9'b111111111;
assign micromatrizz[97][461] = 9'b111111111;
assign micromatrizz[97][462] = 9'b111111111;
assign micromatrizz[97][463] = 9'b111111111;
assign micromatrizz[97][464] = 9'b111111111;
assign micromatrizz[97][465] = 9'b111111111;
assign micromatrizz[97][466] = 9'b111111111;
assign micromatrizz[97][467] = 9'b111111111;
assign micromatrizz[97][468] = 9'b111111111;
assign micromatrizz[97][469] = 9'b111111111;
assign micromatrizz[97][470] = 9'b111111111;
assign micromatrizz[97][471] = 9'b111111111;
assign micromatrizz[97][472] = 9'b111111111;
assign micromatrizz[97][473] = 9'b111111111;
assign micromatrizz[97][474] = 9'b111111111;
assign micromatrizz[97][475] = 9'b111111111;
assign micromatrizz[97][476] = 9'b111111111;
assign micromatrizz[97][477] = 9'b111111111;
assign micromatrizz[97][478] = 9'b111111111;
assign micromatrizz[97][479] = 9'b111111111;
assign micromatrizz[97][480] = 9'b111111111;
assign micromatrizz[97][481] = 9'b111111111;
assign micromatrizz[97][482] = 9'b111111111;
assign micromatrizz[97][483] = 9'b111111111;
assign micromatrizz[97][484] = 9'b111111111;
assign micromatrizz[97][485] = 9'b111111111;
assign micromatrizz[97][486] = 9'b111111111;
assign micromatrizz[97][487] = 9'b111111111;
assign micromatrizz[97][488] = 9'b111111111;
assign micromatrizz[97][489] = 9'b111111111;
assign micromatrizz[97][490] = 9'b111111111;
assign micromatrizz[97][491] = 9'b111111111;
assign micromatrizz[97][492] = 9'b111111111;
assign micromatrizz[97][493] = 9'b111111111;
assign micromatrizz[97][494] = 9'b111111111;
assign micromatrizz[97][495] = 9'b111111111;
assign micromatrizz[97][496] = 9'b111111111;
assign micromatrizz[97][497] = 9'b111111111;
assign micromatrizz[97][498] = 9'b111111111;
assign micromatrizz[97][499] = 9'b111111111;
assign micromatrizz[97][500] = 9'b111111111;
assign micromatrizz[97][501] = 9'b111111111;
assign micromatrizz[97][502] = 9'b111111111;
assign micromatrizz[97][503] = 9'b111111111;
assign micromatrizz[97][504] = 9'b111111111;
assign micromatrizz[97][505] = 9'b111111111;
assign micromatrizz[97][506] = 9'b111111111;
assign micromatrizz[97][507] = 9'b111111111;
assign micromatrizz[97][508] = 9'b111111111;
assign micromatrizz[97][509] = 9'b111111111;
assign micromatrizz[97][510] = 9'b111111111;
assign micromatrizz[97][511] = 9'b111111111;
assign micromatrizz[97][512] = 9'b111111111;
assign micromatrizz[97][513] = 9'b111111111;
assign micromatrizz[97][514] = 9'b111111111;
assign micromatrizz[97][515] = 9'b111111111;
assign micromatrizz[97][516] = 9'b111111111;
assign micromatrizz[97][517] = 9'b111111111;
assign micromatrizz[97][518] = 9'b111111111;
assign micromatrizz[97][519] = 9'b111111111;
assign micromatrizz[97][520] = 9'b111111111;
assign micromatrizz[97][521] = 9'b111111111;
assign micromatrizz[97][522] = 9'b111111111;
assign micromatrizz[97][523] = 9'b111111111;
assign micromatrizz[97][524] = 9'b111111111;
assign micromatrizz[97][525] = 9'b111111111;
assign micromatrizz[97][526] = 9'b111111111;
assign micromatrizz[97][527] = 9'b111111111;
assign micromatrizz[97][528] = 9'b111111111;
assign micromatrizz[97][529] = 9'b111111111;
assign micromatrizz[97][530] = 9'b111111111;
assign micromatrizz[97][531] = 9'b111111111;
assign micromatrizz[97][532] = 9'b111111111;
assign micromatrizz[97][533] = 9'b111111111;
assign micromatrizz[97][534] = 9'b111111111;
assign micromatrizz[97][535] = 9'b111111111;
assign micromatrizz[97][536] = 9'b111111111;
assign micromatrizz[97][537] = 9'b111111111;
assign micromatrizz[97][538] = 9'b111111111;
assign micromatrizz[97][539] = 9'b111111111;
assign micromatrizz[97][540] = 9'b111111111;
assign micromatrizz[97][541] = 9'b111111111;
assign micromatrizz[97][542] = 9'b111111111;
assign micromatrizz[97][543] = 9'b111111111;
assign micromatrizz[97][544] = 9'b111111111;
assign micromatrizz[97][545] = 9'b111111111;
assign micromatrizz[97][546] = 9'b111111111;
assign micromatrizz[97][547] = 9'b111111111;
assign micromatrizz[97][548] = 9'b111111111;
assign micromatrizz[97][549] = 9'b111111111;
assign micromatrizz[97][550] = 9'b111111111;
assign micromatrizz[97][551] = 9'b111111111;
assign micromatrizz[97][552] = 9'b111111111;
assign micromatrizz[97][553] = 9'b111111111;
assign micromatrizz[97][554] = 9'b111111111;
assign micromatrizz[97][555] = 9'b111111111;
assign micromatrizz[97][556] = 9'b111111111;
assign micromatrizz[97][557] = 9'b111111111;
assign micromatrizz[97][558] = 9'b111111111;
assign micromatrizz[97][559] = 9'b111111111;
assign micromatrizz[97][560] = 9'b111111111;
assign micromatrizz[97][561] = 9'b111111111;
assign micromatrizz[97][562] = 9'b111111111;
assign micromatrizz[97][563] = 9'b111111111;
assign micromatrizz[97][564] = 9'b111111111;
assign micromatrizz[97][565] = 9'b111111111;
assign micromatrizz[97][566] = 9'b111111111;
assign micromatrizz[97][567] = 9'b111111111;
assign micromatrizz[97][568] = 9'b111111111;
assign micromatrizz[97][569] = 9'b111111111;
assign micromatrizz[97][570] = 9'b111111111;
assign micromatrizz[97][571] = 9'b111111111;
assign micromatrizz[97][572] = 9'b111111111;
assign micromatrizz[97][573] = 9'b111111111;
assign micromatrizz[97][574] = 9'b111111111;
assign micromatrizz[97][575] = 9'b111111111;
assign micromatrizz[97][576] = 9'b111111111;
assign micromatrizz[97][577] = 9'b111111111;
assign micromatrizz[97][578] = 9'b111111111;
assign micromatrizz[97][579] = 9'b111111111;
assign micromatrizz[97][580] = 9'b111111111;
assign micromatrizz[97][581] = 9'b111111111;
assign micromatrizz[97][582] = 9'b111111111;
assign micromatrizz[97][583] = 9'b111111111;
assign micromatrizz[97][584] = 9'b111111111;
assign micromatrizz[97][585] = 9'b111111111;
assign micromatrizz[97][586] = 9'b111111111;
assign micromatrizz[97][587] = 9'b111111111;
assign micromatrizz[97][588] = 9'b111111111;
assign micromatrizz[97][589] = 9'b111111111;
assign micromatrizz[97][590] = 9'b111111111;
assign micromatrizz[97][591] = 9'b111111111;
assign micromatrizz[97][592] = 9'b111111111;
assign micromatrizz[97][593] = 9'b111111111;
assign micromatrizz[97][594] = 9'b111111111;
assign micromatrizz[97][595] = 9'b111111111;
assign micromatrizz[97][596] = 9'b111111111;
assign micromatrizz[97][597] = 9'b111111111;
assign micromatrizz[97][598] = 9'b111111111;
assign micromatrizz[97][599] = 9'b111111111;
assign micromatrizz[97][600] = 9'b111111111;
assign micromatrizz[97][601] = 9'b111111111;
assign micromatrizz[97][602] = 9'b111111111;
assign micromatrizz[97][603] = 9'b111111111;
assign micromatrizz[97][604] = 9'b111111111;
assign micromatrizz[97][605] = 9'b111111111;
assign micromatrizz[97][606] = 9'b111111111;
assign micromatrizz[97][607] = 9'b111111111;
assign micromatrizz[97][608] = 9'b111111111;
assign micromatrizz[97][609] = 9'b111111111;
assign micromatrizz[97][610] = 9'b111111111;
assign micromatrizz[97][611] = 9'b111111111;
assign micromatrizz[97][612] = 9'b111111111;
assign micromatrizz[97][613] = 9'b111111111;
assign micromatrizz[97][614] = 9'b111111111;
assign micromatrizz[97][615] = 9'b111111111;
assign micromatrizz[97][616] = 9'b111111111;
assign micromatrizz[97][617] = 9'b111111111;
assign micromatrizz[97][618] = 9'b111111111;
assign micromatrizz[97][619] = 9'b111111111;
assign micromatrizz[97][620] = 9'b111111111;
assign micromatrizz[97][621] = 9'b111111111;
assign micromatrizz[97][622] = 9'b111111111;
assign micromatrizz[97][623] = 9'b111111111;
assign micromatrizz[97][624] = 9'b111111111;
assign micromatrizz[97][625] = 9'b111111111;
assign micromatrizz[97][626] = 9'b111111111;
assign micromatrizz[97][627] = 9'b111111111;
assign micromatrizz[97][628] = 9'b111111111;
assign micromatrizz[97][629] = 9'b111111111;
assign micromatrizz[97][630] = 9'b111111111;
assign micromatrizz[97][631] = 9'b111111111;
assign micromatrizz[97][632] = 9'b111111111;
assign micromatrizz[97][633] = 9'b111111111;
assign micromatrizz[97][634] = 9'b111111111;
assign micromatrizz[97][635] = 9'b111111111;
assign micromatrizz[97][636] = 9'b111111111;
assign micromatrizz[97][637] = 9'b111111111;
assign micromatrizz[97][638] = 9'b111111111;
assign micromatrizz[97][639] = 9'b111111111;
assign micromatrizz[98][0] = 9'b111111111;
assign micromatrizz[98][1] = 9'b111111111;
assign micromatrizz[98][2] = 9'b111111111;
assign micromatrizz[98][3] = 9'b111111111;
assign micromatrizz[98][4] = 9'b111111111;
assign micromatrizz[98][5] = 9'b111111111;
assign micromatrizz[98][6] = 9'b111111111;
assign micromatrizz[98][7] = 9'b111111111;
assign micromatrizz[98][8] = 9'b111111111;
assign micromatrizz[98][9] = 9'b111111111;
assign micromatrizz[98][10] = 9'b111111111;
assign micromatrizz[98][11] = 9'b111111111;
assign micromatrizz[98][12] = 9'b111111111;
assign micromatrizz[98][13] = 9'b111111111;
assign micromatrizz[98][14] = 9'b111111111;
assign micromatrizz[98][15] = 9'b111111111;
assign micromatrizz[98][16] = 9'b111111111;
assign micromatrizz[98][17] = 9'b111111111;
assign micromatrizz[98][18] = 9'b111111111;
assign micromatrizz[98][19] = 9'b111111111;
assign micromatrizz[98][20] = 9'b111111111;
assign micromatrizz[98][21] = 9'b111111111;
assign micromatrizz[98][22] = 9'b111111111;
assign micromatrizz[98][23] = 9'b111111111;
assign micromatrizz[98][24] = 9'b111111111;
assign micromatrizz[98][25] = 9'b111111111;
assign micromatrizz[98][26] = 9'b111111111;
assign micromatrizz[98][27] = 9'b111111111;
assign micromatrizz[98][28] = 9'b111111111;
assign micromatrizz[98][29] = 9'b111111111;
assign micromatrizz[98][30] = 9'b111111111;
assign micromatrizz[98][31] = 9'b111111111;
assign micromatrizz[98][32] = 9'b111111111;
assign micromatrizz[98][33] = 9'b111111111;
assign micromatrizz[98][34] = 9'b111111111;
assign micromatrizz[98][35] = 9'b111111111;
assign micromatrizz[98][36] = 9'b111111111;
assign micromatrizz[98][37] = 9'b111111111;
assign micromatrizz[98][38] = 9'b111111111;
assign micromatrizz[98][39] = 9'b111111111;
assign micromatrizz[98][40] = 9'b111111111;
assign micromatrizz[98][41] = 9'b111111111;
assign micromatrizz[98][42] = 9'b111111111;
assign micromatrizz[98][43] = 9'b111111111;
assign micromatrizz[98][44] = 9'b111111111;
assign micromatrizz[98][45] = 9'b111111111;
assign micromatrizz[98][46] = 9'b111111111;
assign micromatrizz[98][47] = 9'b111111111;
assign micromatrizz[98][48] = 9'b111111111;
assign micromatrizz[98][49] = 9'b111111111;
assign micromatrizz[98][50] = 9'b111111111;
assign micromatrizz[98][51] = 9'b111111111;
assign micromatrizz[98][52] = 9'b111111111;
assign micromatrizz[98][53] = 9'b111111111;
assign micromatrizz[98][54] = 9'b111111111;
assign micromatrizz[98][55] = 9'b111111111;
assign micromatrizz[98][56] = 9'b111111111;
assign micromatrizz[98][57] = 9'b111111111;
assign micromatrizz[98][58] = 9'b111111111;
assign micromatrizz[98][59] = 9'b111111111;
assign micromatrizz[98][60] = 9'b111111111;
assign micromatrizz[98][61] = 9'b111111111;
assign micromatrizz[98][62] = 9'b111111111;
assign micromatrizz[98][63] = 9'b111111111;
assign micromatrizz[98][64] = 9'b111111111;
assign micromatrizz[98][65] = 9'b111111111;
assign micromatrizz[98][66] = 9'b111111111;
assign micromatrizz[98][67] = 9'b111111111;
assign micromatrizz[98][68] = 9'b111111111;
assign micromatrizz[98][69] = 9'b111111111;
assign micromatrizz[98][70] = 9'b111111111;
assign micromatrizz[98][71] = 9'b111111111;
assign micromatrizz[98][72] = 9'b111111111;
assign micromatrizz[98][73] = 9'b111111111;
assign micromatrizz[98][74] = 9'b111111111;
assign micromatrizz[98][75] = 9'b111111111;
assign micromatrizz[98][76] = 9'b111111111;
assign micromatrizz[98][77] = 9'b111111111;
assign micromatrizz[98][78] = 9'b111111111;
assign micromatrizz[98][79] = 9'b111111111;
assign micromatrizz[98][80] = 9'b111111111;
assign micromatrizz[98][81] = 9'b111111111;
assign micromatrizz[98][82] = 9'b111111111;
assign micromatrizz[98][83] = 9'b111111111;
assign micromatrizz[98][84] = 9'b111111111;
assign micromatrizz[98][85] = 9'b111111111;
assign micromatrizz[98][86] = 9'b111111111;
assign micromatrizz[98][87] = 9'b111111111;
assign micromatrizz[98][88] = 9'b111111111;
assign micromatrizz[98][89] = 9'b111111111;
assign micromatrizz[98][90] = 9'b111111111;
assign micromatrizz[98][91] = 9'b111111111;
assign micromatrizz[98][92] = 9'b111111111;
assign micromatrizz[98][93] = 9'b111111111;
assign micromatrizz[98][94] = 9'b111111111;
assign micromatrizz[98][95] = 9'b111111111;
assign micromatrizz[98][96] = 9'b111111111;
assign micromatrizz[98][97] = 9'b111111111;
assign micromatrizz[98][98] = 9'b111111111;
assign micromatrizz[98][99] = 9'b111111111;
assign micromatrizz[98][100] = 9'b111111111;
assign micromatrizz[98][101] = 9'b111111111;
assign micromatrizz[98][102] = 9'b111111111;
assign micromatrizz[98][103] = 9'b111111111;
assign micromatrizz[98][104] = 9'b111111111;
assign micromatrizz[98][105] = 9'b111111111;
assign micromatrizz[98][106] = 9'b111111111;
assign micromatrizz[98][107] = 9'b111111111;
assign micromatrizz[98][108] = 9'b111111111;
assign micromatrizz[98][109] = 9'b111111111;
assign micromatrizz[98][110] = 9'b111111111;
assign micromatrizz[98][111] = 9'b111111111;
assign micromatrizz[98][112] = 9'b111111111;
assign micromatrizz[98][113] = 9'b111111111;
assign micromatrizz[98][114] = 9'b111111111;
assign micromatrizz[98][115] = 9'b111111111;
assign micromatrizz[98][116] = 9'b111111111;
assign micromatrizz[98][117] = 9'b111111111;
assign micromatrizz[98][118] = 9'b111111111;
assign micromatrizz[98][119] = 9'b111111111;
assign micromatrizz[98][120] = 9'b111111111;
assign micromatrizz[98][121] = 9'b111111111;
assign micromatrizz[98][122] = 9'b111111111;
assign micromatrizz[98][123] = 9'b111111111;
assign micromatrizz[98][124] = 9'b111111111;
assign micromatrizz[98][125] = 9'b111111111;
assign micromatrizz[98][126] = 9'b111111111;
assign micromatrizz[98][127] = 9'b111111111;
assign micromatrizz[98][128] = 9'b111111111;
assign micromatrizz[98][129] = 9'b111111111;
assign micromatrizz[98][130] = 9'b111111111;
assign micromatrizz[98][131] = 9'b111111111;
assign micromatrizz[98][132] = 9'b111111111;
assign micromatrizz[98][133] = 9'b111111111;
assign micromatrizz[98][134] = 9'b111111111;
assign micromatrizz[98][135] = 9'b111111111;
assign micromatrizz[98][136] = 9'b111111111;
assign micromatrizz[98][137] = 9'b111111111;
assign micromatrizz[98][138] = 9'b111111111;
assign micromatrizz[98][139] = 9'b111111111;
assign micromatrizz[98][140] = 9'b111111111;
assign micromatrizz[98][141] = 9'b111111111;
assign micromatrizz[98][142] = 9'b111111111;
assign micromatrizz[98][143] = 9'b111111111;
assign micromatrizz[98][144] = 9'b111111111;
assign micromatrizz[98][145] = 9'b111111111;
assign micromatrizz[98][146] = 9'b111111111;
assign micromatrizz[98][147] = 9'b111111111;
assign micromatrizz[98][148] = 9'b111111111;
assign micromatrizz[98][149] = 9'b111111111;
assign micromatrizz[98][150] = 9'b111111111;
assign micromatrizz[98][151] = 9'b111111111;
assign micromatrizz[98][152] = 9'b111111111;
assign micromatrizz[98][153] = 9'b111111111;
assign micromatrizz[98][154] = 9'b111111111;
assign micromatrizz[98][155] = 9'b111111111;
assign micromatrizz[98][156] = 9'b111111111;
assign micromatrizz[98][157] = 9'b111111111;
assign micromatrizz[98][158] = 9'b111111111;
assign micromatrizz[98][159] = 9'b111111111;
assign micromatrizz[98][160] = 9'b111111111;
assign micromatrizz[98][161] = 9'b111111111;
assign micromatrizz[98][162] = 9'b111111111;
assign micromatrizz[98][163] = 9'b111111111;
assign micromatrizz[98][164] = 9'b111111111;
assign micromatrizz[98][165] = 9'b111111111;
assign micromatrizz[98][166] = 9'b111111111;
assign micromatrizz[98][167] = 9'b111111111;
assign micromatrizz[98][168] = 9'b111111111;
assign micromatrizz[98][169] = 9'b111111111;
assign micromatrizz[98][170] = 9'b111111111;
assign micromatrizz[98][171] = 9'b111111111;
assign micromatrizz[98][172] = 9'b111111111;
assign micromatrizz[98][173] = 9'b111111111;
assign micromatrizz[98][174] = 9'b111111111;
assign micromatrizz[98][175] = 9'b111111111;
assign micromatrizz[98][176] = 9'b111111111;
assign micromatrizz[98][177] = 9'b111111111;
assign micromatrizz[98][178] = 9'b111111111;
assign micromatrizz[98][179] = 9'b111111111;
assign micromatrizz[98][180] = 9'b111111111;
assign micromatrizz[98][181] = 9'b111111111;
assign micromatrizz[98][182] = 9'b111111111;
assign micromatrizz[98][183] = 9'b111111111;
assign micromatrizz[98][184] = 9'b111111111;
assign micromatrizz[98][185] = 9'b111111111;
assign micromatrizz[98][186] = 9'b111111111;
assign micromatrizz[98][187] = 9'b111111111;
assign micromatrizz[98][188] = 9'b111111111;
assign micromatrizz[98][189] = 9'b111111111;
assign micromatrizz[98][190] = 9'b111111111;
assign micromatrizz[98][191] = 9'b111111111;
assign micromatrizz[98][192] = 9'b111111111;
assign micromatrizz[98][193] = 9'b111111111;
assign micromatrizz[98][194] = 9'b111111111;
assign micromatrizz[98][195] = 9'b111111111;
assign micromatrizz[98][196] = 9'b111111111;
assign micromatrizz[98][197] = 9'b111111111;
assign micromatrizz[98][198] = 9'b111111111;
assign micromatrizz[98][199] = 9'b111111111;
assign micromatrizz[98][200] = 9'b111111111;
assign micromatrizz[98][201] = 9'b111111111;
assign micromatrizz[98][202] = 9'b111111111;
assign micromatrizz[98][203] = 9'b111111111;
assign micromatrizz[98][204] = 9'b111111111;
assign micromatrizz[98][205] = 9'b111111111;
assign micromatrizz[98][206] = 9'b111111111;
assign micromatrizz[98][207] = 9'b111111111;
assign micromatrizz[98][208] = 9'b111111111;
assign micromatrizz[98][209] = 9'b111111111;
assign micromatrizz[98][210] = 9'b111111111;
assign micromatrizz[98][211] = 9'b111111111;
assign micromatrizz[98][212] = 9'b111111111;
assign micromatrizz[98][213] = 9'b111111111;
assign micromatrizz[98][214] = 9'b111111111;
assign micromatrizz[98][215] = 9'b111111111;
assign micromatrizz[98][216] = 9'b111111111;
assign micromatrizz[98][217] = 9'b111111111;
assign micromatrizz[98][218] = 9'b111111111;
assign micromatrizz[98][219] = 9'b111111111;
assign micromatrizz[98][220] = 9'b111111111;
assign micromatrizz[98][221] = 9'b111111111;
assign micromatrizz[98][222] = 9'b111111111;
assign micromatrizz[98][223] = 9'b111111111;
assign micromatrizz[98][224] = 9'b111111111;
assign micromatrizz[98][225] = 9'b111111111;
assign micromatrizz[98][226] = 9'b111111111;
assign micromatrizz[98][227] = 9'b111111111;
assign micromatrizz[98][228] = 9'b111111111;
assign micromatrizz[98][229] = 9'b111111111;
assign micromatrizz[98][230] = 9'b111111111;
assign micromatrizz[98][231] = 9'b111111111;
assign micromatrizz[98][232] = 9'b111111111;
assign micromatrizz[98][233] = 9'b111111111;
assign micromatrizz[98][234] = 9'b111111111;
assign micromatrizz[98][235] = 9'b111111111;
assign micromatrizz[98][236] = 9'b111111111;
assign micromatrizz[98][237] = 9'b111111111;
assign micromatrizz[98][238] = 9'b111111111;
assign micromatrizz[98][239] = 9'b111111111;
assign micromatrizz[98][240] = 9'b111111111;
assign micromatrizz[98][241] = 9'b111111111;
assign micromatrizz[98][242] = 9'b111111111;
assign micromatrizz[98][243] = 9'b111111111;
assign micromatrizz[98][244] = 9'b111111111;
assign micromatrizz[98][245] = 9'b111111111;
assign micromatrizz[98][246] = 9'b111111111;
assign micromatrizz[98][247] = 9'b111111111;
assign micromatrizz[98][248] = 9'b111111111;
assign micromatrizz[98][249] = 9'b111111111;
assign micromatrizz[98][250] = 9'b111111111;
assign micromatrizz[98][251] = 9'b111111111;
assign micromatrizz[98][252] = 9'b111111111;
assign micromatrizz[98][253] = 9'b111111111;
assign micromatrizz[98][254] = 9'b111111111;
assign micromatrizz[98][255] = 9'b111111111;
assign micromatrizz[98][256] = 9'b111111111;
assign micromatrizz[98][257] = 9'b111111111;
assign micromatrizz[98][258] = 9'b111111111;
assign micromatrizz[98][259] = 9'b111111111;
assign micromatrizz[98][260] = 9'b111111111;
assign micromatrizz[98][261] = 9'b111111111;
assign micromatrizz[98][262] = 9'b111111111;
assign micromatrizz[98][263] = 9'b111111111;
assign micromatrizz[98][264] = 9'b111111111;
assign micromatrizz[98][265] = 9'b111111111;
assign micromatrizz[98][266] = 9'b111111111;
assign micromatrizz[98][267] = 9'b111111111;
assign micromatrizz[98][268] = 9'b111111111;
assign micromatrizz[98][269] = 9'b111111111;
assign micromatrizz[98][270] = 9'b111111111;
assign micromatrizz[98][271] = 9'b111111111;
assign micromatrizz[98][272] = 9'b111111111;
assign micromatrizz[98][273] = 9'b111111111;
assign micromatrizz[98][274] = 9'b111111111;
assign micromatrizz[98][275] = 9'b111111111;
assign micromatrizz[98][276] = 9'b111111111;
assign micromatrizz[98][277] = 9'b111111111;
assign micromatrizz[98][278] = 9'b111111111;
assign micromatrizz[98][279] = 9'b111111111;
assign micromatrizz[98][280] = 9'b111111111;
assign micromatrizz[98][281] = 9'b111111111;
assign micromatrizz[98][282] = 9'b111111111;
assign micromatrizz[98][283] = 9'b111111111;
assign micromatrizz[98][284] = 9'b111111111;
assign micromatrizz[98][285] = 9'b111111111;
assign micromatrizz[98][286] = 9'b111111111;
assign micromatrizz[98][287] = 9'b111111111;
assign micromatrizz[98][288] = 9'b111111111;
assign micromatrizz[98][289] = 9'b111111111;
assign micromatrizz[98][290] = 9'b111111111;
assign micromatrizz[98][291] = 9'b111111111;
assign micromatrizz[98][292] = 9'b111111111;
assign micromatrizz[98][293] = 9'b111111111;
assign micromatrizz[98][294] = 9'b111111111;
assign micromatrizz[98][295] = 9'b111111111;
assign micromatrizz[98][296] = 9'b111111111;
assign micromatrizz[98][297] = 9'b111111111;
assign micromatrizz[98][298] = 9'b111111111;
assign micromatrizz[98][299] = 9'b111111111;
assign micromatrizz[98][300] = 9'b111111111;
assign micromatrizz[98][301] = 9'b111111111;
assign micromatrizz[98][302] = 9'b111111111;
assign micromatrizz[98][303] = 9'b111111111;
assign micromatrizz[98][304] = 9'b111111111;
assign micromatrizz[98][305] = 9'b111111111;
assign micromatrizz[98][306] = 9'b111111111;
assign micromatrizz[98][307] = 9'b111111111;
assign micromatrizz[98][308] = 9'b111111111;
assign micromatrizz[98][309] = 9'b111111111;
assign micromatrizz[98][310] = 9'b111111111;
assign micromatrizz[98][311] = 9'b111111111;
assign micromatrizz[98][312] = 9'b111111111;
assign micromatrizz[98][313] = 9'b111111111;
assign micromatrizz[98][314] = 9'b111111111;
assign micromatrizz[98][315] = 9'b111111111;
assign micromatrizz[98][316] = 9'b111111111;
assign micromatrizz[98][317] = 9'b111111111;
assign micromatrizz[98][318] = 9'b111111111;
assign micromatrizz[98][319] = 9'b111111111;
assign micromatrizz[98][320] = 9'b111111111;
assign micromatrizz[98][321] = 9'b111111111;
assign micromatrizz[98][322] = 9'b111111111;
assign micromatrizz[98][323] = 9'b111111111;
assign micromatrizz[98][324] = 9'b111111111;
assign micromatrizz[98][325] = 9'b111111111;
assign micromatrizz[98][326] = 9'b111111111;
assign micromatrizz[98][327] = 9'b111111111;
assign micromatrizz[98][328] = 9'b111111111;
assign micromatrizz[98][329] = 9'b111111111;
assign micromatrizz[98][330] = 9'b111111111;
assign micromatrizz[98][331] = 9'b111111111;
assign micromatrizz[98][332] = 9'b111111111;
assign micromatrizz[98][333] = 9'b111111111;
assign micromatrizz[98][334] = 9'b111111111;
assign micromatrizz[98][335] = 9'b111111111;
assign micromatrizz[98][336] = 9'b111111111;
assign micromatrizz[98][337] = 9'b111111111;
assign micromatrizz[98][338] = 9'b111111111;
assign micromatrizz[98][339] = 9'b111111111;
assign micromatrizz[98][340] = 9'b111111111;
assign micromatrizz[98][341] = 9'b111111111;
assign micromatrizz[98][342] = 9'b111111111;
assign micromatrizz[98][343] = 9'b111111111;
assign micromatrizz[98][344] = 9'b111111111;
assign micromatrizz[98][345] = 9'b111111111;
assign micromatrizz[98][346] = 9'b111111111;
assign micromatrizz[98][347] = 9'b111111111;
assign micromatrizz[98][348] = 9'b111111111;
assign micromatrizz[98][349] = 9'b111111111;
assign micromatrizz[98][350] = 9'b111111111;
assign micromatrizz[98][351] = 9'b111111111;
assign micromatrizz[98][352] = 9'b111111111;
assign micromatrizz[98][353] = 9'b111111111;
assign micromatrizz[98][354] = 9'b111111111;
assign micromatrizz[98][355] = 9'b111111111;
assign micromatrizz[98][356] = 9'b111111111;
assign micromatrizz[98][357] = 9'b111111111;
assign micromatrizz[98][358] = 9'b111111111;
assign micromatrizz[98][359] = 9'b111111111;
assign micromatrizz[98][360] = 9'b111111111;
assign micromatrizz[98][361] = 9'b111111111;
assign micromatrizz[98][362] = 9'b111111111;
assign micromatrizz[98][363] = 9'b111111111;
assign micromatrizz[98][364] = 9'b111111111;
assign micromatrizz[98][365] = 9'b111111111;
assign micromatrizz[98][366] = 9'b111111111;
assign micromatrizz[98][367] = 9'b111111111;
assign micromatrizz[98][368] = 9'b111111111;
assign micromatrizz[98][369] = 9'b111111111;
assign micromatrizz[98][370] = 9'b111111111;
assign micromatrizz[98][371] = 9'b111111111;
assign micromatrizz[98][372] = 9'b111111111;
assign micromatrizz[98][373] = 9'b111111111;
assign micromatrizz[98][374] = 9'b111111111;
assign micromatrizz[98][375] = 9'b111111111;
assign micromatrizz[98][376] = 9'b111111111;
assign micromatrizz[98][377] = 9'b111111111;
assign micromatrizz[98][378] = 9'b111111111;
assign micromatrizz[98][379] = 9'b111111111;
assign micromatrizz[98][380] = 9'b111111111;
assign micromatrizz[98][381] = 9'b111111111;
assign micromatrizz[98][382] = 9'b111111111;
assign micromatrizz[98][383] = 9'b111111111;
assign micromatrizz[98][384] = 9'b111111111;
assign micromatrizz[98][385] = 9'b111111111;
assign micromatrizz[98][386] = 9'b111111111;
assign micromatrizz[98][387] = 9'b111111111;
assign micromatrizz[98][388] = 9'b111111111;
assign micromatrizz[98][389] = 9'b111111111;
assign micromatrizz[98][390] = 9'b111111111;
assign micromatrizz[98][391] = 9'b111111111;
assign micromatrizz[98][392] = 9'b111111111;
assign micromatrizz[98][393] = 9'b111111111;
assign micromatrizz[98][394] = 9'b111111111;
assign micromatrizz[98][395] = 9'b111111111;
assign micromatrizz[98][396] = 9'b111111111;
assign micromatrizz[98][397] = 9'b111111111;
assign micromatrizz[98][398] = 9'b111111111;
assign micromatrizz[98][399] = 9'b111111111;
assign micromatrizz[98][400] = 9'b111111111;
assign micromatrizz[98][401] = 9'b111111111;
assign micromatrizz[98][402] = 9'b111111111;
assign micromatrizz[98][403] = 9'b111111111;
assign micromatrizz[98][404] = 9'b111111111;
assign micromatrizz[98][405] = 9'b111111111;
assign micromatrizz[98][406] = 9'b111111111;
assign micromatrizz[98][407] = 9'b111111111;
assign micromatrizz[98][408] = 9'b111111111;
assign micromatrizz[98][409] = 9'b111111111;
assign micromatrizz[98][410] = 9'b111111111;
assign micromatrizz[98][411] = 9'b111111111;
assign micromatrizz[98][412] = 9'b111111111;
assign micromatrizz[98][413] = 9'b111111111;
assign micromatrizz[98][414] = 9'b111111111;
assign micromatrizz[98][415] = 9'b111111111;
assign micromatrizz[98][416] = 9'b111111111;
assign micromatrizz[98][417] = 9'b111111111;
assign micromatrizz[98][418] = 9'b111111111;
assign micromatrizz[98][419] = 9'b111111111;
assign micromatrizz[98][420] = 9'b111111111;
assign micromatrizz[98][421] = 9'b111111111;
assign micromatrizz[98][422] = 9'b111111111;
assign micromatrizz[98][423] = 9'b111111111;
assign micromatrizz[98][424] = 9'b111111111;
assign micromatrizz[98][425] = 9'b111111111;
assign micromatrizz[98][426] = 9'b111111111;
assign micromatrizz[98][427] = 9'b111111111;
assign micromatrizz[98][428] = 9'b111111111;
assign micromatrizz[98][429] = 9'b111111111;
assign micromatrizz[98][430] = 9'b111111111;
assign micromatrizz[98][431] = 9'b111111111;
assign micromatrizz[98][432] = 9'b111111111;
assign micromatrizz[98][433] = 9'b111111111;
assign micromatrizz[98][434] = 9'b111111111;
assign micromatrizz[98][435] = 9'b111111111;
assign micromatrizz[98][436] = 9'b111111111;
assign micromatrizz[98][437] = 9'b111111111;
assign micromatrizz[98][438] = 9'b111111111;
assign micromatrizz[98][439] = 9'b111111111;
assign micromatrizz[98][440] = 9'b111111111;
assign micromatrizz[98][441] = 9'b111111111;
assign micromatrizz[98][442] = 9'b111111111;
assign micromatrizz[98][443] = 9'b111111111;
assign micromatrizz[98][444] = 9'b111111111;
assign micromatrizz[98][445] = 9'b111111111;
assign micromatrizz[98][446] = 9'b111111111;
assign micromatrizz[98][447] = 9'b111111111;
assign micromatrizz[98][448] = 9'b111111111;
assign micromatrizz[98][449] = 9'b111111111;
assign micromatrizz[98][450] = 9'b111111111;
assign micromatrizz[98][451] = 9'b111111111;
assign micromatrizz[98][452] = 9'b111111111;
assign micromatrizz[98][453] = 9'b111111111;
assign micromatrizz[98][454] = 9'b111111111;
assign micromatrizz[98][455] = 9'b111111111;
assign micromatrizz[98][456] = 9'b111111111;
assign micromatrizz[98][457] = 9'b111111111;
assign micromatrizz[98][458] = 9'b111111111;
assign micromatrizz[98][459] = 9'b111111111;
assign micromatrizz[98][460] = 9'b111111111;
assign micromatrizz[98][461] = 9'b111111111;
assign micromatrizz[98][462] = 9'b111111111;
assign micromatrizz[98][463] = 9'b111111111;
assign micromatrizz[98][464] = 9'b111111111;
assign micromatrizz[98][465] = 9'b111111111;
assign micromatrizz[98][466] = 9'b111111111;
assign micromatrizz[98][467] = 9'b111111111;
assign micromatrizz[98][468] = 9'b111111111;
assign micromatrizz[98][469] = 9'b111111111;
assign micromatrizz[98][470] = 9'b111111111;
assign micromatrizz[98][471] = 9'b111111111;
assign micromatrizz[98][472] = 9'b111111111;
assign micromatrizz[98][473] = 9'b111111111;
assign micromatrizz[98][474] = 9'b111111111;
assign micromatrizz[98][475] = 9'b111111111;
assign micromatrizz[98][476] = 9'b111111111;
assign micromatrizz[98][477] = 9'b111111111;
assign micromatrizz[98][478] = 9'b111111111;
assign micromatrizz[98][479] = 9'b111111111;
assign micromatrizz[98][480] = 9'b111111111;
assign micromatrizz[98][481] = 9'b111111111;
assign micromatrizz[98][482] = 9'b111111111;
assign micromatrizz[98][483] = 9'b111111111;
assign micromatrizz[98][484] = 9'b111111111;
assign micromatrizz[98][485] = 9'b111111111;
assign micromatrizz[98][486] = 9'b111111111;
assign micromatrizz[98][487] = 9'b111111111;
assign micromatrizz[98][488] = 9'b111111111;
assign micromatrizz[98][489] = 9'b111111111;
assign micromatrizz[98][490] = 9'b111111111;
assign micromatrizz[98][491] = 9'b111111111;
assign micromatrizz[98][492] = 9'b111111111;
assign micromatrizz[98][493] = 9'b111111111;
assign micromatrizz[98][494] = 9'b111111111;
assign micromatrizz[98][495] = 9'b111111111;
assign micromatrizz[98][496] = 9'b111111111;
assign micromatrizz[98][497] = 9'b111111111;
assign micromatrizz[98][498] = 9'b111111111;
assign micromatrizz[98][499] = 9'b111111111;
assign micromatrizz[98][500] = 9'b111111111;
assign micromatrizz[98][501] = 9'b111111111;
assign micromatrizz[98][502] = 9'b111111111;
assign micromatrizz[98][503] = 9'b111111111;
assign micromatrizz[98][504] = 9'b111111111;
assign micromatrizz[98][505] = 9'b111111111;
assign micromatrizz[98][506] = 9'b111111111;
assign micromatrizz[98][507] = 9'b111111111;
assign micromatrizz[98][508] = 9'b111111111;
assign micromatrizz[98][509] = 9'b111111111;
assign micromatrizz[98][510] = 9'b111111111;
assign micromatrizz[98][511] = 9'b111111111;
assign micromatrizz[98][512] = 9'b111111111;
assign micromatrizz[98][513] = 9'b111111111;
assign micromatrizz[98][514] = 9'b111111111;
assign micromatrizz[98][515] = 9'b111111111;
assign micromatrizz[98][516] = 9'b111111111;
assign micromatrizz[98][517] = 9'b111111111;
assign micromatrizz[98][518] = 9'b111111111;
assign micromatrizz[98][519] = 9'b111111111;
assign micromatrizz[98][520] = 9'b111111111;
assign micromatrizz[98][521] = 9'b111111111;
assign micromatrizz[98][522] = 9'b111111111;
assign micromatrizz[98][523] = 9'b111111111;
assign micromatrizz[98][524] = 9'b111111111;
assign micromatrizz[98][525] = 9'b111111111;
assign micromatrizz[98][526] = 9'b111111111;
assign micromatrizz[98][527] = 9'b111111111;
assign micromatrizz[98][528] = 9'b111111111;
assign micromatrizz[98][529] = 9'b111111111;
assign micromatrizz[98][530] = 9'b111111111;
assign micromatrizz[98][531] = 9'b111111111;
assign micromatrizz[98][532] = 9'b111111111;
assign micromatrizz[98][533] = 9'b111111111;
assign micromatrizz[98][534] = 9'b111111111;
assign micromatrizz[98][535] = 9'b111111111;
assign micromatrizz[98][536] = 9'b111111111;
assign micromatrizz[98][537] = 9'b111111111;
assign micromatrizz[98][538] = 9'b111111111;
assign micromatrizz[98][539] = 9'b111111111;
assign micromatrizz[98][540] = 9'b111111111;
assign micromatrizz[98][541] = 9'b111111111;
assign micromatrizz[98][542] = 9'b111111111;
assign micromatrizz[98][543] = 9'b111111111;
assign micromatrizz[98][544] = 9'b111111111;
assign micromatrizz[98][545] = 9'b111111111;
assign micromatrizz[98][546] = 9'b111111111;
assign micromatrizz[98][547] = 9'b111111111;
assign micromatrizz[98][548] = 9'b111111111;
assign micromatrizz[98][549] = 9'b111111111;
assign micromatrizz[98][550] = 9'b111111111;
assign micromatrizz[98][551] = 9'b111111111;
assign micromatrizz[98][552] = 9'b111111111;
assign micromatrizz[98][553] = 9'b111111111;
assign micromatrizz[98][554] = 9'b111111111;
assign micromatrizz[98][555] = 9'b111111111;
assign micromatrizz[98][556] = 9'b111111111;
assign micromatrizz[98][557] = 9'b111111111;
assign micromatrizz[98][558] = 9'b111111111;
assign micromatrizz[98][559] = 9'b111111111;
assign micromatrizz[98][560] = 9'b111111111;
assign micromatrizz[98][561] = 9'b111111111;
assign micromatrizz[98][562] = 9'b111111111;
assign micromatrizz[98][563] = 9'b111111111;
assign micromatrizz[98][564] = 9'b111111111;
assign micromatrizz[98][565] = 9'b111111111;
assign micromatrizz[98][566] = 9'b111111111;
assign micromatrizz[98][567] = 9'b111111111;
assign micromatrizz[98][568] = 9'b111111111;
assign micromatrizz[98][569] = 9'b111111111;
assign micromatrizz[98][570] = 9'b111111111;
assign micromatrizz[98][571] = 9'b111111111;
assign micromatrizz[98][572] = 9'b111111111;
assign micromatrizz[98][573] = 9'b111111111;
assign micromatrizz[98][574] = 9'b111111111;
assign micromatrizz[98][575] = 9'b111111111;
assign micromatrizz[98][576] = 9'b111111111;
assign micromatrizz[98][577] = 9'b111111111;
assign micromatrizz[98][578] = 9'b111111111;
assign micromatrizz[98][579] = 9'b111111111;
assign micromatrizz[98][580] = 9'b111111111;
assign micromatrizz[98][581] = 9'b111111111;
assign micromatrizz[98][582] = 9'b111111111;
assign micromatrizz[98][583] = 9'b111111111;
assign micromatrizz[98][584] = 9'b111111111;
assign micromatrizz[98][585] = 9'b111111111;
assign micromatrizz[98][586] = 9'b111111111;
assign micromatrizz[98][587] = 9'b111111111;
assign micromatrizz[98][588] = 9'b111111111;
assign micromatrizz[98][589] = 9'b111111111;
assign micromatrizz[98][590] = 9'b111111111;
assign micromatrizz[98][591] = 9'b111111111;
assign micromatrizz[98][592] = 9'b111111111;
assign micromatrizz[98][593] = 9'b111111111;
assign micromatrizz[98][594] = 9'b111111111;
assign micromatrizz[98][595] = 9'b111111111;
assign micromatrizz[98][596] = 9'b111111111;
assign micromatrizz[98][597] = 9'b111111111;
assign micromatrizz[98][598] = 9'b111111111;
assign micromatrizz[98][599] = 9'b111111111;
assign micromatrizz[98][600] = 9'b111111111;
assign micromatrizz[98][601] = 9'b111111111;
assign micromatrizz[98][602] = 9'b111111111;
assign micromatrizz[98][603] = 9'b111111111;
assign micromatrizz[98][604] = 9'b111111111;
assign micromatrizz[98][605] = 9'b111111111;
assign micromatrizz[98][606] = 9'b111111111;
assign micromatrizz[98][607] = 9'b111111111;
assign micromatrizz[98][608] = 9'b111111111;
assign micromatrizz[98][609] = 9'b111111111;
assign micromatrizz[98][610] = 9'b111111111;
assign micromatrizz[98][611] = 9'b111111111;
assign micromatrizz[98][612] = 9'b111111111;
assign micromatrizz[98][613] = 9'b111111111;
assign micromatrizz[98][614] = 9'b111111111;
assign micromatrizz[98][615] = 9'b111111111;
assign micromatrizz[98][616] = 9'b111111111;
assign micromatrizz[98][617] = 9'b111111111;
assign micromatrizz[98][618] = 9'b111111111;
assign micromatrizz[98][619] = 9'b111111111;
assign micromatrizz[98][620] = 9'b111111111;
assign micromatrizz[98][621] = 9'b111111111;
assign micromatrizz[98][622] = 9'b111111111;
assign micromatrizz[98][623] = 9'b111111111;
assign micromatrizz[98][624] = 9'b111111111;
assign micromatrizz[98][625] = 9'b111111111;
assign micromatrizz[98][626] = 9'b111111111;
assign micromatrizz[98][627] = 9'b111111111;
assign micromatrizz[98][628] = 9'b111111111;
assign micromatrizz[98][629] = 9'b111111111;
assign micromatrizz[98][630] = 9'b111111111;
assign micromatrizz[98][631] = 9'b111111111;
assign micromatrizz[98][632] = 9'b111111111;
assign micromatrizz[98][633] = 9'b111111111;
assign micromatrizz[98][634] = 9'b111111111;
assign micromatrizz[98][635] = 9'b111111111;
assign micromatrizz[98][636] = 9'b111111111;
assign micromatrizz[98][637] = 9'b111111111;
assign micromatrizz[98][638] = 9'b111111111;
assign micromatrizz[98][639] = 9'b111111111;
assign micromatrizz[99][0] = 9'b111111111;
assign micromatrizz[99][1] = 9'b111111111;
assign micromatrizz[99][2] = 9'b111111111;
assign micromatrizz[99][3] = 9'b111111111;
assign micromatrizz[99][4] = 9'b111111111;
assign micromatrizz[99][5] = 9'b111111111;
assign micromatrizz[99][6] = 9'b111111111;
assign micromatrizz[99][7] = 9'b111111111;
assign micromatrizz[99][8] = 9'b111111111;
assign micromatrizz[99][9] = 9'b111111111;
assign micromatrizz[99][10] = 9'b111111111;
assign micromatrizz[99][11] = 9'b111111111;
assign micromatrizz[99][12] = 9'b111111111;
assign micromatrizz[99][13] = 9'b111111111;
assign micromatrizz[99][14] = 9'b111111111;
assign micromatrizz[99][15] = 9'b111111111;
assign micromatrizz[99][16] = 9'b111111111;
assign micromatrizz[99][17] = 9'b111111111;
assign micromatrizz[99][18] = 9'b111111111;
assign micromatrizz[99][19] = 9'b111111111;
assign micromatrizz[99][20] = 9'b111111111;
assign micromatrizz[99][21] = 9'b111111111;
assign micromatrizz[99][22] = 9'b111111111;
assign micromatrizz[99][23] = 9'b111111111;
assign micromatrizz[99][24] = 9'b111111111;
assign micromatrizz[99][25] = 9'b111111111;
assign micromatrizz[99][26] = 9'b111111111;
assign micromatrizz[99][27] = 9'b111111111;
assign micromatrizz[99][28] = 9'b111111111;
assign micromatrizz[99][29] = 9'b111111111;
assign micromatrizz[99][30] = 9'b111111111;
assign micromatrizz[99][31] = 9'b111111111;
assign micromatrizz[99][32] = 9'b111111111;
assign micromatrizz[99][33] = 9'b111111111;
assign micromatrizz[99][34] = 9'b111111111;
assign micromatrizz[99][35] = 9'b111111111;
assign micromatrizz[99][36] = 9'b111111111;
assign micromatrizz[99][37] = 9'b111111111;
assign micromatrizz[99][38] = 9'b111111111;
assign micromatrizz[99][39] = 9'b111111111;
assign micromatrizz[99][40] = 9'b111111111;
assign micromatrizz[99][41] = 9'b111111111;
assign micromatrizz[99][42] = 9'b111111111;
assign micromatrizz[99][43] = 9'b111111111;
assign micromatrizz[99][44] = 9'b111111111;
assign micromatrizz[99][45] = 9'b111111111;
assign micromatrizz[99][46] = 9'b111111111;
assign micromatrizz[99][47] = 9'b111111111;
assign micromatrizz[99][48] = 9'b111111111;
assign micromatrizz[99][49] = 9'b111111111;
assign micromatrizz[99][50] = 9'b111111111;
assign micromatrizz[99][51] = 9'b111111111;
assign micromatrizz[99][52] = 9'b111111111;
assign micromatrizz[99][53] = 9'b111111111;
assign micromatrizz[99][54] = 9'b111111111;
assign micromatrizz[99][55] = 9'b111111111;
assign micromatrizz[99][56] = 9'b111111111;
assign micromatrizz[99][57] = 9'b111111111;
assign micromatrizz[99][58] = 9'b111111111;
assign micromatrizz[99][59] = 9'b111111111;
assign micromatrizz[99][60] = 9'b111111111;
assign micromatrizz[99][61] = 9'b111111111;
assign micromatrizz[99][62] = 9'b111111111;
assign micromatrizz[99][63] = 9'b111111111;
assign micromatrizz[99][64] = 9'b111111111;
assign micromatrizz[99][65] = 9'b111111111;
assign micromatrizz[99][66] = 9'b111111111;
assign micromatrizz[99][67] = 9'b111111111;
assign micromatrizz[99][68] = 9'b111111111;
assign micromatrizz[99][69] = 9'b111111111;
assign micromatrizz[99][70] = 9'b111111111;
assign micromatrizz[99][71] = 9'b111111111;
assign micromatrizz[99][72] = 9'b111111111;
assign micromatrizz[99][73] = 9'b111111111;
assign micromatrizz[99][74] = 9'b111111111;
assign micromatrizz[99][75] = 9'b111111111;
assign micromatrizz[99][76] = 9'b111111111;
assign micromatrizz[99][77] = 9'b111111111;
assign micromatrizz[99][78] = 9'b111111111;
assign micromatrizz[99][79] = 9'b111111111;
assign micromatrizz[99][80] = 9'b111111111;
assign micromatrizz[99][81] = 9'b111111111;
assign micromatrizz[99][82] = 9'b111111111;
assign micromatrizz[99][83] = 9'b111111111;
assign micromatrizz[99][84] = 9'b111111111;
assign micromatrizz[99][85] = 9'b111111111;
assign micromatrizz[99][86] = 9'b111111111;
assign micromatrizz[99][87] = 9'b111111111;
assign micromatrizz[99][88] = 9'b111111111;
assign micromatrizz[99][89] = 9'b111111111;
assign micromatrizz[99][90] = 9'b111111111;
assign micromatrizz[99][91] = 9'b111111111;
assign micromatrizz[99][92] = 9'b111111111;
assign micromatrizz[99][93] = 9'b111111111;
assign micromatrizz[99][94] = 9'b111111111;
assign micromatrizz[99][95] = 9'b111111111;
assign micromatrizz[99][96] = 9'b111111111;
assign micromatrizz[99][97] = 9'b111111111;
assign micromatrizz[99][98] = 9'b111111111;
assign micromatrizz[99][99] = 9'b111111111;
assign micromatrizz[99][100] = 9'b111111111;
assign micromatrizz[99][101] = 9'b111111111;
assign micromatrizz[99][102] = 9'b111111111;
assign micromatrizz[99][103] = 9'b111111111;
assign micromatrizz[99][104] = 9'b111111111;
assign micromatrizz[99][105] = 9'b111111111;
assign micromatrizz[99][106] = 9'b111111111;
assign micromatrizz[99][107] = 9'b111111111;
assign micromatrizz[99][108] = 9'b111111111;
assign micromatrizz[99][109] = 9'b111111111;
assign micromatrizz[99][110] = 9'b111111111;
assign micromatrizz[99][111] = 9'b111111111;
assign micromatrizz[99][112] = 9'b111111111;
assign micromatrizz[99][113] = 9'b111111111;
assign micromatrizz[99][114] = 9'b111111111;
assign micromatrizz[99][115] = 9'b111111111;
assign micromatrizz[99][116] = 9'b111111111;
assign micromatrizz[99][117] = 9'b111111111;
assign micromatrizz[99][118] = 9'b111111111;
assign micromatrizz[99][119] = 9'b111111111;
assign micromatrizz[99][120] = 9'b111111111;
assign micromatrizz[99][121] = 9'b111111111;
assign micromatrizz[99][122] = 9'b111111111;
assign micromatrizz[99][123] = 9'b111111111;
assign micromatrizz[99][124] = 9'b111111111;
assign micromatrizz[99][125] = 9'b111111111;
assign micromatrizz[99][126] = 9'b111111111;
assign micromatrizz[99][127] = 9'b111111111;
assign micromatrizz[99][128] = 9'b111111111;
assign micromatrizz[99][129] = 9'b111111111;
assign micromatrizz[99][130] = 9'b111111111;
assign micromatrizz[99][131] = 9'b111111111;
assign micromatrizz[99][132] = 9'b111111111;
assign micromatrizz[99][133] = 9'b111111111;
assign micromatrizz[99][134] = 9'b111111111;
assign micromatrizz[99][135] = 9'b111111111;
assign micromatrizz[99][136] = 9'b111111111;
assign micromatrizz[99][137] = 9'b111111111;
assign micromatrizz[99][138] = 9'b111111111;
assign micromatrizz[99][139] = 9'b111111111;
assign micromatrizz[99][140] = 9'b111111111;
assign micromatrizz[99][141] = 9'b111111111;
assign micromatrizz[99][142] = 9'b111111111;
assign micromatrizz[99][143] = 9'b111111111;
assign micromatrizz[99][144] = 9'b111111111;
assign micromatrizz[99][145] = 9'b111111111;
assign micromatrizz[99][146] = 9'b111111111;
assign micromatrizz[99][147] = 9'b111111111;
assign micromatrizz[99][148] = 9'b111111111;
assign micromatrizz[99][149] = 9'b111111111;
assign micromatrizz[99][150] = 9'b111111111;
assign micromatrizz[99][151] = 9'b111111111;
assign micromatrizz[99][152] = 9'b111111111;
assign micromatrizz[99][153] = 9'b111111111;
assign micromatrizz[99][154] = 9'b111111111;
assign micromatrizz[99][155] = 9'b111111111;
assign micromatrizz[99][156] = 9'b111111111;
assign micromatrizz[99][157] = 9'b111111111;
assign micromatrizz[99][158] = 9'b111111111;
assign micromatrizz[99][159] = 9'b111111111;
assign micromatrizz[99][160] = 9'b111111111;
assign micromatrizz[99][161] = 9'b111111111;
assign micromatrizz[99][162] = 9'b111111111;
assign micromatrizz[99][163] = 9'b111111111;
assign micromatrizz[99][164] = 9'b111111111;
assign micromatrizz[99][165] = 9'b111111111;
assign micromatrizz[99][166] = 9'b111111111;
assign micromatrizz[99][167] = 9'b111111111;
assign micromatrizz[99][168] = 9'b111111111;
assign micromatrizz[99][169] = 9'b111111111;
assign micromatrizz[99][170] = 9'b111111111;
assign micromatrizz[99][171] = 9'b111111111;
assign micromatrizz[99][172] = 9'b111111111;
assign micromatrizz[99][173] = 9'b111111111;
assign micromatrizz[99][174] = 9'b111111111;
assign micromatrizz[99][175] = 9'b111111111;
assign micromatrizz[99][176] = 9'b111111111;
assign micromatrizz[99][177] = 9'b111111111;
assign micromatrizz[99][178] = 9'b111111111;
assign micromatrizz[99][179] = 9'b111111111;
assign micromatrizz[99][180] = 9'b111111111;
assign micromatrizz[99][181] = 9'b111111111;
assign micromatrizz[99][182] = 9'b111111111;
assign micromatrizz[99][183] = 9'b111111111;
assign micromatrizz[99][184] = 9'b111111111;
assign micromatrizz[99][185] = 9'b111111111;
assign micromatrizz[99][186] = 9'b111111111;
assign micromatrizz[99][187] = 9'b111111111;
assign micromatrizz[99][188] = 9'b111111111;
assign micromatrizz[99][189] = 9'b111111111;
assign micromatrizz[99][190] = 9'b111111111;
assign micromatrizz[99][191] = 9'b111111111;
assign micromatrizz[99][192] = 9'b111111111;
assign micromatrizz[99][193] = 9'b111111111;
assign micromatrizz[99][194] = 9'b111111111;
assign micromatrizz[99][195] = 9'b111111111;
assign micromatrizz[99][196] = 9'b111111111;
assign micromatrizz[99][197] = 9'b111111111;
assign micromatrizz[99][198] = 9'b111111111;
assign micromatrizz[99][199] = 9'b111111111;
assign micromatrizz[99][200] = 9'b111111111;
assign micromatrizz[99][201] = 9'b111111111;
assign micromatrizz[99][202] = 9'b111111111;
assign micromatrizz[99][203] = 9'b111111111;
assign micromatrizz[99][204] = 9'b111111111;
assign micromatrizz[99][205] = 9'b111111111;
assign micromatrizz[99][206] = 9'b111111111;
assign micromatrizz[99][207] = 9'b111111111;
assign micromatrizz[99][208] = 9'b111111111;
assign micromatrizz[99][209] = 9'b111111111;
assign micromatrizz[99][210] = 9'b111111111;
assign micromatrizz[99][211] = 9'b111111111;
assign micromatrizz[99][212] = 9'b111111111;
assign micromatrizz[99][213] = 9'b111111111;
assign micromatrizz[99][214] = 9'b111111111;
assign micromatrizz[99][215] = 9'b111111111;
assign micromatrizz[99][216] = 9'b111111111;
assign micromatrizz[99][217] = 9'b111111111;
assign micromatrizz[99][218] = 9'b111111111;
assign micromatrizz[99][219] = 9'b111111111;
assign micromatrizz[99][220] = 9'b111111111;
assign micromatrizz[99][221] = 9'b111111111;
assign micromatrizz[99][222] = 9'b111111111;
assign micromatrizz[99][223] = 9'b111111111;
assign micromatrizz[99][224] = 9'b111111111;
assign micromatrizz[99][225] = 9'b111111111;
assign micromatrizz[99][226] = 9'b111111111;
assign micromatrizz[99][227] = 9'b111111111;
assign micromatrizz[99][228] = 9'b111111111;
assign micromatrizz[99][229] = 9'b111111111;
assign micromatrizz[99][230] = 9'b111111111;
assign micromatrizz[99][231] = 9'b111111111;
assign micromatrizz[99][232] = 9'b111111111;
assign micromatrizz[99][233] = 9'b111111111;
assign micromatrizz[99][234] = 9'b111111111;
assign micromatrizz[99][235] = 9'b111111111;
assign micromatrizz[99][236] = 9'b111111111;
assign micromatrizz[99][237] = 9'b111111111;
assign micromatrizz[99][238] = 9'b111111111;
assign micromatrizz[99][239] = 9'b111111111;
assign micromatrizz[99][240] = 9'b111111111;
assign micromatrizz[99][241] = 9'b111111111;
assign micromatrizz[99][242] = 9'b111111111;
assign micromatrizz[99][243] = 9'b111111111;
assign micromatrizz[99][244] = 9'b111111111;
assign micromatrizz[99][245] = 9'b111111111;
assign micromatrizz[99][246] = 9'b111111111;
assign micromatrizz[99][247] = 9'b111111111;
assign micromatrizz[99][248] = 9'b111111111;
assign micromatrizz[99][249] = 9'b111111111;
assign micromatrizz[99][250] = 9'b111111111;
assign micromatrizz[99][251] = 9'b111111111;
assign micromatrizz[99][252] = 9'b111111111;
assign micromatrizz[99][253] = 9'b111111111;
assign micromatrizz[99][254] = 9'b111111111;
assign micromatrizz[99][255] = 9'b111111111;
assign micromatrizz[99][256] = 9'b111111111;
assign micromatrizz[99][257] = 9'b111111111;
assign micromatrizz[99][258] = 9'b111111111;
assign micromatrizz[99][259] = 9'b111111111;
assign micromatrizz[99][260] = 9'b111111111;
assign micromatrizz[99][261] = 9'b111111111;
assign micromatrizz[99][262] = 9'b111111111;
assign micromatrizz[99][263] = 9'b111111111;
assign micromatrizz[99][264] = 9'b111111111;
assign micromatrizz[99][265] = 9'b111111111;
assign micromatrizz[99][266] = 9'b111111111;
assign micromatrizz[99][267] = 9'b111111111;
assign micromatrizz[99][268] = 9'b111111111;
assign micromatrizz[99][269] = 9'b111111111;
assign micromatrizz[99][270] = 9'b111111111;
assign micromatrizz[99][271] = 9'b111111111;
assign micromatrizz[99][272] = 9'b111111111;
assign micromatrizz[99][273] = 9'b111111111;
assign micromatrizz[99][274] = 9'b111111111;
assign micromatrizz[99][275] = 9'b111111111;
assign micromatrizz[99][276] = 9'b111111111;
assign micromatrizz[99][277] = 9'b111111111;
assign micromatrizz[99][278] = 9'b111111111;
assign micromatrizz[99][279] = 9'b111111111;
assign micromatrizz[99][280] = 9'b111111111;
assign micromatrizz[99][281] = 9'b111111111;
assign micromatrizz[99][282] = 9'b111111111;
assign micromatrizz[99][283] = 9'b111111111;
assign micromatrizz[99][284] = 9'b111111111;
assign micromatrizz[99][285] = 9'b111111111;
assign micromatrizz[99][286] = 9'b111111111;
assign micromatrizz[99][287] = 9'b111111111;
assign micromatrizz[99][288] = 9'b111111111;
assign micromatrizz[99][289] = 9'b111111111;
assign micromatrizz[99][290] = 9'b111111111;
assign micromatrizz[99][291] = 9'b111111111;
assign micromatrizz[99][292] = 9'b111111111;
assign micromatrizz[99][293] = 9'b111111111;
assign micromatrizz[99][294] = 9'b111111111;
assign micromatrizz[99][295] = 9'b111111111;
assign micromatrizz[99][296] = 9'b111111111;
assign micromatrizz[99][297] = 9'b111111111;
assign micromatrizz[99][298] = 9'b111111111;
assign micromatrizz[99][299] = 9'b111111111;
assign micromatrizz[99][300] = 9'b111111111;
assign micromatrizz[99][301] = 9'b111111111;
assign micromatrizz[99][302] = 9'b111111111;
assign micromatrizz[99][303] = 9'b111111111;
assign micromatrizz[99][304] = 9'b111111111;
assign micromatrizz[99][305] = 9'b111111111;
assign micromatrizz[99][306] = 9'b111111111;
assign micromatrizz[99][307] = 9'b111111111;
assign micromatrizz[99][308] = 9'b111111111;
assign micromatrizz[99][309] = 9'b111111111;
assign micromatrizz[99][310] = 9'b111111111;
assign micromatrizz[99][311] = 9'b111111111;
assign micromatrizz[99][312] = 9'b111111111;
assign micromatrizz[99][313] = 9'b111111111;
assign micromatrizz[99][314] = 9'b111111111;
assign micromatrizz[99][315] = 9'b111111111;
assign micromatrizz[99][316] = 9'b111111111;
assign micromatrizz[99][317] = 9'b111111111;
assign micromatrizz[99][318] = 9'b111111111;
assign micromatrizz[99][319] = 9'b111111111;
assign micromatrizz[99][320] = 9'b111111111;
assign micromatrizz[99][321] = 9'b111111111;
assign micromatrizz[99][322] = 9'b111111111;
assign micromatrizz[99][323] = 9'b111111111;
assign micromatrizz[99][324] = 9'b111111111;
assign micromatrizz[99][325] = 9'b111111111;
assign micromatrizz[99][326] = 9'b111111111;
assign micromatrizz[99][327] = 9'b111111111;
assign micromatrizz[99][328] = 9'b111111111;
assign micromatrizz[99][329] = 9'b111111111;
assign micromatrizz[99][330] = 9'b111111111;
assign micromatrizz[99][331] = 9'b111111111;
assign micromatrizz[99][332] = 9'b111111111;
assign micromatrizz[99][333] = 9'b111111111;
assign micromatrizz[99][334] = 9'b111111111;
assign micromatrizz[99][335] = 9'b111111111;
assign micromatrizz[99][336] = 9'b111111111;
assign micromatrizz[99][337] = 9'b111111111;
assign micromatrizz[99][338] = 9'b111111111;
assign micromatrizz[99][339] = 9'b111111111;
assign micromatrizz[99][340] = 9'b111111111;
assign micromatrizz[99][341] = 9'b111111111;
assign micromatrizz[99][342] = 9'b111111111;
assign micromatrizz[99][343] = 9'b111111111;
assign micromatrizz[99][344] = 9'b111111111;
assign micromatrizz[99][345] = 9'b111111111;
assign micromatrizz[99][346] = 9'b111111111;
assign micromatrizz[99][347] = 9'b111111111;
assign micromatrizz[99][348] = 9'b111111111;
assign micromatrizz[99][349] = 9'b111111111;
assign micromatrizz[99][350] = 9'b111111111;
assign micromatrizz[99][351] = 9'b111111111;
assign micromatrizz[99][352] = 9'b111111111;
assign micromatrizz[99][353] = 9'b111111111;
assign micromatrizz[99][354] = 9'b111111111;
assign micromatrizz[99][355] = 9'b111111111;
assign micromatrizz[99][356] = 9'b111111111;
assign micromatrizz[99][357] = 9'b111111111;
assign micromatrizz[99][358] = 9'b111111111;
assign micromatrizz[99][359] = 9'b111111111;
assign micromatrizz[99][360] = 9'b111111111;
assign micromatrizz[99][361] = 9'b111111111;
assign micromatrizz[99][362] = 9'b111111111;
assign micromatrizz[99][363] = 9'b111111111;
assign micromatrizz[99][364] = 9'b111111111;
assign micromatrizz[99][365] = 9'b111111111;
assign micromatrizz[99][366] = 9'b111111111;
assign micromatrizz[99][367] = 9'b111111111;
assign micromatrizz[99][368] = 9'b111111111;
assign micromatrizz[99][369] = 9'b111111111;
assign micromatrizz[99][370] = 9'b111111111;
assign micromatrizz[99][371] = 9'b111111111;
assign micromatrizz[99][372] = 9'b111111111;
assign micromatrizz[99][373] = 9'b111111111;
assign micromatrizz[99][374] = 9'b111111111;
assign micromatrizz[99][375] = 9'b111111111;
assign micromatrizz[99][376] = 9'b111111111;
assign micromatrizz[99][377] = 9'b111111111;
assign micromatrizz[99][378] = 9'b111111111;
assign micromatrizz[99][379] = 9'b111111111;
assign micromatrizz[99][380] = 9'b111111111;
assign micromatrizz[99][381] = 9'b111111111;
assign micromatrizz[99][382] = 9'b111111111;
assign micromatrizz[99][383] = 9'b111111111;
assign micromatrizz[99][384] = 9'b111111111;
assign micromatrizz[99][385] = 9'b111111111;
assign micromatrizz[99][386] = 9'b111111111;
assign micromatrizz[99][387] = 9'b111111111;
assign micromatrizz[99][388] = 9'b111111111;
assign micromatrizz[99][389] = 9'b111111111;
assign micromatrizz[99][390] = 9'b111111111;
assign micromatrizz[99][391] = 9'b111111111;
assign micromatrizz[99][392] = 9'b111111111;
assign micromatrizz[99][393] = 9'b111111111;
assign micromatrizz[99][394] = 9'b111111111;
assign micromatrizz[99][395] = 9'b111111111;
assign micromatrizz[99][396] = 9'b111111111;
assign micromatrizz[99][397] = 9'b111111111;
assign micromatrizz[99][398] = 9'b111111111;
assign micromatrizz[99][399] = 9'b111111111;
assign micromatrizz[99][400] = 9'b111111111;
assign micromatrizz[99][401] = 9'b111111111;
assign micromatrizz[99][402] = 9'b111111111;
assign micromatrizz[99][403] = 9'b111111111;
assign micromatrizz[99][404] = 9'b111111111;
assign micromatrizz[99][405] = 9'b111111111;
assign micromatrizz[99][406] = 9'b111111111;
assign micromatrizz[99][407] = 9'b111111111;
assign micromatrizz[99][408] = 9'b111111111;
assign micromatrizz[99][409] = 9'b111111111;
assign micromatrizz[99][410] = 9'b111111111;
assign micromatrizz[99][411] = 9'b111111111;
assign micromatrizz[99][412] = 9'b111111111;
assign micromatrizz[99][413] = 9'b111111111;
assign micromatrizz[99][414] = 9'b111111111;
assign micromatrizz[99][415] = 9'b111111111;
assign micromatrizz[99][416] = 9'b111111111;
assign micromatrizz[99][417] = 9'b111111111;
assign micromatrizz[99][418] = 9'b111111111;
assign micromatrizz[99][419] = 9'b111111111;
assign micromatrizz[99][420] = 9'b111111111;
assign micromatrizz[99][421] = 9'b111111111;
assign micromatrizz[99][422] = 9'b111111111;
assign micromatrizz[99][423] = 9'b111111111;
assign micromatrizz[99][424] = 9'b111111111;
assign micromatrizz[99][425] = 9'b111111111;
assign micromatrizz[99][426] = 9'b111111111;
assign micromatrizz[99][427] = 9'b111111111;
assign micromatrizz[99][428] = 9'b111111111;
assign micromatrizz[99][429] = 9'b111111111;
assign micromatrizz[99][430] = 9'b111111111;
assign micromatrizz[99][431] = 9'b111111111;
assign micromatrizz[99][432] = 9'b111111111;
assign micromatrizz[99][433] = 9'b111111111;
assign micromatrizz[99][434] = 9'b111111111;
assign micromatrizz[99][435] = 9'b111111111;
assign micromatrizz[99][436] = 9'b111111111;
assign micromatrizz[99][437] = 9'b111111111;
assign micromatrizz[99][438] = 9'b111111111;
assign micromatrizz[99][439] = 9'b111111111;
assign micromatrizz[99][440] = 9'b111111111;
assign micromatrizz[99][441] = 9'b111111111;
assign micromatrizz[99][442] = 9'b111111111;
assign micromatrizz[99][443] = 9'b111111111;
assign micromatrizz[99][444] = 9'b111111111;
assign micromatrizz[99][445] = 9'b111111111;
assign micromatrizz[99][446] = 9'b111111111;
assign micromatrizz[99][447] = 9'b111111111;
assign micromatrizz[99][448] = 9'b111111111;
assign micromatrizz[99][449] = 9'b111111111;
assign micromatrizz[99][450] = 9'b111111111;
assign micromatrizz[99][451] = 9'b111111111;
assign micromatrizz[99][452] = 9'b111111111;
assign micromatrizz[99][453] = 9'b111111111;
assign micromatrizz[99][454] = 9'b111111111;
assign micromatrizz[99][455] = 9'b111111111;
assign micromatrizz[99][456] = 9'b111111111;
assign micromatrizz[99][457] = 9'b111111111;
assign micromatrizz[99][458] = 9'b111111111;
assign micromatrizz[99][459] = 9'b111111111;
assign micromatrizz[99][460] = 9'b111111111;
assign micromatrizz[99][461] = 9'b111111111;
assign micromatrizz[99][462] = 9'b111111111;
assign micromatrizz[99][463] = 9'b111111111;
assign micromatrizz[99][464] = 9'b111111111;
assign micromatrizz[99][465] = 9'b111111111;
assign micromatrizz[99][466] = 9'b111111111;
assign micromatrizz[99][467] = 9'b111111111;
assign micromatrizz[99][468] = 9'b111111111;
assign micromatrizz[99][469] = 9'b111111111;
assign micromatrizz[99][470] = 9'b111111111;
assign micromatrizz[99][471] = 9'b111111111;
assign micromatrizz[99][472] = 9'b111111111;
assign micromatrizz[99][473] = 9'b111111111;
assign micromatrizz[99][474] = 9'b111111111;
assign micromatrizz[99][475] = 9'b111111111;
assign micromatrizz[99][476] = 9'b111111111;
assign micromatrizz[99][477] = 9'b111111111;
assign micromatrizz[99][478] = 9'b111111111;
assign micromatrizz[99][479] = 9'b111111111;
assign micromatrizz[99][480] = 9'b111111111;
assign micromatrizz[99][481] = 9'b111111111;
assign micromatrizz[99][482] = 9'b111111111;
assign micromatrizz[99][483] = 9'b111111111;
assign micromatrizz[99][484] = 9'b111111111;
assign micromatrizz[99][485] = 9'b111111111;
assign micromatrizz[99][486] = 9'b111111111;
assign micromatrizz[99][487] = 9'b111111111;
assign micromatrizz[99][488] = 9'b111111111;
assign micromatrizz[99][489] = 9'b111111111;
assign micromatrizz[99][490] = 9'b111111111;
assign micromatrizz[99][491] = 9'b111111111;
assign micromatrizz[99][492] = 9'b111111111;
assign micromatrizz[99][493] = 9'b111111111;
assign micromatrizz[99][494] = 9'b111111111;
assign micromatrizz[99][495] = 9'b111111111;
assign micromatrizz[99][496] = 9'b111111111;
assign micromatrizz[99][497] = 9'b111111111;
assign micromatrizz[99][498] = 9'b111111111;
assign micromatrizz[99][499] = 9'b111111111;
assign micromatrizz[99][500] = 9'b111111111;
assign micromatrizz[99][501] = 9'b111111111;
assign micromatrizz[99][502] = 9'b111111111;
assign micromatrizz[99][503] = 9'b111111111;
assign micromatrizz[99][504] = 9'b111111111;
assign micromatrizz[99][505] = 9'b111111111;
assign micromatrizz[99][506] = 9'b111111111;
assign micromatrizz[99][507] = 9'b111111111;
assign micromatrizz[99][508] = 9'b111111111;
assign micromatrizz[99][509] = 9'b111111111;
assign micromatrizz[99][510] = 9'b111111111;
assign micromatrizz[99][511] = 9'b111111111;
assign micromatrizz[99][512] = 9'b111111111;
assign micromatrizz[99][513] = 9'b111111111;
assign micromatrizz[99][514] = 9'b111111111;
assign micromatrizz[99][515] = 9'b111111111;
assign micromatrizz[99][516] = 9'b111111111;
assign micromatrizz[99][517] = 9'b111111111;
assign micromatrizz[99][518] = 9'b111111111;
assign micromatrizz[99][519] = 9'b111111111;
assign micromatrizz[99][520] = 9'b111111111;
assign micromatrizz[99][521] = 9'b111111111;
assign micromatrizz[99][522] = 9'b111111111;
assign micromatrizz[99][523] = 9'b111111111;
assign micromatrizz[99][524] = 9'b111111111;
assign micromatrizz[99][525] = 9'b111111111;
assign micromatrizz[99][526] = 9'b111111111;
assign micromatrizz[99][527] = 9'b111111111;
assign micromatrizz[99][528] = 9'b111111111;
assign micromatrizz[99][529] = 9'b111111111;
assign micromatrizz[99][530] = 9'b111111111;
assign micromatrizz[99][531] = 9'b111111111;
assign micromatrizz[99][532] = 9'b111111111;
assign micromatrizz[99][533] = 9'b111111111;
assign micromatrizz[99][534] = 9'b111111111;
assign micromatrizz[99][535] = 9'b111111111;
assign micromatrizz[99][536] = 9'b111111111;
assign micromatrizz[99][537] = 9'b111111111;
assign micromatrizz[99][538] = 9'b111111111;
assign micromatrizz[99][539] = 9'b111111111;
assign micromatrizz[99][540] = 9'b111111111;
assign micromatrizz[99][541] = 9'b111111111;
assign micromatrizz[99][542] = 9'b111111111;
assign micromatrizz[99][543] = 9'b111111111;
assign micromatrizz[99][544] = 9'b111111111;
assign micromatrizz[99][545] = 9'b111111111;
assign micromatrizz[99][546] = 9'b111111111;
assign micromatrizz[99][547] = 9'b111111111;
assign micromatrizz[99][548] = 9'b111111111;
assign micromatrizz[99][549] = 9'b111111111;
assign micromatrizz[99][550] = 9'b111111111;
assign micromatrizz[99][551] = 9'b111111111;
assign micromatrizz[99][552] = 9'b111111111;
assign micromatrizz[99][553] = 9'b111111111;
assign micromatrizz[99][554] = 9'b111111111;
assign micromatrizz[99][555] = 9'b111111111;
assign micromatrizz[99][556] = 9'b111111111;
assign micromatrizz[99][557] = 9'b111111111;
assign micromatrizz[99][558] = 9'b111111111;
assign micromatrizz[99][559] = 9'b111111111;
assign micromatrizz[99][560] = 9'b111111111;
assign micromatrizz[99][561] = 9'b111111111;
assign micromatrizz[99][562] = 9'b111111111;
assign micromatrizz[99][563] = 9'b111111111;
assign micromatrizz[99][564] = 9'b111111111;
assign micromatrizz[99][565] = 9'b111111111;
assign micromatrizz[99][566] = 9'b111111111;
assign micromatrizz[99][567] = 9'b111111111;
assign micromatrizz[99][568] = 9'b111111111;
assign micromatrizz[99][569] = 9'b111111111;
assign micromatrizz[99][570] = 9'b111111111;
assign micromatrizz[99][571] = 9'b111111111;
assign micromatrizz[99][572] = 9'b111111111;
assign micromatrizz[99][573] = 9'b111111111;
assign micromatrizz[99][574] = 9'b111111111;
assign micromatrizz[99][575] = 9'b111111111;
assign micromatrizz[99][576] = 9'b111111111;
assign micromatrizz[99][577] = 9'b111111111;
assign micromatrizz[99][578] = 9'b111111111;
assign micromatrizz[99][579] = 9'b111111111;
assign micromatrizz[99][580] = 9'b111111111;
assign micromatrizz[99][581] = 9'b111111111;
assign micromatrizz[99][582] = 9'b111111111;
assign micromatrizz[99][583] = 9'b111111111;
assign micromatrizz[99][584] = 9'b111111111;
assign micromatrizz[99][585] = 9'b111111111;
assign micromatrizz[99][586] = 9'b111111111;
assign micromatrizz[99][587] = 9'b111111111;
assign micromatrizz[99][588] = 9'b111111111;
assign micromatrizz[99][589] = 9'b111111111;
assign micromatrizz[99][590] = 9'b111111111;
assign micromatrizz[99][591] = 9'b111111111;
assign micromatrizz[99][592] = 9'b111111111;
assign micromatrizz[99][593] = 9'b111111111;
assign micromatrizz[99][594] = 9'b111111111;
assign micromatrizz[99][595] = 9'b111111111;
assign micromatrizz[99][596] = 9'b111111111;
assign micromatrizz[99][597] = 9'b111111111;
assign micromatrizz[99][598] = 9'b111111111;
assign micromatrizz[99][599] = 9'b111111111;
assign micromatrizz[99][600] = 9'b111111111;
assign micromatrizz[99][601] = 9'b111111111;
assign micromatrizz[99][602] = 9'b111111111;
assign micromatrizz[99][603] = 9'b111111111;
assign micromatrizz[99][604] = 9'b111111111;
assign micromatrizz[99][605] = 9'b111111111;
assign micromatrizz[99][606] = 9'b111111111;
assign micromatrizz[99][607] = 9'b111111111;
assign micromatrizz[99][608] = 9'b111111111;
assign micromatrizz[99][609] = 9'b111111111;
assign micromatrizz[99][610] = 9'b111111111;
assign micromatrizz[99][611] = 9'b111111111;
assign micromatrizz[99][612] = 9'b111111111;
assign micromatrizz[99][613] = 9'b111111111;
assign micromatrizz[99][614] = 9'b111111111;
assign micromatrizz[99][615] = 9'b111111111;
assign micromatrizz[99][616] = 9'b111111111;
assign micromatrizz[99][617] = 9'b111111111;
assign micromatrizz[99][618] = 9'b111111111;
assign micromatrizz[99][619] = 9'b111111111;
assign micromatrizz[99][620] = 9'b111111111;
assign micromatrizz[99][621] = 9'b111111111;
assign micromatrizz[99][622] = 9'b111111111;
assign micromatrizz[99][623] = 9'b111111111;
assign micromatrizz[99][624] = 9'b111111111;
assign micromatrizz[99][625] = 9'b111111111;
assign micromatrizz[99][626] = 9'b111111111;
assign micromatrizz[99][627] = 9'b111111111;
assign micromatrizz[99][628] = 9'b111111111;
assign micromatrizz[99][629] = 9'b111111111;
assign micromatrizz[99][630] = 9'b111111111;
assign micromatrizz[99][631] = 9'b111111111;
assign micromatrizz[99][632] = 9'b111111111;
assign micromatrizz[99][633] = 9'b111111111;
assign micromatrizz[99][634] = 9'b111111111;
assign micromatrizz[99][635] = 9'b111111111;
assign micromatrizz[99][636] = 9'b111111111;
assign micromatrizz[99][637] = 9'b111111111;
assign micromatrizz[99][638] = 9'b111111111;
assign micromatrizz[99][639] = 9'b111111111;
//Total de Lineas = 64000
endmodule*/


