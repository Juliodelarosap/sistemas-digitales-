/*`timescale 1ns / 1ps
module boton_de_inicio (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (F[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= F[vcount- posy][hcount- posx][7:5];
				green <= F[vcount- posy][hcount- posx][4:2];
            blue 	<= F[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 50;
parameter RESOLUCION_Y = 100;
wire [8:0] F[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign F[35][4] = 9'b110011111;
assign F[35][5] = 9'b110011111;
assign F[35][6] = 9'b110011111;
assign F[35][7] = 9'b110011111;
assign F[35][8] = 9'b110011111;
assign F[35][9] = 9'b110011111;
assign F[35][10] = 9'b110011111;
assign F[35][11] = 9'b110011111;
assign F[35][12] = 9'b110011111;
assign F[35][13] = 9'b110011111;
assign F[35][14] = 9'b110011111;
assign F[35][15] = 9'b110011111;
assign F[35][16] = 9'b110011111;
assign F[35][17] = 9'b110011111;
assign F[35][18] = 9'b110011111;
assign F[35][19] = 9'b110011111;
assign F[35][20] = 9'b110011111;
assign F[35][21] = 9'b110011111;
assign F[35][22] = 9'b110011111;
assign F[35][23] = 9'b110011111;
assign F[35][24] = 9'b110011111;
assign F[35][25] = 9'b110011111;
assign F[35][26] = 9'b110011111;
assign F[35][27] = 9'b110011111;
assign F[35][28] = 9'b110011111;
assign F[35][29] = 9'b110011111;
assign F[35][30] = 9'b110011111;
assign F[35][31] = 9'b110011111;
assign F[35][32] = 9'b110011111;
assign F[35][33] = 9'b110011111;
assign F[35][34] = 9'b110011111;
assign F[35][35] = 9'b110011111;
assign F[35][36] = 9'b110011111;
assign F[35][37] = 9'b110011111;
assign F[35][38] = 9'b110011111;
assign F[35][39] = 9'b110011111;
assign F[35][40] = 9'b110011111;
assign F[35][41] = 9'b110011111;
assign F[35][42] = 9'b110011111;
assign F[35][43] = 9'b110011111;
assign F[35][44] = 9'b110011111;
assign F[35][45] = 9'b110011111;
assign F[36][2] = 9'b101001000;
assign F[36][3] = 9'b110010010;
assign F[36][4] = 9'b110111111;
assign F[36][5] = 9'b110111111;
assign F[36][6] = 9'b110111111;
assign F[36][7] = 9'b110111111;
assign F[36][8] = 9'b110111111;
assign F[36][9] = 9'b110111111;
assign F[36][10] = 9'b110111111;
assign F[36][11] = 9'b110111111;
assign F[36][12] = 9'b110111111;
assign F[36][13] = 9'b110111111;
assign F[36][14] = 9'b110111111;
assign F[36][15] = 9'b110111111;
assign F[36][16] = 9'b110111111;
assign F[36][17] = 9'b110111111;
assign F[36][18] = 9'b110111111;
assign F[36][19] = 9'b110111111;
assign F[36][20] = 9'b110111111;
assign F[36][21] = 9'b110111111;
assign F[36][22] = 9'b110111111;
assign F[36][23] = 9'b110111111;
assign F[36][24] = 9'b110111111;
assign F[36][25] = 9'b110111111;
assign F[36][26] = 9'b110111111;
assign F[36][27] = 9'b110111111;
assign F[36][28] = 9'b110111111;
assign F[36][29] = 9'b110111111;
assign F[36][30] = 9'b110111111;
assign F[36][31] = 9'b110111111;
assign F[36][32] = 9'b110111111;
assign F[36][33] = 9'b110111111;
assign F[36][34] = 9'b110111111;
assign F[36][35] = 9'b110111111;
assign F[36][36] = 9'b110111111;
assign F[36][37] = 9'b110111111;
assign F[36][38] = 9'b110111111;
assign F[36][39] = 9'b110111111;
assign F[36][40] = 9'b110111111;
assign F[36][41] = 9'b110111111;
assign F[36][42] = 9'b110111111;
assign F[36][43] = 9'b110111111;
assign F[36][44] = 9'b110111111;
assign F[36][45] = 9'b110111111;
assign F[36][46] = 9'b110010111;
assign F[36][47] = 9'b101001001;
assign F[37][2] = 9'b101001001;
assign F[37][3] = 9'b110011111;
assign F[37][4] = 9'b110011111;
assign F[37][5] = 9'b110011111;
assign F[37][6] = 9'b110011111;
assign F[37][7] = 9'b110011111;
assign F[37][8] = 9'b110011111;
assign F[37][9] = 9'b110011111;
assign F[37][10] = 9'b110011111;
assign F[37][11] = 9'b110011111;
assign F[37][12] = 9'b110011111;
assign F[37][13] = 9'b110011111;
assign F[37][14] = 9'b110011111;
assign F[37][15] = 9'b110011111;
assign F[37][16] = 9'b110011111;
assign F[37][17] = 9'b110011111;
assign F[37][18] = 9'b110011111;
assign F[37][19] = 9'b110011111;
assign F[37][20] = 9'b110011111;
assign F[37][21] = 9'b110011111;
assign F[37][22] = 9'b110011111;
assign F[37][23] = 9'b110011111;
assign F[37][24] = 9'b110011111;
assign F[37][25] = 9'b110011111;
assign F[37][26] = 9'b110011111;
assign F[37][27] = 9'b110011111;
assign F[37][28] = 9'b110011111;
assign F[37][29] = 9'b110011111;
assign F[37][30] = 9'b110011111;
assign F[37][31] = 9'b110011111;
assign F[37][32] = 9'b110011111;
assign F[37][33] = 9'b110011111;
assign F[37][34] = 9'b110011111;
assign F[37][35] = 9'b110011111;
assign F[37][36] = 9'b110011111;
assign F[37][37] = 9'b110011111;
assign F[37][38] = 9'b110011111;
assign F[37][39] = 9'b110011111;
assign F[37][40] = 9'b110011111;
assign F[37][41] = 9'b110011111;
assign F[37][42] = 9'b110011111;
assign F[37][43] = 9'b110011111;
assign F[37][44] = 9'b110011111;
assign F[37][45] = 9'b110011111;
assign F[37][46] = 9'b110111111;
assign F[37][47] = 9'b101101101;
assign F[38][2] = 9'b101001101;
assign F[38][3] = 9'b110011111;
assign F[38][4] = 9'b110011111;
assign F[38][5] = 9'b110011111;
assign F[38][6] = 9'b110011111;
assign F[38][7] = 9'b110011111;
assign F[38][8] = 9'b110011111;
assign F[38][9] = 9'b110011111;
assign F[38][10] = 9'b110011111;
assign F[38][11] = 9'b110011111;
assign F[38][12] = 9'b110011111;
assign F[38][13] = 9'b110011111;
assign F[38][14] = 9'b110011111;
assign F[38][15] = 9'b110011111;
assign F[38][16] = 9'b110011111;
assign F[38][17] = 9'b110011111;
assign F[38][18] = 9'b110011111;
assign F[38][19] = 9'b110011111;
assign F[38][20] = 9'b110011111;
assign F[38][21] = 9'b110011111;
assign F[38][22] = 9'b110011111;
assign F[38][23] = 9'b110011111;
assign F[38][24] = 9'b110011111;
assign F[38][25] = 9'b110011111;
assign F[38][26] = 9'b110011111;
assign F[38][27] = 9'b110011111;
assign F[38][28] = 9'b110011111;
assign F[38][29] = 9'b110011111;
assign F[38][30] = 9'b110011111;
assign F[38][31] = 9'b110011111;
assign F[38][32] = 9'b110011111;
assign F[38][33] = 9'b110011111;
assign F[38][34] = 9'b110011111;
assign F[38][35] = 9'b110011111;
assign F[38][36] = 9'b110011111;
assign F[38][37] = 9'b110011111;
assign F[38][38] = 9'b110011111;
assign F[38][39] = 9'b110011111;
assign F[38][40] = 9'b110011111;
assign F[38][41] = 9'b110011111;
assign F[38][42] = 9'b110011111;
assign F[38][43] = 9'b110011111;
assign F[38][44] = 9'b110011111;
assign F[38][45] = 9'b110011111;
assign F[38][46] = 9'b110011111;
assign F[38][47] = 9'b101101101;
assign F[38][48] = 9'b100100000;
assign F[39][2] = 9'b101001001;
assign F[39][3] = 9'b110011111;
assign F[39][4] = 9'b110011111;
assign F[39][5] = 9'b110011111;
assign F[39][6] = 9'b110011111;
assign F[39][7] = 9'b110011111;
assign F[39][8] = 9'b110011111;
assign F[39][9] = 9'b110011111;
assign F[39][10] = 9'b110011111;
assign F[39][11] = 9'b110011111;
assign F[39][12] = 9'b110010111;
assign F[39][13] = 9'b110010111;
assign F[39][14] = 9'b110010111;
assign F[39][15] = 9'b110011111;
assign F[39][16] = 9'b110010111;
assign F[39][17] = 9'b110010111;
assign F[39][18] = 9'b110010111;
assign F[39][19] = 9'b110010111;
assign F[39][20] = 9'b110010111;
assign F[39][21] = 9'b110011111;
assign F[39][22] = 9'b110011111;
assign F[39][23] = 9'b101110011;
assign F[39][24] = 9'b110011111;
assign F[39][25] = 9'b110011111;
assign F[39][26] = 9'b110011111;
assign F[39][27] = 9'b110011111;
assign F[39][28] = 9'b110010111;
assign F[39][29] = 9'b110010111;
assign F[39][30] = 9'b110010111;
assign F[39][31] = 9'b110011111;
assign F[39][32] = 9'b110011111;
assign F[39][33] = 9'b110010111;
assign F[39][34] = 9'b110010111;
assign F[39][35] = 9'b110010111;
assign F[39][36] = 9'b110010111;
assign F[39][37] = 9'b110010111;
assign F[39][38] = 9'b110011111;
assign F[39][39] = 9'b110011111;
assign F[39][40] = 9'b110011111;
assign F[39][41] = 9'b110011111;
assign F[39][42] = 9'b110011111;
assign F[39][43] = 9'b110011111;
assign F[39][44] = 9'b110011111;
assign F[39][45] = 9'b110011111;
assign F[39][46] = 9'b110011111;
assign F[39][47] = 9'b101101101;
assign F[40][2] = 9'b101001001;
assign F[40][3] = 9'b110011111;
assign F[40][4] = 9'b110011111;
assign F[40][5] = 9'b110011111;
assign F[40][6] = 9'b110011111;
assign F[40][7] = 9'b110011111;
assign F[40][8] = 9'b110011111;
assign F[40][9] = 9'b110011111;
assign F[40][10] = 9'b110011111;
assign F[40][11] = 9'b101110010;
assign F[40][12] = 9'b110010001;
assign F[40][13] = 9'b110010001;
assign F[40][14] = 9'b101101101;
assign F[40][15] = 9'b101001001;
assign F[40][16] = 9'b101101101;
assign F[40][17] = 9'b110010001;
assign F[40][18] = 9'b110010010;
assign F[40][19] = 9'b110010001;
assign F[40][20] = 9'b101101001;
assign F[40][21] = 9'b110010111;
assign F[40][22] = 9'b101110001;
assign F[40][23] = 9'b110010001;
assign F[40][24] = 9'b101101101;
assign F[40][25] = 9'b110011111;
assign F[40][26] = 9'b110011111;
assign F[40][27] = 9'b101101101;
assign F[40][28] = 9'b110010001;
assign F[40][29] = 9'b110010001;
assign F[40][30] = 9'b110010001;
assign F[40][31] = 9'b101110010;
assign F[40][32] = 9'b101110010;
assign F[40][33] = 9'b101101101;
assign F[40][34] = 9'b110010001;
assign F[40][35] = 9'b110010010;
assign F[40][36] = 9'b110010001;
assign F[40][37] = 9'b101101101;
assign F[40][38] = 9'b110010111;
assign F[40][39] = 9'b110011111;
assign F[40][40] = 9'b110011111;
assign F[40][41] = 9'b110011111;
assign F[40][42] = 9'b110011111;
assign F[40][43] = 9'b110011111;
assign F[40][44] = 9'b110011111;
assign F[40][45] = 9'b110011111;
assign F[40][46] = 9'b110011111;
assign F[40][47] = 9'b101101101;
assign F[41][2] = 9'b101001001;
assign F[41][3] = 9'b110011111;
assign F[41][4] = 9'b110011111;
assign F[41][5] = 9'b110011111;
assign F[41][6] = 9'b110011111;
assign F[41][7] = 9'b110011111;
assign F[41][8] = 9'b110011111;
assign F[41][9] = 9'b110011111;
assign F[41][10] = 9'b110010111;
assign F[41][11] = 9'b110010001;
assign F[41][12] = 9'b110010010;
assign F[41][13] = 9'b101110001;
assign F[41][14] = 9'b110010010;
assign F[41][15] = 9'b101110010;
assign F[41][16] = 9'b110010010;
assign F[41][17] = 9'b101110001;
assign F[41][18] = 9'b111111111;
assign F[41][19] = 9'b101101101;
assign F[41][20] = 9'b110010010;
assign F[41][21] = 9'b101110010;
assign F[41][22] = 9'b110010001;
assign F[41][23] = 9'b110001101;
assign F[41][24] = 9'b110010001;
assign F[41][25] = 9'b101110010;
assign F[41][26] = 9'b110011111;
assign F[41][27] = 9'b110010010;
assign F[41][28] = 9'b111110110;
assign F[41][29] = 9'b101110001;
assign F[41][30] = 9'b110010010;
assign F[41][31] = 9'b110110110;
assign F[41][32] = 9'b101101101;
assign F[41][33] = 9'b110010010;
assign F[41][34] = 9'b101110001;
assign F[41][35] = 9'b111111111;
assign F[41][36] = 9'b101101101;
assign F[41][37] = 9'b101110010;
assign F[41][38] = 9'b110011111;
assign F[41][39] = 9'b110011111;
assign F[41][40] = 9'b110011111;
assign F[41][41] = 9'b110011111;
assign F[41][42] = 9'b110011111;
assign F[41][43] = 9'b110011111;
assign F[41][44] = 9'b110011111;
assign F[41][45] = 9'b110011111;
assign F[41][46] = 9'b110011111;
assign F[41][47] = 9'b101101101;
assign F[42][2] = 9'b101001001;
assign F[42][3] = 9'b101110111;
assign F[42][4] = 9'b101110111;
assign F[42][5] = 9'b101110111;
assign F[42][6] = 9'b101110111;
assign F[42][7] = 9'b101110111;
assign F[42][8] = 9'b101110111;
assign F[42][9] = 9'b101110111;
assign F[42][10] = 9'b101110111;
assign F[42][11] = 9'b101101101;
assign F[42][12] = 9'b110110110;
assign F[42][13] = 9'b110010001;
assign F[42][14] = 9'b101110010;
assign F[42][15] = 9'b110011111;
assign F[42][16] = 9'b110011111;
assign F[42][17] = 9'b101110001;
assign F[42][18] = 9'b110110110;
assign F[42][19] = 9'b101110010;
assign F[42][20] = 9'b110011111;
assign F[42][21] = 9'b101110010;
assign F[42][22] = 9'b110010001;
assign F[42][23] = 9'b101001001;
assign F[42][24] = 9'b110010001;
assign F[42][25] = 9'b101110001;
assign F[42][26] = 9'b110011111;
assign F[42][27] = 9'b101110001;
assign F[42][28] = 9'b110110110;
assign F[42][29] = 9'b101101101;
assign F[42][30] = 9'b110010010;
assign F[42][31] = 9'b110010001;
assign F[42][32] = 9'b101110010;
assign F[42][33] = 9'b110111111;
assign F[42][34] = 9'b101110010;
assign F[42][35] = 9'b110110010;
assign F[42][36] = 9'b101110010;
assign F[42][37] = 9'b110111111;
assign F[42][38] = 9'b110011111;
assign F[42][39] = 9'b110011111;
assign F[42][40] = 9'b110011111;
assign F[42][41] = 9'b110011111;
assign F[42][42] = 9'b110011111;
assign F[42][43] = 9'b110011111;
assign F[42][44] = 9'b110011111;
assign F[42][45] = 9'b110011111;
assign F[42][46] = 9'b110011111;
assign F[42][47] = 9'b101101101;
assign F[43][2] = 9'b101001001;
assign F[43][3] = 9'b101110111;
assign F[43][4] = 9'b101110111;
assign F[43][5] = 9'b101110111;
assign F[43][6] = 9'b101110111;
assign F[43][7] = 9'b101110111;
assign F[43][8] = 9'b101110111;
assign F[43][9] = 9'b101110111;
assign F[43][10] = 9'b101110111;
assign F[43][11] = 9'b101010011;
assign F[43][12] = 9'b101001101;
assign F[43][13] = 9'b110010010;
assign F[43][14] = 9'b110010001;
assign F[43][15] = 9'b101001101;
assign F[43][16] = 9'b101110111;
assign F[43][17] = 9'b101001101;
assign F[43][18] = 9'b111110110;
assign F[43][19] = 9'b101001101;
assign F[43][20] = 9'b101010011;
assign F[43][21] = 9'b101110001;
assign F[43][22] = 9'b111111110;
assign F[43][23] = 9'b101001101;
assign F[43][24] = 9'b110110110;
assign F[43][25] = 9'b110010010;
assign F[43][26] = 9'b101010011;
assign F[43][27] = 9'b101110001;
assign F[43][28] = 9'b111111111;
assign F[43][29] = 9'b110010001;
assign F[43][30] = 9'b111110110;
assign F[43][31] = 9'b101001101;
assign F[43][32] = 9'b101111111;
assign F[43][33] = 9'b101111111;
assign F[43][34] = 9'b101110010;
assign F[43][35] = 9'b110110010;
assign F[43][36] = 9'b101110010;
assign F[43][37] = 9'b110011111;
assign F[43][38] = 9'b110011111;
assign F[43][39] = 9'b110011111;
assign F[43][40] = 9'b110011111;
assign F[43][41] = 9'b110011111;
assign F[43][42] = 9'b110011111;
assign F[43][43] = 9'b110011111;
assign F[43][44] = 9'b110011111;
assign F[43][45] = 9'b110011111;
assign F[43][46] = 9'b110011111;
assign F[43][47] = 9'b101101101;
assign F[44][2] = 9'b101001001;
assign F[44][3] = 9'b101110111;
assign F[44][4] = 9'b101110111;
assign F[44][5] = 9'b101110111;
assign F[44][6] = 9'b101110111;
assign F[44][7] = 9'b101110111;
assign F[44][8] = 9'b101110111;
assign F[44][9] = 9'b101110111;
assign F[44][10] = 9'b101110011;
assign F[44][11] = 9'b101001101;
assign F[44][12] = 9'b101010011;
assign F[44][13] = 9'b101001101;
assign F[44][14] = 9'b111111110;
assign F[44][15] = 9'b101101101;
assign F[44][16] = 9'b101110111;
assign F[44][17] = 9'b101101101;
assign F[44][18] = 9'b111111110;
assign F[44][19] = 9'b101010010;
assign F[44][20] = 9'b101010010;
assign F[44][21] = 9'b110110110;
assign F[44][22] = 9'b110010010;
assign F[44][23] = 9'b101110001;
assign F[44][24] = 9'b110010001;
assign F[44][25] = 9'b111111110;
assign F[44][26] = 9'b101001101;
assign F[44][27] = 9'b101110010;
assign F[44][28] = 9'b110110110;
assign F[44][29] = 9'b100101001;
assign F[44][30] = 9'b110010001;
assign F[44][31] = 9'b110010001;
assign F[44][32] = 9'b101010011;
assign F[44][33] = 9'b101110111;
assign F[44][34] = 9'b101001101;
assign F[44][35] = 9'b111110110;
assign F[44][36] = 9'b101001110;
assign F[44][37] = 9'b101110111;
assign F[44][38] = 9'b101110111;
assign F[44][39] = 9'b110011111;
assign F[44][40] = 9'b110011111;
assign F[44][41] = 9'b110011111;
assign F[44][42] = 9'b110011111;
assign F[44][43] = 9'b110011111;
assign F[44][44] = 9'b110011111;
assign F[44][45] = 9'b110011111;
assign F[44][46] = 9'b110011111;
assign F[44][47] = 9'b101101101;
assign F[45][2] = 9'b101001001;
assign F[45][3] = 9'b101110111;
assign F[45][4] = 9'b101110111;
assign F[45][5] = 9'b101110111;
assign F[45][6] = 9'b101110111;
assign F[45][7] = 9'b101110111;
assign F[45][8] = 9'b101110111;
assign F[45][9] = 9'b101110111;
assign F[45][10] = 9'b101010011;
assign F[45][11] = 9'b101101101;
assign F[45][12] = 9'b110010001;
assign F[45][13] = 9'b110010001;
assign F[45][14] = 9'b110010001;
assign F[45][15] = 9'b101010010;
assign F[45][16] = 9'b101110111;
assign F[45][17] = 9'b101001101;
assign F[45][18] = 9'b110001101;
assign F[45][19] = 9'b101001110;
assign F[45][20] = 9'b101001101;
assign F[45][21] = 9'b110010001;
assign F[45][22] = 9'b101001101;
assign F[45][23] = 9'b101110111;
assign F[45][24] = 9'b101001110;
assign F[45][25] = 9'b110010001;
assign F[45][26] = 9'b101001101;
assign F[45][27] = 9'b101001101;
assign F[45][28] = 9'b110001101;
assign F[45][29] = 9'b101010011;
assign F[45][30] = 9'b101001110;
assign F[45][31] = 9'b110010001;
assign F[45][32] = 9'b101001001;
assign F[45][33] = 9'b101110111;
assign F[45][34] = 9'b101001101;
assign F[45][35] = 9'b110001101;
assign F[45][36] = 9'b101001110;
assign F[45][37] = 9'b101110111;
assign F[45][38] = 9'b101110111;
assign F[45][39] = 9'b101110111;
assign F[45][40] = 9'b101110111;
assign F[45][41] = 9'b101110111;
assign F[45][42] = 9'b110011111;
assign F[45][43] = 9'b110011111;
assign F[45][44] = 9'b110011111;
assign F[45][45] = 9'b110011111;
assign F[45][46] = 9'b110011111;
assign F[45][47] = 9'b101101101;
assign F[46][2] = 9'b101001001;
assign F[46][3] = 9'b101110111;
assign F[46][4] = 9'b101110111;
assign F[46][5] = 9'b101110111;
assign F[46][6] = 9'b101110111;
assign F[46][7] = 9'b101110111;
assign F[46][8] = 9'b101110111;
assign F[46][9] = 9'b101110111;
assign F[46][10] = 9'b101110111;
assign F[46][11] = 9'b101010011;
assign F[46][12] = 9'b101010010;
assign F[46][13] = 9'b101010010;
assign F[46][14] = 9'b101010011;
assign F[46][15] = 9'b101110111;
assign F[46][16] = 9'b101110111;
assign F[46][17] = 9'b101110011;
assign F[46][18] = 9'b101010010;
assign F[46][19] = 9'b101110011;
assign F[46][20] = 9'b101110011;
assign F[46][21] = 9'b101010010;
assign F[46][22] = 9'b101110011;
assign F[46][23] = 9'b101110111;
assign F[46][24] = 9'b101110111;
assign F[46][25] = 9'b101010010;
assign F[46][26] = 9'b101010010;
assign F[46][27] = 9'b101010011;
assign F[46][28] = 9'b101010010;
assign F[46][29] = 9'b101110111;
assign F[46][30] = 9'b101110111;
assign F[46][31] = 9'b101010010;
assign F[46][32] = 9'b101010010;
assign F[46][33] = 9'b101110111;
assign F[46][34] = 9'b101110011;
assign F[46][35] = 9'b101010010;
assign F[46][36] = 9'b101110011;
assign F[46][37] = 9'b101110111;
assign F[46][38] = 9'b101110111;
assign F[46][39] = 9'b101110111;
assign F[46][40] = 9'b101110111;
assign F[46][41] = 9'b101110111;
assign F[46][42] = 9'b101110111;
assign F[46][43] = 9'b101110111;
assign F[46][44] = 9'b110011111;
assign F[46][45] = 9'b110011111;
assign F[46][46] = 9'b110111111;
assign F[46][47] = 9'b101101101;
assign F[47][2] = 9'b101001001;
assign F[47][3] = 9'b101110111;
assign F[47][4] = 9'b101110111;
assign F[47][5] = 9'b101110111;
assign F[47][6] = 9'b101110111;
assign F[47][7] = 9'b101110111;
assign F[47][8] = 9'b101110111;
assign F[47][9] = 9'b101110111;
assign F[47][10] = 9'b101110111;
assign F[47][11] = 9'b101110111;
assign F[47][12] = 9'b101110111;
assign F[47][13] = 9'b101110111;
assign F[47][14] = 9'b101110111;
assign F[47][15] = 9'b101110111;
assign F[47][16] = 9'b101110111;
assign F[47][17] = 9'b101110111;
assign F[47][18] = 9'b101110111;
assign F[47][19] = 9'b101110111;
assign F[47][20] = 9'b101110111;
assign F[47][21] = 9'b101110111;
assign F[47][22] = 9'b101110111;
assign F[47][23] = 9'b101110111;
assign F[47][24] = 9'b101110111;
assign F[47][25] = 9'b101110111;
assign F[47][26] = 9'b101110111;
assign F[47][27] = 9'b101110111;
assign F[47][28] = 9'b101110111;
assign F[47][29] = 9'b101110111;
assign F[47][30] = 9'b101110111;
assign F[47][31] = 9'b101110111;
assign F[47][32] = 9'b101110111;
assign F[47][33] = 9'b101110111;
assign F[47][34] = 9'b101110111;
assign F[47][35] = 9'b101110111;
assign F[47][36] = 9'b101110111;
assign F[47][37] = 9'b101110111;
assign F[47][38] = 9'b101110111;
assign F[47][39] = 9'b101110111;
assign F[47][40] = 9'b101110111;
assign F[47][41] = 9'b101110111;
assign F[47][42] = 9'b101110111;
assign F[47][43] = 9'b101110111;
assign F[47][44] = 9'b101110111;
assign F[47][45] = 9'b101110111;
assign F[47][46] = 9'b110011111;
assign F[47][47] = 9'b101101101;
assign F[48][2] = 9'b101001001;
assign F[48][3] = 9'b101110111;
assign F[48][4] = 9'b101110111;
assign F[48][5] = 9'b101110111;
assign F[48][6] = 9'b101110111;
assign F[48][7] = 9'b101110111;
assign F[48][8] = 9'b101110111;
assign F[48][9] = 9'b101110111;
assign F[48][10] = 9'b101110111;
assign F[48][11] = 9'b101110111;
assign F[48][12] = 9'b101110111;
assign F[48][13] = 9'b101110111;
assign F[48][14] = 9'b101110111;
assign F[48][15] = 9'b101110111;
assign F[48][16] = 9'b101110111;
assign F[48][17] = 9'b101110111;
assign F[48][18] = 9'b101110111;
assign F[48][19] = 9'b101110111;
assign F[48][20] = 9'b101110111;
assign F[48][21] = 9'b101110111;
assign F[48][22] = 9'b101110111;
assign F[48][23] = 9'b101110111;
assign F[48][24] = 9'b101110111;
assign F[48][25] = 9'b101110111;
assign F[48][26] = 9'b101110111;
assign F[48][27] = 9'b101110111;
assign F[48][28] = 9'b101110111;
assign F[48][29] = 9'b101110111;
assign F[48][30] = 9'b101110111;
assign F[48][31] = 9'b101110111;
assign F[48][32] = 9'b101110111;
assign F[48][33] = 9'b101110111;
assign F[48][34] = 9'b101110111;
assign F[48][35] = 9'b101110111;
assign F[48][36] = 9'b101110111;
assign F[48][37] = 9'b101110111;
assign F[48][38] = 9'b101110111;
assign F[48][39] = 9'b101110111;
assign F[48][40] = 9'b101110111;
assign F[48][41] = 9'b101110111;
assign F[48][42] = 9'b101110111;
assign F[48][43] = 9'b101110111;
assign F[48][44] = 9'b101110111;
assign F[48][45] = 9'b101110111;
assign F[48][46] = 9'b101110111;
assign F[48][47] = 9'b101001101;
assign F[49][2] = 9'b101001001;
assign F[49][3] = 9'b101110111;
assign F[49][4] = 9'b101110111;
assign F[49][5] = 9'b101110111;
assign F[49][6] = 9'b101110111;
assign F[49][7] = 9'b101110111;
assign F[49][8] = 9'b101110111;
assign F[49][9] = 9'b101110111;
assign F[49][10] = 9'b101110111;
assign F[49][11] = 9'b101110111;
assign F[49][12] = 9'b101110111;
assign F[49][13] = 9'b101110111;
assign F[49][14] = 9'b101110111;
assign F[49][15] = 9'b101110111;
assign F[49][16] = 9'b101110111;
assign F[49][17] = 9'b101110111;
assign F[49][18] = 9'b101110111;
assign F[49][19] = 9'b101110111;
assign F[49][20] = 9'b101110111;
assign F[49][21] = 9'b101110111;
assign F[49][22] = 9'b101110111;
assign F[49][23] = 9'b101110111;
assign F[49][24] = 9'b101110111;
assign F[49][25] = 9'b101110111;
assign F[49][26] = 9'b101110111;
assign F[49][27] = 9'b101110111;
assign F[49][28] = 9'b101110111;
assign F[49][29] = 9'b101110111;
assign F[49][30] = 9'b101110111;
assign F[49][31] = 9'b101110111;
assign F[49][32] = 9'b101110111;
assign F[49][33] = 9'b101110111;
assign F[49][34] = 9'b101110111;
assign F[49][35] = 9'b101110111;
assign F[49][36] = 9'b101110111;
assign F[49][37] = 9'b101110111;
assign F[49][38] = 9'b101110111;
assign F[49][39] = 9'b101110111;
assign F[49][40] = 9'b101110111;
assign F[49][41] = 9'b101110111;
assign F[49][42] = 9'b101110111;
assign F[49][43] = 9'b101110111;
assign F[49][44] = 9'b101110111;
assign F[49][45] = 9'b101110111;
assign F[49][46] = 9'b101110111;
assign F[49][47] = 9'b101001101;
assign F[50][2] = 9'b101001001;
assign F[50][3] = 9'b101010010;
assign F[50][4] = 9'b101110011;
assign F[50][5] = 9'b101110111;
assign F[50][6] = 9'b101110111;
assign F[50][7] = 9'b101110111;
assign F[50][8] = 9'b101110111;
assign F[50][9] = 9'b101110111;
assign F[50][10] = 9'b101110111;
assign F[50][11] = 9'b101110111;
assign F[50][12] = 9'b101110111;
assign F[50][13] = 9'b101110111;
assign F[50][14] = 9'b101110111;
assign F[50][15] = 9'b101110111;
assign F[50][16] = 9'b101110111;
assign F[50][17] = 9'b101110111;
assign F[50][18] = 9'b101110111;
assign F[50][19] = 9'b101110111;
assign F[50][20] = 9'b101110111;
assign F[50][21] = 9'b101110111;
assign F[50][22] = 9'b101110111;
assign F[50][23] = 9'b101110111;
assign F[50][24] = 9'b101110111;
assign F[50][25] = 9'b101110111;
assign F[50][26] = 9'b101110111;
assign F[50][27] = 9'b101110111;
assign F[50][28] = 9'b101110111;
assign F[50][29] = 9'b101110111;
assign F[50][30] = 9'b101110111;
assign F[50][31] = 9'b101110111;
assign F[50][32] = 9'b101110111;
assign F[50][33] = 9'b101110111;
assign F[50][34] = 9'b101110111;
assign F[50][35] = 9'b101110111;
assign F[50][36] = 9'b101110111;
assign F[50][37] = 9'b101110111;
assign F[50][38] = 9'b101110111;
assign F[50][39] = 9'b101110111;
assign F[50][40] = 9'b101110111;
assign F[50][41] = 9'b101110111;
assign F[50][42] = 9'b101110111;
assign F[50][43] = 9'b101110111;
assign F[50][44] = 9'b101110111;
assign F[50][45] = 9'b101110011;
assign F[50][46] = 9'b101010011;
assign F[50][47] = 9'b101001001;
assign F[50][48] = 9'b101000100;
assign F[51][2] = 9'b101000100;
assign F[51][3] = 9'b101001001;
assign F[51][4] = 9'b101001110;
assign F[51][5] = 9'b101001110;
assign F[51][6] = 9'b101001110;
assign F[51][7] = 9'b101001110;
assign F[51][8] = 9'b101001110;
assign F[51][9] = 9'b101001110;
assign F[51][10] = 9'b101001110;
assign F[51][11] = 9'b101001110;
assign F[51][12] = 9'b101001110;
assign F[51][13] = 9'b101001110;
assign F[51][14] = 9'b101001110;
assign F[51][15] = 9'b101001110;
assign F[51][16] = 9'b101001110;
assign F[51][17] = 9'b101001110;
assign F[51][18] = 9'b101001110;
assign F[51][19] = 9'b101001110;
assign F[51][20] = 9'b101001110;
assign F[51][21] = 9'b101001110;
assign F[51][22] = 9'b101001110;
assign F[51][23] = 9'b101001110;
assign F[51][24] = 9'b101001110;
assign F[51][25] = 9'b101001110;
assign F[51][26] = 9'b101001110;
assign F[51][27] = 9'b101001110;
assign F[51][28] = 9'b101001110;
assign F[51][29] = 9'b101001110;
assign F[51][30] = 9'b101001110;
assign F[51][31] = 9'b101001110;
assign F[51][32] = 9'b101001110;
assign F[51][33] = 9'b101001110;
assign F[51][34] = 9'b101001110;
assign F[51][35] = 9'b101001110;
assign F[51][36] = 9'b101001110;
assign F[51][37] = 9'b101001110;
assign F[51][38] = 9'b101001110;
assign F[51][39] = 9'b101001110;
assign F[51][40] = 9'b101001110;
assign F[51][41] = 9'b101001110;
assign F[51][42] = 9'b101001110;
assign F[51][43] = 9'b101001110;
assign F[51][44] = 9'b101001110;
assign F[51][45] = 9'b101001110;
assign F[51][46] = 9'b101001101;
assign F[51][47] = 9'b101001000;
assign F[52][2] = 9'b101001000;
assign F[52][3] = 9'b101001000;
assign F[52][4] = 9'b101001001;
assign F[52][5] = 9'b101001001;
assign F[52][6] = 9'b101001001;
assign F[52][7] = 9'b101001001;
assign F[52][8] = 9'b101001001;
assign F[52][9] = 9'b101001001;
assign F[52][10] = 9'b101001001;
assign F[52][11] = 9'b101001001;
assign F[52][12] = 9'b101001001;
assign F[52][13] = 9'b101001001;
assign F[52][14] = 9'b101001001;
assign F[52][15] = 9'b101001001;
assign F[52][16] = 9'b101001001;
assign F[52][17] = 9'b101001001;
assign F[52][18] = 9'b101001001;
assign F[52][19] = 9'b101001001;
assign F[52][20] = 9'b101001001;
assign F[52][21] = 9'b101001001;
assign F[52][22] = 9'b101001001;
assign F[52][23] = 9'b101001001;
assign F[52][24] = 9'b101001001;
assign F[52][25] = 9'b101001001;
assign F[52][26] = 9'b101001001;
assign F[52][27] = 9'b101001001;
assign F[52][28] = 9'b101001001;
assign F[52][29] = 9'b101001001;
assign F[52][30] = 9'b101001001;
assign F[52][31] = 9'b101001001;
assign F[52][32] = 9'b101001001;
assign F[52][33] = 9'b101001001;
assign F[52][34] = 9'b101001001;
assign F[52][35] = 9'b101001001;
assign F[52][36] = 9'b101001001;
assign F[52][37] = 9'b101001001;
assign F[52][38] = 9'b101001001;
assign F[52][39] = 9'b101001001;
assign F[52][40] = 9'b101001001;
assign F[52][41] = 9'b101001001;
assign F[52][42] = 9'b101001001;
assign F[52][43] = 9'b101001001;
assign F[52][44] = 9'b101001001;
assign F[52][45] = 9'b101001001;
assign F[52][46] = 9'b101001000;
assign F[52][47] = 9'b101001000;
assign F[53][3] = 9'b101001000;
assign F[53][4] = 9'b101000100;
assign F[53][5] = 9'b101000100;
assign F[53][6] = 9'b101000100;
assign F[53][7] = 9'b101000100;
assign F[53][8] = 9'b101000100;
assign F[53][9] = 9'b101000100;
assign F[53][10] = 9'b101000100;
assign F[53][11] = 9'b101000100;
assign F[53][12] = 9'b101000100;
assign F[53][13] = 9'b101000100;
assign F[53][14] = 9'b101000100;
assign F[53][15] = 9'b101000100;
assign F[53][16] = 9'b101000100;
assign F[53][17] = 9'b101000100;
assign F[53][18] = 9'b101000100;
assign F[53][19] = 9'b101000100;
assign F[53][20] = 9'b101000100;
assign F[53][21] = 9'b101000100;
assign F[53][22] = 9'b101000100;
assign F[53][23] = 9'b101000100;
assign F[53][24] = 9'b101000100;
assign F[53][25] = 9'b101000100;
assign F[53][26] = 9'b101000100;
assign F[53][27] = 9'b101000100;
assign F[53][28] = 9'b101000100;
assign F[53][29] = 9'b101000100;
assign F[53][30] = 9'b101000100;
assign F[53][31] = 9'b101000100;
assign F[53][32] = 9'b101000100;
assign F[53][33] = 9'b101000100;
assign F[53][34] = 9'b101000100;
assign F[53][35] = 9'b101000100;
assign F[53][36] = 9'b101000100;
assign F[53][37] = 9'b101000100;
assign F[53][38] = 9'b101000100;
assign F[53][39] = 9'b101000100;
assign F[53][40] = 9'b101000100;
assign F[53][41] = 9'b101000100;
assign F[53][42] = 9'b101000100;
assign F[53][43] = 9'b101000100;
assign F[53][44] = 9'b101000100;
assign F[53][45] = 9'b101000100;
assign F[53][46] = 9'b101001000;
//Total de Lineas = 870
endmodule*/

