`timescale 1ns / 1ps
/*module el_nano (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (F[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= F[vcount- posy][hcount- posx][7:5];
				green <= F[vcount- posy][hcount- posx][4:2];
            blue 	<= F[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 100;
parameter RESOLUCION_Y = 100;
wire [8:0] F[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign F[13][38] = 9'b101101001;
assign F[13][39] = 9'b101101000;
assign F[13][40] = 9'b100100000;
assign F[13][41] = 9'b101101000;
assign F[13][42] = 9'b101101000;
assign F[13][43] = 9'b101001000;
assign F[13][44] = 9'b101000100;
assign F[13][45] = 9'b101000100;
assign F[13][46] = 9'b100100000;
assign F[13][47] = 9'b100000000;
assign F[13][48] = 9'b100000000;
assign F[13][49] = 9'b100000000;
assign F[13][50] = 9'b100000000;
assign F[13][51] = 9'b100000000;
assign F[13][52] = 9'b100000000;
assign F[13][53] = 9'b100000000;
assign F[13][54] = 9'b100100000;
assign F[13][55] = 9'b100100100;
assign F[13][56] = 9'b100100100;
assign F[13][57] = 9'b100000000;
assign F[13][58] = 9'b100000000;
assign F[13][59] = 9'b100100000;
assign F[13][60] = 9'b101000100;
assign F[13][61] = 9'b100000000;
assign F[13][62] = 9'b100000000;
assign F[14][37] = 9'b101101101;
assign F[14][38] = 9'b101001000;
assign F[14][39] = 9'b101101000;
assign F[14][40] = 9'b101000100;
assign F[14][41] = 9'b101101000;
assign F[14][42] = 9'b101101000;
assign F[14][43] = 9'b101000100;
assign F[14][44] = 9'b101000100;
assign F[14][45] = 9'b101000100;
assign F[14][46] = 9'b100100100;
assign F[14][47] = 9'b100100100;
assign F[14][48] = 9'b100100100;
assign F[14][49] = 9'b100100100;
assign F[14][50] = 9'b100100000;
assign F[14][51] = 9'b100100000;
assign F[14][52] = 9'b100100000;
assign F[14][53] = 9'b100100000;
assign F[14][54] = 9'b100100000;
assign F[14][55] = 9'b101000100;
assign F[14][56] = 9'b101000100;
assign F[14][57] = 9'b100100100;
assign F[14][58] = 9'b100100000;
assign F[14][59] = 9'b100100100;
assign F[14][60] = 9'b101000100;
assign F[14][61] = 9'b100100000;
assign F[14][62] = 9'b100000000;
assign F[14][63] = 9'b100000000;
assign F[15][36] = 9'b101101000;
assign F[15][37] = 9'b101101000;
assign F[15][38] = 9'b101000100;
assign F[15][39] = 9'b101000100;
assign F[15][40] = 9'b101101000;
assign F[15][41] = 9'b101101000;
assign F[15][42] = 9'b101001000;
assign F[15][43] = 9'b101000100;
assign F[15][44] = 9'b100100100;
assign F[15][45] = 9'b100100100;
assign F[15][46] = 9'b100100100;
assign F[15][47] = 9'b100100100;
assign F[15][48] = 9'b100100100;
assign F[15][49] = 9'b100100100;
assign F[15][50] = 9'b100100000;
assign F[15][51] = 9'b100100000;
assign F[15][52] = 9'b100100000;
assign F[15][53] = 9'b100100000;
assign F[15][54] = 9'b100100000;
assign F[15][55] = 9'b100100100;
assign F[15][56] = 9'b100100100;
assign F[15][57] = 9'b100100100;
assign F[15][58] = 9'b101000100;
assign F[15][59] = 9'b101000100;
assign F[15][60] = 9'b100100100;
assign F[15][61] = 9'b101000100;
assign F[15][62] = 9'b100100100;
assign F[15][63] = 9'b100000000;
assign F[15][64] = 9'b100000000;
assign F[16][35] = 9'b101101000;
assign F[16][36] = 9'b101101000;
assign F[16][37] = 9'b101000100;
assign F[16][38] = 9'b101101000;
assign F[16][39] = 9'b101101000;
assign F[16][40] = 9'b101101000;
assign F[16][41] = 9'b101000100;
assign F[16][42] = 9'b100100100;
assign F[16][43] = 9'b101000100;
assign F[16][44] = 9'b100100000;
assign F[16][45] = 9'b100000000;
assign F[16][46] = 9'b100100000;
assign F[16][47] = 9'b100100000;
assign F[16][48] = 9'b100100000;
assign F[16][49] = 9'b100100000;
assign F[16][50] = 9'b100100000;
assign F[16][51] = 9'b100100000;
assign F[16][52] = 9'b100100000;
assign F[16][53] = 9'b100100000;
assign F[16][54] = 9'b100100000;
assign F[16][55] = 9'b100100000;
assign F[16][56] = 9'b100000000;
assign F[16][57] = 9'b100100000;
assign F[16][58] = 9'b101000100;
assign F[16][59] = 9'b101000100;
assign F[16][60] = 9'b101000100;
assign F[16][61] = 9'b101000100;
assign F[16][62] = 9'b101000100;
assign F[16][63] = 9'b100100100;
assign F[16][64] = 9'b100000000;
assign F[16][65] = 9'b100000000;
assign F[17][33] = 9'b101101000;
assign F[17][34] = 9'b101101000;
assign F[17][35] = 9'b101101000;
assign F[17][36] = 9'b101101000;
assign F[17][37] = 9'b101101000;
assign F[17][38] = 9'b101101000;
assign F[17][39] = 9'b101101000;
assign F[17][40] = 9'b101000100;
assign F[17][41] = 9'b101000100;
assign F[17][42] = 9'b100100100;
assign F[17][43] = 9'b100100100;
assign F[17][44] = 9'b100100000;
assign F[17][45] = 9'b100100000;
assign F[17][46] = 9'b100100000;
assign F[17][47] = 9'b100100000;
assign F[17][48] = 9'b100100000;
assign F[17][49] = 9'b100100000;
assign F[17][50] = 9'b100100000;
assign F[17][51] = 9'b100000000;
assign F[17][52] = 9'b100000000;
assign F[17][53] = 9'b100100000;
assign F[17][54] = 9'b100100000;
assign F[17][55] = 9'b100000000;
assign F[17][56] = 9'b100000000;
assign F[17][57] = 9'b100100000;
assign F[17][58] = 9'b100100100;
assign F[17][59] = 9'b101000100;
assign F[17][60] = 9'b101000100;
assign F[17][61] = 9'b100100000;
assign F[17][62] = 9'b100000000;
assign F[17][63] = 9'b100000000;
assign F[17][64] = 9'b100000000;
assign F[17][65] = 9'b100000000;
assign F[18][32] = 9'b101101000;
assign F[18][33] = 9'b101101000;
assign F[18][34] = 9'b101101000;
assign F[18][35] = 9'b101101000;
assign F[18][36] = 9'b101101000;
assign F[18][37] = 9'b101101000;
assign F[18][38] = 9'b101000100;
assign F[18][39] = 9'b100100100;
assign F[18][40] = 9'b101000100;
assign F[18][41] = 9'b100100100;
assign F[18][42] = 9'b100100100;
assign F[18][43] = 9'b100100100;
assign F[18][44] = 9'b100100100;
assign F[18][45] = 9'b101000100;
assign F[18][46] = 9'b101101000;
assign F[18][47] = 9'b101101000;
assign F[18][48] = 9'b101101000;
assign F[18][49] = 9'b101101000;
assign F[18][50] = 9'b101000100;
assign F[18][51] = 9'b100100000;
assign F[18][52] = 9'b100100100;
assign F[18][53] = 9'b100100100;
assign F[18][54] = 9'b100100100;
assign F[18][55] = 9'b100100100;
assign F[18][56] = 9'b100100100;
assign F[18][57] = 9'b100100100;
assign F[18][58] = 9'b101000100;
assign F[18][59] = 9'b101000100;
assign F[18][60] = 9'b101000100;
assign F[18][61] = 9'b100100100;
assign F[18][62] = 9'b100100000;
assign F[18][63] = 9'b100000000;
assign F[18][64] = 9'b100100100;
assign F[18][65] = 9'b100100100;
assign F[18][66] = 9'b100000000;
assign F[18][67] = 9'b100000000;
assign F[18][68] = 9'b100000000;
assign F[19][32] = 9'b101101000;
assign F[19][33] = 9'b101101000;
assign F[19][34] = 9'b101101000;
assign F[19][35] = 9'b101101000;
assign F[19][36] = 9'b101101000;
assign F[19][37] = 9'b101000100;
assign F[19][38] = 9'b100100100;
assign F[19][39] = 9'b100100100;
assign F[19][40] = 9'b100100100;
assign F[19][41] = 9'b101000100;
assign F[19][42] = 9'b101101000;
assign F[19][43] = 9'b101101000;
assign F[19][44] = 9'b101101000;
assign F[19][45] = 9'b101101000;
assign F[19][46] = 9'b101101000;
assign F[19][47] = 9'b101101000;
assign F[19][48] = 9'b101101000;
assign F[19][49] = 9'b101101000;
assign F[19][50] = 9'b101101000;
assign F[19][51] = 9'b101101000;
assign F[19][52] = 9'b101101000;
assign F[19][53] = 9'b101101000;
assign F[19][54] = 9'b101101000;
assign F[19][55] = 9'b101101000;
assign F[19][56] = 9'b101101000;
assign F[19][57] = 9'b101101000;
assign F[19][58] = 9'b101101000;
assign F[19][59] = 9'b101101000;
assign F[19][60] = 9'b101101000;
assign F[19][61] = 9'b101101000;
assign F[19][62] = 9'b101000100;
assign F[19][63] = 9'b100000000;
assign F[19][64] = 9'b100100000;
assign F[19][65] = 9'b100100000;
assign F[19][66] = 9'b100100100;
assign F[19][67] = 9'b100000000;
assign F[19][68] = 9'b100000000;
assign F[20][31] = 9'b101101001;
assign F[20][32] = 9'b101101000;
assign F[20][33] = 9'b101101000;
assign F[20][34] = 9'b101101000;
assign F[20][35] = 9'b101001000;
assign F[20][36] = 9'b101000100;
assign F[20][37] = 9'b100100100;
assign F[20][38] = 9'b100100100;
assign F[20][39] = 9'b100100100;
assign F[20][40] = 9'b100100100;
assign F[20][41] = 9'b101101000;
assign F[20][42] = 9'b110001000;
assign F[20][43] = 9'b110001101;
assign F[20][44] = 9'b110001101;
assign F[20][45] = 9'b110001101;
assign F[20][46] = 9'b101101000;
assign F[20][47] = 9'b101101000;
assign F[20][48] = 9'b101101000;
assign F[20][49] = 9'b110001101;
assign F[20][50] = 9'b110001101;
assign F[20][51] = 9'b110001101;
assign F[20][52] = 9'b110001101;
assign F[20][53] = 9'b110001101;
assign F[20][54] = 9'b110001101;
assign F[20][55] = 9'b110001101;
assign F[20][56] = 9'b110001101;
assign F[20][57] = 9'b110001101;
assign F[20][58] = 9'b110001101;
assign F[20][59] = 9'b110001101;
assign F[20][60] = 9'b110001101;
assign F[20][61] = 9'b110001101;
assign F[20][62] = 9'b101101000;
assign F[20][63] = 9'b101000100;
assign F[20][64] = 9'b100100000;
assign F[20][65] = 9'b100100000;
assign F[20][66] = 9'b100100100;
assign F[20][67] = 9'b100100000;
assign F[20][68] = 9'b100000000;
assign F[20][69] = 9'b100000000;
assign F[21][30] = 9'b101001000;
assign F[21][31] = 9'b101101000;
assign F[21][32] = 9'b101101000;
assign F[21][33] = 9'b101001000;
assign F[21][34] = 9'b101101000;
assign F[21][35] = 9'b101000100;
assign F[21][36] = 9'b100100100;
assign F[21][37] = 9'b100100100;
assign F[21][38] = 9'b101000100;
assign F[21][39] = 9'b101000100;
assign F[21][40] = 9'b101000100;
assign F[21][41] = 9'b101101000;
assign F[21][42] = 9'b110001101;
assign F[21][43] = 9'b110101101;
assign F[21][44] = 9'b110101101;
assign F[21][45] = 9'b110101101;
assign F[21][46] = 9'b110001000;
assign F[21][47] = 9'b110001001;
assign F[21][48] = 9'b110001101;
assign F[21][49] = 9'b110101101;
assign F[21][50] = 9'b110101101;
assign F[21][51] = 9'b110101101;
assign F[21][52] = 9'b110101101;
assign F[21][53] = 9'b110101101;
assign F[21][54] = 9'b110101101;
assign F[21][55] = 9'b110101101;
assign F[21][56] = 9'b110101101;
assign F[21][57] = 9'b110101101;
assign F[21][58] = 9'b110101101;
assign F[21][59] = 9'b110101101;
assign F[21][60] = 9'b110101101;
assign F[21][61] = 9'b110101101;
assign F[21][62] = 9'b110101101;
assign F[21][63] = 9'b110001101;
assign F[21][64] = 9'b100100100;
assign F[21][65] = 9'b100000000;
assign F[21][66] = 9'b100100000;
assign F[21][67] = 9'b100100000;
assign F[21][68] = 9'b100100000;
assign F[21][69] = 9'b100000000;
assign F[21][70] = 9'b100000000;
assign F[21][71] = 9'b100000000;
assign F[22][30] = 9'b100100100;
assign F[22][31] = 9'b101000100;
assign F[22][32] = 9'b100100100;
assign F[22][33] = 9'b100100100;
assign F[22][34] = 9'b100100100;
assign F[22][35] = 9'b101000100;
assign F[22][36] = 9'b101000100;
assign F[22][37] = 9'b101000100;
assign F[22][38] = 9'b101101000;
assign F[22][39] = 9'b101101000;
assign F[22][40] = 9'b101101000;
assign F[22][41] = 9'b110101101;
assign F[22][42] = 9'b110110001;
assign F[22][43] = 9'b110101101;
assign F[22][44] = 9'b110101101;
assign F[22][45] = 9'b110101101;
assign F[22][46] = 9'b111110001;
assign F[22][47] = 9'b110101101;
assign F[22][48] = 9'b110101101;
assign F[22][49] = 9'b110101101;
assign F[22][50] = 9'b110101101;
assign F[22][51] = 9'b110101101;
assign F[22][52] = 9'b110101101;
assign F[22][53] = 9'b110101101;
assign F[22][54] = 9'b110101101;
assign F[22][55] = 9'b110101101;
assign F[22][56] = 9'b110101101;
assign F[22][57] = 9'b110101101;
assign F[22][58] = 9'b110101101;
assign F[22][59] = 9'b110101101;
assign F[22][60] = 9'b110101101;
assign F[22][61] = 9'b110101101;
assign F[22][62] = 9'b110101101;
assign F[22][63] = 9'b110101101;
assign F[22][64] = 9'b101000100;
assign F[22][65] = 9'b100000000;
assign F[22][66] = 9'b100100000;
assign F[22][67] = 9'b100100000;
assign F[22][68] = 9'b100100000;
assign F[22][70] = 9'b100000000;
assign F[22][71] = 9'b100000000;
assign F[23][30] = 9'b100100100;
assign F[23][31] = 9'b101000100;
assign F[23][32] = 9'b101000100;
assign F[23][33] = 9'b100100100;
assign F[23][34] = 9'b101000100;
assign F[23][35] = 9'b101000100;
assign F[23][36] = 9'b101000100;
assign F[23][37] = 9'b101101000;
assign F[23][38] = 9'b101101000;
assign F[23][39] = 9'b110001000;
assign F[23][40] = 9'b110101101;
assign F[23][41] = 9'b111110001;
assign F[23][42] = 9'b111110001;
assign F[23][43] = 9'b110101101;
assign F[23][44] = 9'b110101101;
assign F[23][45] = 9'b110101101;
assign F[23][46] = 9'b111110001;
assign F[23][47] = 9'b111110001;
assign F[23][48] = 9'b110101101;
assign F[23][49] = 9'b111110001;
assign F[23][50] = 9'b111110001;
assign F[23][51] = 9'b111110001;
assign F[23][52] = 9'b111110001;
assign F[23][53] = 9'b111110001;
assign F[23][54] = 9'b111110001;
assign F[23][55] = 9'b110101101;
assign F[23][56] = 9'b110101101;
assign F[23][57] = 9'b110101101;
assign F[23][58] = 9'b110101101;
assign F[23][59] = 9'b110101101;
assign F[23][60] = 9'b110101101;
assign F[23][61] = 9'b110101101;
assign F[23][62] = 9'b110101101;
assign F[23][63] = 9'b110101101;
assign F[23][64] = 9'b101101000;
assign F[23][65] = 9'b100100100;
assign F[23][66] = 9'b100000000;
assign F[23][67] = 9'b100100000;
assign F[23][68] = 9'b100100000;
assign F[23][69] = 9'b100100100;
assign F[23][70] = 9'b100000000;
assign F[23][71] = 9'b100000000;
assign F[24][30] = 9'b100100100;
assign F[24][31] = 9'b101000100;
assign F[24][32] = 9'b101000100;
assign F[24][33] = 9'b100100100;
assign F[24][34] = 9'b101000100;
assign F[24][35] = 9'b101000100;
assign F[24][36] = 9'b101101000;
assign F[24][37] = 9'b110001101;
assign F[24][38] = 9'b110001101;
assign F[24][39] = 9'b110101101;
assign F[24][40] = 9'b111110001;
assign F[24][41] = 9'b111110001;
assign F[24][42] = 9'b111110001;
assign F[24][43] = 9'b111110001;
assign F[24][44] = 9'b111110001;
assign F[24][45] = 9'b111110001;
assign F[24][46] = 9'b111110001;
assign F[24][47] = 9'b111110001;
assign F[24][48] = 9'b111110001;
assign F[24][49] = 9'b111110001;
assign F[24][50] = 9'b111110001;
assign F[24][51] = 9'b111110001;
assign F[24][52] = 9'b111110001;
assign F[24][53] = 9'b111110001;
assign F[24][54] = 9'b111110001;
assign F[24][55] = 9'b110101101;
assign F[24][56] = 9'b110101101;
assign F[24][57] = 9'b110101101;
assign F[24][58] = 9'b110101101;
assign F[24][59] = 9'b110101101;
assign F[24][60] = 9'b110101101;
assign F[24][61] = 9'b110101101;
assign F[24][62] = 9'b110101101;
assign F[24][63] = 9'b110101101;
assign F[24][64] = 9'b110001000;
assign F[24][65] = 9'b101000100;
assign F[24][66] = 9'b100000000;
assign F[24][67] = 9'b100100000;
assign F[24][68] = 9'b100000000;
assign F[24][69] = 9'b100000000;
assign F[24][70] = 9'b100000000;
assign F[25][30] = 9'b100100100;
assign F[25][31] = 9'b101000100;
assign F[25][32] = 9'b101000100;
assign F[25][33] = 9'b101000100;
assign F[25][34] = 9'b100100100;
assign F[25][35] = 9'b110001000;
assign F[25][36] = 9'b110101101;
assign F[25][37] = 9'b111110001;
assign F[25][38] = 9'b111110001;
assign F[25][39] = 9'b111110001;
assign F[25][40] = 9'b111110001;
assign F[25][41] = 9'b111110001;
assign F[25][42] = 9'b111110001;
assign F[25][43] = 9'b111110001;
assign F[25][44] = 9'b111110001;
assign F[25][45] = 9'b111110001;
assign F[25][46] = 9'b111110001;
assign F[25][47] = 9'b111110001;
assign F[25][48] = 9'b111110001;
assign F[25][49] = 9'b111110001;
assign F[25][50] = 9'b111110001;
assign F[25][51] = 9'b110101101;
assign F[25][52] = 9'b110101101;
assign F[25][53] = 9'b111110001;
assign F[25][54] = 9'b111110001;
assign F[25][55] = 9'b111110001;
assign F[25][56] = 9'b111110001;
assign F[25][57] = 9'b110101101;
assign F[25][58] = 9'b110101101;
assign F[25][59] = 9'b110101101;
assign F[25][60] = 9'b110101101;
assign F[25][61] = 9'b110101101;
assign F[25][62] = 9'b110101101;
assign F[25][63] = 9'b110101101;
assign F[25][64] = 9'b110001000;
assign F[25][65] = 9'b101000100;
assign F[25][66] = 9'b100000000;
assign F[25][67] = 9'b100100000;
assign F[25][68] = 9'b100100000;
assign F[25][69] = 9'b100000000;
assign F[25][70] = 9'b100000000;
assign F[25][71] = 9'b100000000;
assign F[26][30] = 9'b100100100;
assign F[26][31] = 9'b101000100;
assign F[26][32] = 9'b101000100;
assign F[26][33] = 9'b101000100;
assign F[26][34] = 9'b101101000;
assign F[26][35] = 9'b110101101;
assign F[26][36] = 9'b111110001;
assign F[26][37] = 9'b111110001;
assign F[26][38] = 9'b111110001;
assign F[26][39] = 9'b111110001;
assign F[26][40] = 9'b111110001;
assign F[26][41] = 9'b111110001;
assign F[26][42] = 9'b111110001;
assign F[26][43] = 9'b111110001;
assign F[26][44] = 9'b111110001;
assign F[26][45] = 9'b111110001;
assign F[26][46] = 9'b111110001;
assign F[26][47] = 9'b111110001;
assign F[26][48] = 9'b111110001;
assign F[26][49] = 9'b111110001;
assign F[26][50] = 9'b111110001;
assign F[26][51] = 9'b111110001;
assign F[26][52] = 9'b110001101;
assign F[26][53] = 9'b111110001;
assign F[26][54] = 9'b111110001;
assign F[26][55] = 9'b111110101;
assign F[26][56] = 9'b111110001;
assign F[26][57] = 9'b110101101;
assign F[26][58] = 9'b110101101;
assign F[26][59] = 9'b110101101;
assign F[26][60] = 9'b110101101;
assign F[26][61] = 9'b110101101;
assign F[26][62] = 9'b110101101;
assign F[26][63] = 9'b110101101;
assign F[26][64] = 9'b110101101;
assign F[26][65] = 9'b101101000;
assign F[26][66] = 9'b100000000;
assign F[26][67] = 9'b100100000;
assign F[26][68] = 9'b100100000;
assign F[26][69] = 9'b100100000;
assign F[26][70] = 9'b100000000;
assign F[26][71] = 9'b100000000;
assign F[27][30] = 9'b100100100;
assign F[27][31] = 9'b101000100;
assign F[27][32] = 9'b101000100;
assign F[27][33] = 9'b101000100;
assign F[27][34] = 9'b101000100;
assign F[27][35] = 9'b111110001;
assign F[27][36] = 9'b111110101;
assign F[27][37] = 9'b111110001;
assign F[27][38] = 9'b111110001;
assign F[27][39] = 9'b111110001;
assign F[27][40] = 9'b111110001;
assign F[27][41] = 9'b111110001;
assign F[27][42] = 9'b111110001;
assign F[27][43] = 9'b111110001;
assign F[27][44] = 9'b111110101;
assign F[27][45] = 9'b111110101;
assign F[27][46] = 9'b111110101;
assign F[27][47] = 9'b111110101;
assign F[27][48] = 9'b111110001;
assign F[27][49] = 9'b111110101;
assign F[27][50] = 9'b111110101;
assign F[27][51] = 9'b111110001;
assign F[27][52] = 9'b111110001;
assign F[27][53] = 9'b111110001;
assign F[27][54] = 9'b111110001;
assign F[27][55] = 9'b111110101;
assign F[27][56] = 9'b111110001;
assign F[27][57] = 9'b110101101;
assign F[27][58] = 9'b110001101;
assign F[27][59] = 9'b110001101;
assign F[27][60] = 9'b110001101;
assign F[27][61] = 9'b110001101;
assign F[27][62] = 9'b110001101;
assign F[27][63] = 9'b110001101;
assign F[27][64] = 9'b110101101;
assign F[27][65] = 9'b110001101;
assign F[27][66] = 9'b100000000;
assign F[27][67] = 9'b100100000;
assign F[27][68] = 9'b100100000;
assign F[27][69] = 9'b100100000;
assign F[27][70] = 9'b100000000;
assign F[27][71] = 9'b100000000;
assign F[28][30] = 9'b100100100;
assign F[28][31] = 9'b101000100;
assign F[28][32] = 9'b101000100;
assign F[28][33] = 9'b101000100;
assign F[28][34] = 9'b100100100;
assign F[28][35] = 9'b110101101;
assign F[28][36] = 9'b111110001;
assign F[28][37] = 9'b111110001;
assign F[28][38] = 9'b111110001;
assign F[28][39] = 9'b111110001;
assign F[28][40] = 9'b111110001;
assign F[28][41] = 9'b111110001;
assign F[28][42] = 9'b111110001;
assign F[28][43] = 9'b111110001;
assign F[28][44] = 9'b111110001;
assign F[28][45] = 9'b110110001;
assign F[28][46] = 9'b111110001;
assign F[28][47] = 9'b111110001;
assign F[28][48] = 9'b111110001;
assign F[28][49] = 9'b111110001;
assign F[28][50] = 9'b111110001;
assign F[28][51] = 9'b111110001;
assign F[28][52] = 9'b111110001;
assign F[28][53] = 9'b111110001;
assign F[28][54] = 9'b111110001;
assign F[28][55] = 9'b111110001;
assign F[28][56] = 9'b111110001;
assign F[28][57] = 9'b110001101;
assign F[28][58] = 9'b101101000;
assign F[28][59] = 9'b101000100;
assign F[28][60] = 9'b101000100;
assign F[28][61] = 9'b101000100;
assign F[28][62] = 9'b101000100;
assign F[28][63] = 9'b101000100;
assign F[28][64] = 9'b110001101;
assign F[28][65] = 9'b101101000;
assign F[28][66] = 9'b100000000;
assign F[28][67] = 9'b100100000;
assign F[28][68] = 9'b100100000;
assign F[28][69] = 9'b100100000;
assign F[28][70] = 9'b100000000;
assign F[28][71] = 9'b100000000;
assign F[28][72] = 9'b100000000;
assign F[29][29] = 9'b101000100;
assign F[29][30] = 9'b101000100;
assign F[29][31] = 9'b101000100;
assign F[29][32] = 9'b101000100;
assign F[29][33] = 9'b101000100;
assign F[29][34] = 9'b100100100;
assign F[29][35] = 9'b110001101;
assign F[29][36] = 9'b111110001;
assign F[29][37] = 9'b111110001;
assign F[29][38] = 9'b111110001;
assign F[29][39] = 9'b111110001;
assign F[29][40] = 9'b111110001;
assign F[29][41] = 9'b111110001;
assign F[29][42] = 9'b111110001;
assign F[29][43] = 9'b110001101;
assign F[29][44] = 9'b101101000;
assign F[29][45] = 9'b101000100;
assign F[29][46] = 9'b101101000;
assign F[29][47] = 9'b101101000;
assign F[29][48] = 9'b101101000;
assign F[29][49] = 9'b101100100;
assign F[29][50] = 9'b110001000;
assign F[29][51] = 9'b110101101;
assign F[29][52] = 9'b111110001;
assign F[29][53] = 9'b111110001;
assign F[29][54] = 9'b110101101;
assign F[29][55] = 9'b110001101;
assign F[29][56] = 9'b110001001;
assign F[29][57] = 9'b101101000;
assign F[29][58] = 9'b101000100;
assign F[29][59] = 9'b100100000;
assign F[29][60] = 9'b100100100;
assign F[29][61] = 9'b100100100;
assign F[29][62] = 9'b100100100;
assign F[29][63] = 9'b100100100;
assign F[29][64] = 9'b101001000;
assign F[29][65] = 9'b101000100;
assign F[29][66] = 9'b100100000;
assign F[29][67] = 9'b100000000;
assign F[29][68] = 9'b100000000;
assign F[29][69] = 9'b100000000;
assign F[29][70] = 9'b100100100;
assign F[29][71] = 9'b101000100;
assign F[29][72] = 9'b100000000;
assign F[29][73] = 9'b100000000;
assign F[30][29] = 9'b101000100;
assign F[30][30] = 9'b101000100;
assign F[30][31] = 9'b101000100;
assign F[30][32] = 9'b101000100;
assign F[30][33] = 9'b101000100;
assign F[30][34] = 9'b100100100;
assign F[30][35] = 9'b110001101;
assign F[30][36] = 9'b111110001;
assign F[30][37] = 9'b111110001;
assign F[30][38] = 9'b111110001;
assign F[30][39] = 9'b111110001;
assign F[30][40] = 9'b110101101;
assign F[30][41] = 9'b101101000;
assign F[30][42] = 9'b101101000;
assign F[30][43] = 9'b101101000;
assign F[30][44] = 9'b101101000;
assign F[30][45] = 9'b101001000;
assign F[30][46] = 9'b100100100;
assign F[30][47] = 9'b100100100;
assign F[30][48] = 9'b100100100;
assign F[30][49] = 9'b100100000;
assign F[30][50] = 9'b101000100;
assign F[30][51] = 9'b101101000;
assign F[30][52] = 9'b111110001;
assign F[30][53] = 9'b111110001;
assign F[30][54] = 9'b111110001;
assign F[30][55] = 9'b110001000;
assign F[30][56] = 9'b101000100;
assign F[30][57] = 9'b100100000;
assign F[30][58] = 9'b101001000;
assign F[30][59] = 9'b101101000;
assign F[30][60] = 9'b101101001;
assign F[30][61] = 9'b101101000;
assign F[30][62] = 9'b101101000;
assign F[30][63] = 9'b101101000;
assign F[30][64] = 9'b110001000;
assign F[30][65] = 9'b101101000;
assign F[30][66] = 9'b100100000;
assign F[30][67] = 9'b100100000;
assign F[30][68] = 9'b100000000;
assign F[30][69] = 9'b100000000;
assign F[30][70] = 9'b100100100;
assign F[30][71] = 9'b100100100;
assign F[30][72] = 9'b100000000;
assign F[30][73] = 9'b100000000;
assign F[31][29] = 9'b101000100;
assign F[31][30] = 9'b101000100;
assign F[31][31] = 9'b101000100;
assign F[31][32] = 9'b101000100;
assign F[31][33] = 9'b101000100;
assign F[31][34] = 9'b100100100;
assign F[31][35] = 9'b110001101;
assign F[31][36] = 9'b111110001;
assign F[31][37] = 9'b111110001;
assign F[31][38] = 9'b111110001;
assign F[31][39] = 9'b111110001;
assign F[31][40] = 9'b110001101;
assign F[31][41] = 9'b110001101;
assign F[31][42] = 9'b110001101;
assign F[31][43] = 9'b111110001;
assign F[31][44] = 9'b111110001;
assign F[31][45] = 9'b110110001;
assign F[31][46] = 9'b110001101;
assign F[31][47] = 9'b101101000;
assign F[31][48] = 9'b101001000;
assign F[31][49] = 9'b101000100;
assign F[31][50] = 9'b110001001;
assign F[31][51] = 9'b110101101;
assign F[31][52] = 9'b111110001;
assign F[31][53] = 9'b111110001;
assign F[31][54] = 9'b111110001;
assign F[31][55] = 9'b101101000;
assign F[31][56] = 9'b101000100;
assign F[31][57] = 9'b100100000;
assign F[31][58] = 9'b100100100;
assign F[31][59] = 9'b100100100;
assign F[31][60] = 9'b100100100;
assign F[31][61] = 9'b100100100;
assign F[31][62] = 9'b101000100;
assign F[31][63] = 9'b101101000;
assign F[31][64] = 9'b110001000;
assign F[31][65] = 9'b101101000;
assign F[31][66] = 9'b100100000;
assign F[31][67] = 9'b100100000;
assign F[31][68] = 9'b100100000;
assign F[31][69] = 9'b100100000;
assign F[31][70] = 9'b100000000;
assign F[31][71] = 9'b100000000;
assign F[32][29] = 9'b100100100;
assign F[32][30] = 9'b101000100;
assign F[32][31] = 9'b101000100;
assign F[32][32] = 9'b101000100;
assign F[32][33] = 9'b101000100;
assign F[32][34] = 9'b101000100;
assign F[32][35] = 9'b101101000;
assign F[32][36] = 9'b110001101;
assign F[32][37] = 9'b111110001;
assign F[32][38] = 9'b111110001;
assign F[32][39] = 9'b111110001;
assign F[32][40] = 9'b111110001;
assign F[32][41] = 9'b111110001;
assign F[32][42] = 9'b111110001;
assign F[32][43] = 9'b110101101;
assign F[32][44] = 9'b101101000;
assign F[32][45] = 9'b101000100;
assign F[32][46] = 9'b101000100;
assign F[32][47] = 9'b101001000;
assign F[32][48] = 9'b101101000;
assign F[32][49] = 9'b101101000;
assign F[32][50] = 9'b110001101;
assign F[32][51] = 9'b110101101;
assign F[32][52] = 9'b111110001;
assign F[32][53] = 9'b111110001;
assign F[32][54] = 9'b111110001;
assign F[32][55] = 9'b110101101;
assign F[32][56] = 9'b101101000;
assign F[32][57] = 9'b100100000;
assign F[32][58] = 9'b100100100;
assign F[32][59] = 9'b100100100;
assign F[32][60] = 9'b100100000;
assign F[32][61] = 9'b100100000;
assign F[32][62] = 9'b100100000;
assign F[32][63] = 9'b100100100;
assign F[32][64] = 9'b101101000;
assign F[32][65] = 9'b101101000;
assign F[32][66] = 9'b100100000;
assign F[32][67] = 9'b100100000;
assign F[32][68] = 9'b100100000;
assign F[32][69] = 9'b100100000;
assign F[32][70] = 9'b100000000;
assign F[32][71] = 9'b100000000;
assign F[33][29] = 9'b100100100;
assign F[33][30] = 9'b100100100;
assign F[33][31] = 9'b101000100;
assign F[33][32] = 9'b101000100;
assign F[33][33] = 9'b101000100;
assign F[33][34] = 9'b101000100;
assign F[33][35] = 9'b101101000;
assign F[33][36] = 9'b110001101;
assign F[33][37] = 9'b111110101;
assign F[33][38] = 9'b111110001;
assign F[33][39] = 9'b111110001;
assign F[33][40] = 9'b111110001;
assign F[33][41] = 9'b111110001;
assign F[33][42] = 9'b110101101;
assign F[33][43] = 9'b110001101;
assign F[33][44] = 9'b101101000;
assign F[33][45] = 9'b101001000;
assign F[33][46] = 9'b101000100;
assign F[33][47] = 9'b101001000;
assign F[33][48] = 9'b101101000;
assign F[33][49] = 9'b101101000;
assign F[33][50] = 9'b110001101;
assign F[33][51] = 9'b110101101;
assign F[33][52] = 9'b111110001;
assign F[33][53] = 9'b111110001;
assign F[33][54] = 9'b111110001;
assign F[33][55] = 9'b111110001;
assign F[33][56] = 9'b101101000;
assign F[33][57] = 9'b100100000;
assign F[33][58] = 9'b100100100;
assign F[33][59] = 9'b101000100;
assign F[33][60] = 9'b101000100;
assign F[33][61] = 9'b101000100;
assign F[33][62] = 9'b101000100;
assign F[33][63] = 9'b101000100;
assign F[33][64] = 9'b101101000;
assign F[33][65] = 9'b101101000;
assign F[33][66] = 9'b101000100;
assign F[33][67] = 9'b100100000;
assign F[33][68] = 9'b100100000;
assign F[33][69] = 9'b100100000;
assign F[33][70] = 9'b100000000;
assign F[33][71] = 9'b100000000;
assign F[34][30] = 9'b100100100;
assign F[34][31] = 9'b101000100;
assign F[34][32] = 9'b101000100;
assign F[34][33] = 9'b101000100;
assign F[34][34] = 9'b100100100;
assign F[34][35] = 9'b101000100;
assign F[34][36] = 9'b110001101;
assign F[34][37] = 9'b111110101;
assign F[34][38] = 9'b111110001;
assign F[34][39] = 9'b111110001;
assign F[34][40] = 9'b111110001;
assign F[34][41] = 9'b111110001;
assign F[34][42] = 9'b110110001;
assign F[34][43] = 9'b111110001;
assign F[34][44] = 9'b111110001;
assign F[34][45] = 9'b111110001;
assign F[34][46] = 9'b110001101;
assign F[34][47] = 9'b110001101;
assign F[34][48] = 9'b110001001;
assign F[34][49] = 9'b110001000;
assign F[34][50] = 9'b110001101;
assign F[34][51] = 9'b111110001;
assign F[34][52] = 9'b111110001;
assign F[34][53] = 9'b111110001;
assign F[34][54] = 9'b111110001;
assign F[34][55] = 9'b111101101;
assign F[34][56] = 9'b110001001;
assign F[34][57] = 9'b101000100;
assign F[34][58] = 9'b101000100;
assign F[34][59] = 9'b101101000;
assign F[34][60] = 9'b101101000;
assign F[34][61] = 9'b101101000;
assign F[34][62] = 9'b101101000;
assign F[34][63] = 9'b101101000;
assign F[34][64] = 9'b110001000;
assign F[34][65] = 9'b110001000;
assign F[34][66] = 9'b101101000;
assign F[34][67] = 9'b100100100;
assign F[34][68] = 9'b100000000;
assign F[34][69] = 9'b100000000;
assign F[34][70] = 9'b100000000;
assign F[34][71] = 9'b100000000;
assign F[35][30] = 9'b100100100;
assign F[35][31] = 9'b101000100;
assign F[35][32] = 9'b101000100;
assign F[35][33] = 9'b101000100;
assign F[35][34] = 9'b101000100;
assign F[35][35] = 9'b101000100;
assign F[35][36] = 9'b110001001;
assign F[35][37] = 9'b111110101;
assign F[35][38] = 9'b111110001;
assign F[35][39] = 9'b111110001;
assign F[35][40] = 9'b111110001;
assign F[35][41] = 9'b111110001;
assign F[35][42] = 9'b111110001;
assign F[35][43] = 9'b111110001;
assign F[35][44] = 9'b111110001;
assign F[35][45] = 9'b111110001;
assign F[35][46] = 9'b111110101;
assign F[35][47] = 9'b111110001;
assign F[35][48] = 9'b110101101;
assign F[35][49] = 9'b110110001;
assign F[35][50] = 9'b111110001;
assign F[35][51] = 9'b111110001;
assign F[35][52] = 9'b111110001;
assign F[35][53] = 9'b111110001;
assign F[35][54] = 9'b111110001;
assign F[35][55] = 9'b110101101;
assign F[35][56] = 9'b110001101;
assign F[35][57] = 9'b101101000;
assign F[35][58] = 9'b101101000;
assign F[35][59] = 9'b101101000;
assign F[35][60] = 9'b101101000;
assign F[35][61] = 9'b101101000;
assign F[35][62] = 9'b101101000;
assign F[35][63] = 9'b101101000;
assign F[35][64] = 9'b110001101;
assign F[35][65] = 9'b110101101;
assign F[35][66] = 9'b110001001;
assign F[35][67] = 9'b101000100;
assign F[35][68] = 9'b100000000;
assign F[35][69] = 9'b100000000;
assign F[36][30] = 9'b101000100;
assign F[36][31] = 9'b101000100;
assign F[36][32] = 9'b101101000;
assign F[36][33] = 9'b101101000;
assign F[36][34] = 9'b101101000;
assign F[36][35] = 9'b101101000;
assign F[36][36] = 9'b110001001;
assign F[36][37] = 9'b111110101;
assign F[36][38] = 9'b111110001;
assign F[36][39] = 9'b111110001;
assign F[36][40] = 9'b111110001;
assign F[36][41] = 9'b111110001;
assign F[36][42] = 9'b111110001;
assign F[36][43] = 9'b111110001;
assign F[36][44] = 9'b111110001;
assign F[36][45] = 9'b111110001;
assign F[36][46] = 9'b111110001;
assign F[36][47] = 9'b111110001;
assign F[36][48] = 9'b111110001;
assign F[36][49] = 9'b111110001;
assign F[36][50] = 9'b111110001;
assign F[36][51] = 9'b111110001;
assign F[36][52] = 9'b111110001;
assign F[36][53] = 9'b111110001;
assign F[36][54] = 9'b111110001;
assign F[36][55] = 9'b110101101;
assign F[36][56] = 9'b110001101;
assign F[36][57] = 9'b101101000;
assign F[36][58] = 9'b101101000;
assign F[36][59] = 9'b101101000;
assign F[36][60] = 9'b101101000;
assign F[36][61] = 9'b101101000;
assign F[36][62] = 9'b101101000;
assign F[36][63] = 9'b101101000;
assign F[36][64] = 9'b110001101;
assign F[36][65] = 9'b110101101;
assign F[36][66] = 9'b110110001;
assign F[36][67] = 9'b101000100;
assign F[36][68] = 9'b100000000;
assign F[36][69] = 9'b100000000;
assign F[36][70] = 9'b100000000;
assign F[37][30] = 9'b101101001;
assign F[37][31] = 9'b101101000;
assign F[37][32] = 9'b110001101;
assign F[37][33] = 9'b110001101;
assign F[37][34] = 9'b110101101;
assign F[37][35] = 9'b101101000;
assign F[37][36] = 9'b101101000;
assign F[37][37] = 9'b111110101;
assign F[37][38] = 9'b111110001;
assign F[37][39] = 9'b111110001;
assign F[37][40] = 9'b111110001;
assign F[37][41] = 9'b111110001;
assign F[37][42] = 9'b111110001;
assign F[37][43] = 9'b111110001;
assign F[37][44] = 9'b111110001;
assign F[37][45] = 9'b111110001;
assign F[37][46] = 9'b111110001;
assign F[37][47] = 9'b111110001;
assign F[37][48] = 9'b111110001;
assign F[37][49] = 9'b111110001;
assign F[37][50] = 9'b111110001;
assign F[37][51] = 9'b111110001;
assign F[37][52] = 9'b111110001;
assign F[37][53] = 9'b111110001;
assign F[37][54] = 9'b111110001;
assign F[37][55] = 9'b110101101;
assign F[37][56] = 9'b110101101;
assign F[37][57] = 9'b110101101;
assign F[37][58] = 9'b101101000;
assign F[37][59] = 9'b101101000;
assign F[37][60] = 9'b101101000;
assign F[37][61] = 9'b101101000;
assign F[37][62] = 9'b101101000;
assign F[37][63] = 9'b101101000;
assign F[37][64] = 9'b110001101;
assign F[37][65] = 9'b110101101;
assign F[37][66] = 9'b110101101;
assign F[37][67] = 9'b101000100;
assign F[37][68] = 9'b100000000;
assign F[37][69] = 9'b100000000;
assign F[37][70] = 9'b100000000;
assign F[38][32] = 9'b110101101;
assign F[38][33] = 9'b111101101;
assign F[38][34] = 9'b110101101;
assign F[38][35] = 9'b110001101;
assign F[38][36] = 9'b110001101;
assign F[38][37] = 9'b110101101;
assign F[38][38] = 9'b111110001;
assign F[38][39] = 9'b111110001;
assign F[38][40] = 9'b111110001;
assign F[38][41] = 9'b111110001;
assign F[38][42] = 9'b111110001;
assign F[38][43] = 9'b111110001;
assign F[38][44] = 9'b111110001;
assign F[38][45] = 9'b111110001;
assign F[38][46] = 9'b111110001;
assign F[38][47] = 9'b111110001;
assign F[38][48] = 9'b111110001;
assign F[38][49] = 9'b111110001;
assign F[38][50] = 9'b111110001;
assign F[38][51] = 9'b111110001;
assign F[38][52] = 9'b111110101;
assign F[38][53] = 9'b111110101;
assign F[38][54] = 9'b111110101;
assign F[38][55] = 9'b111110001;
assign F[38][56] = 9'b111110001;
assign F[38][57] = 9'b110101101;
assign F[38][58] = 9'b110101101;
assign F[38][59] = 9'b110001101;
assign F[38][60] = 9'b101101000;
assign F[38][61] = 9'b110001101;
assign F[38][62] = 9'b110001101;
assign F[38][63] = 9'b110001101;
assign F[38][64] = 9'b110101101;
assign F[38][65] = 9'b110101101;
assign F[38][66] = 9'b110101101;
assign F[38][67] = 9'b101000100;
assign F[38][68] = 9'b100000000;
assign F[38][69] = 9'b100000000;
assign F[38][70] = 9'b100000000;
assign F[39][32] = 9'b101101001;
assign F[39][33] = 9'b110001001;
assign F[39][34] = 9'b101101000;
assign F[39][35] = 9'b110001101;
assign F[39][36] = 9'b110001101;
assign F[39][37] = 9'b101101000;
assign F[39][38] = 9'b111110001;
assign F[39][39] = 9'b111110101;
assign F[39][40] = 9'b111110001;
assign F[39][41] = 9'b111110001;
assign F[39][42] = 9'b111110001;
assign F[39][43] = 9'b111110001;
assign F[39][44] = 9'b111110001;
assign F[39][45] = 9'b111110001;
assign F[39][46] = 9'b111110001;
assign F[39][47] = 9'b111110001;
assign F[39][48] = 9'b111110001;
assign F[39][49] = 9'b111110001;
assign F[39][50] = 9'b111110001;
assign F[39][51] = 9'b111110001;
assign F[39][52] = 9'b110001101;
assign F[39][53] = 9'b110001101;
assign F[39][54] = 9'b110001101;
assign F[39][55] = 9'b111110001;
assign F[39][56] = 9'b110101101;
assign F[39][57] = 9'b110001000;
assign F[39][58] = 9'b110001001;
assign F[39][59] = 9'b101101000;
assign F[39][60] = 9'b101101000;
assign F[39][61] = 9'b110001101;
assign F[39][62] = 9'b110001101;
assign F[39][63] = 9'b110001000;
assign F[39][64] = 9'b110001101;
assign F[39][65] = 9'b110101101;
assign F[39][66] = 9'b110101101;
assign F[39][67] = 9'b101000100;
assign F[39][68] = 9'b100100000;
assign F[39][69] = 9'b100000000;
assign F[39][70] = 9'b100000000;
assign F[40][32] = 9'b101001000;
assign F[40][33] = 9'b110001001;
assign F[40][34] = 9'b110101101;
assign F[40][35] = 9'b111110001;
assign F[40][36] = 9'b110001101;
assign F[40][37] = 9'b101000100;
assign F[40][38] = 9'b110001101;
assign F[40][39] = 9'b111110001;
assign F[40][40] = 9'b111110001;
assign F[40][41] = 9'b111110001;
assign F[40][42] = 9'b111110001;
assign F[40][43] = 9'b111110001;
assign F[40][44] = 9'b111110001;
assign F[40][45] = 9'b111110001;
assign F[40][46] = 9'b111110001;
assign F[40][47] = 9'b111110001;
assign F[40][48] = 9'b111110001;
assign F[40][49] = 9'b111110001;
assign F[40][50] = 9'b111110001;
assign F[40][51] = 9'b111110001;
assign F[40][52] = 9'b110001101;
assign F[40][53] = 9'b110001000;
assign F[40][54] = 9'b110001001;
assign F[40][55] = 9'b110001101;
assign F[40][56] = 9'b110001000;
assign F[40][57] = 9'b101101000;
assign F[40][58] = 9'b101000100;
assign F[40][59] = 9'b101000100;
assign F[40][60] = 9'b101101000;
assign F[40][61] = 9'b110001101;
assign F[40][62] = 9'b110101101;
assign F[40][63] = 9'b110001000;
assign F[40][64] = 9'b110001101;
assign F[40][65] = 9'b110101101;
assign F[40][66] = 9'b110101101;
assign F[40][67] = 9'b101000100;
assign F[40][68] = 9'b100000000;
assign F[40][69] = 9'b100000000;
assign F[41][34] = 9'b111111110;
assign F[41][35] = 9'b111110101;
assign F[41][36] = 9'b111110001;
assign F[41][37] = 9'b101101000;
assign F[41][38] = 9'b110001101;
assign F[41][39] = 9'b110101101;
assign F[41][40] = 9'b111110001;
assign F[41][41] = 9'b111110001;
assign F[41][42] = 9'b111110001;
assign F[41][43] = 9'b111110001;
assign F[41][44] = 9'b111110001;
assign F[41][45] = 9'b111110001;
assign F[41][46] = 9'b111110001;
assign F[41][47] = 9'b111110001;
assign F[41][48] = 9'b111110001;
assign F[41][49] = 9'b111110001;
assign F[41][50] = 9'b111110001;
assign F[41][51] = 9'b111110001;
assign F[41][52] = 9'b110101101;
assign F[41][53] = 9'b110101101;
assign F[41][54] = 9'b110101101;
assign F[41][55] = 9'b101101000;
assign F[41][56] = 9'b101101000;
assign F[41][57] = 9'b101101000;
assign F[41][58] = 9'b101000100;
assign F[41][59] = 9'b101000100;
assign F[41][60] = 9'b101101000;
assign F[41][61] = 9'b110001101;
assign F[41][62] = 9'b110001101;
assign F[41][63] = 9'b110101101;
assign F[41][64] = 9'b110101101;
assign F[41][65] = 9'b110101101;
assign F[41][66] = 9'b111110001;
assign F[41][67] = 9'b100100100;
assign F[41][68] = 9'b100000000;
assign F[42][34] = 9'b111110101;
assign F[42][35] = 9'b111110001;
assign F[42][36] = 9'b111110001;
assign F[42][37] = 9'b110101101;
assign F[42][38] = 9'b110101101;
assign F[42][39] = 9'b110101101;
assign F[42][40] = 9'b111110001;
assign F[42][41] = 9'b111110001;
assign F[42][42] = 9'b111110001;
assign F[42][43] = 9'b111110001;
assign F[42][44] = 9'b111110001;
assign F[42][45] = 9'b111110001;
assign F[42][46] = 9'b111110001;
assign F[42][47] = 9'b111110001;
assign F[42][48] = 9'b111110001;
assign F[42][49] = 9'b111110001;
assign F[42][50] = 9'b111110001;
assign F[42][51] = 9'b110001101;
assign F[42][52] = 9'b110101101;
assign F[42][53] = 9'b110101101;
assign F[42][54] = 9'b110101101;
assign F[42][55] = 9'b101101000;
assign F[42][56] = 9'b101101000;
assign F[42][57] = 9'b101101000;
assign F[42][58] = 9'b101000100;
assign F[42][59] = 9'b101000100;
assign F[42][60] = 9'b101000100;
assign F[42][61] = 9'b101001000;
assign F[42][62] = 9'b101101000;
assign F[42][63] = 9'b110101101;
assign F[42][64] = 9'b110101101;
assign F[42][65] = 9'b110101101;
assign F[42][66] = 9'b110110001;
assign F[42][67] = 9'b100100100;
assign F[42][68] = 9'b100000000;
assign F[43][35] = 9'b111110001;
assign F[43][36] = 9'b111110101;
assign F[43][37] = 9'b111110001;
assign F[43][38] = 9'b110101101;
assign F[43][39] = 9'b110101101;
assign F[43][40] = 9'b111110001;
assign F[43][41] = 9'b111110001;
assign F[43][42] = 9'b111110001;
assign F[43][43] = 9'b111110001;
assign F[43][44] = 9'b111110001;
assign F[43][45] = 9'b111110001;
assign F[43][46] = 9'b111110001;
assign F[43][47] = 9'b111110001;
assign F[43][48] = 9'b110001101;
assign F[43][49] = 9'b110101101;
assign F[43][50] = 9'b110101101;
assign F[43][51] = 9'b110101101;
assign F[43][52] = 9'b110101101;
assign F[43][53] = 9'b110101101;
assign F[43][54] = 9'b110101101;
assign F[43][55] = 9'b101101000;
assign F[43][56] = 9'b110001001;
assign F[43][57] = 9'b110101101;
assign F[43][58] = 9'b101101000;
assign F[43][59] = 9'b101101000;
assign F[43][60] = 9'b101101000;
assign F[43][61] = 9'b101000100;
assign F[43][62] = 9'b101000100;
assign F[43][63] = 9'b101101000;
assign F[43][64] = 9'b110101101;
assign F[43][65] = 9'b110101101;
assign F[44][36] = 9'b111110101;
assign F[44][37] = 9'b111110101;
assign F[44][38] = 9'b110101101;
assign F[44][39] = 9'b110101101;
assign F[44][40] = 9'b111110001;
assign F[44][41] = 9'b111110001;
assign F[44][42] = 9'b111110001;
assign F[44][43] = 9'b111110001;
assign F[44][44] = 9'b111110001;
assign F[44][45] = 9'b111110001;
assign F[44][46] = 9'b111110001;
assign F[44][47] = 9'b111110001;
assign F[44][48] = 9'b110001101;
assign F[44][49] = 9'b110101101;
assign F[44][50] = 9'b110101101;
assign F[44][51] = 9'b110101101;
assign F[44][52] = 9'b110101101;
assign F[44][53] = 9'b110101101;
assign F[44][54] = 9'b110101101;
assign F[44][55] = 9'b110101101;
assign F[44][56] = 9'b110001101;
assign F[44][57] = 9'b101101000;
assign F[44][58] = 9'b101101000;
assign F[44][59] = 9'b101101000;
assign F[44][60] = 9'b101101000;
assign F[44][61] = 9'b101000100;
assign F[44][62] = 9'b101000100;
assign F[44][63] = 9'b101101000;
assign F[44][64] = 9'b110001000;
assign F[44][65] = 9'b101101000;
assign F[45][37] = 9'b110110001;
assign F[45][38] = 9'b110101101;
assign F[45][39] = 9'b110101101;
assign F[45][40] = 9'b111110001;
assign F[45][41] = 9'b111110001;
assign F[45][42] = 9'b111110001;
assign F[45][43] = 9'b111110001;
assign F[45][44] = 9'b111110001;
assign F[45][45] = 9'b111110001;
assign F[45][46] = 9'b111110001;
assign F[45][47] = 9'b110001101;
assign F[45][48] = 9'b101101000;
assign F[45][49] = 9'b101101000;
assign F[45][50] = 9'b110001101;
assign F[45][51] = 9'b110101101;
assign F[45][52] = 9'b110101101;
assign F[45][53] = 9'b110101101;
assign F[45][54] = 9'b110101101;
assign F[45][55] = 9'b110101101;
assign F[45][56] = 9'b110001101;
assign F[45][57] = 9'b101101000;
assign F[45][58] = 9'b101101000;
assign F[45][59] = 9'b101101000;
assign F[45][60] = 9'b101101000;
assign F[45][61] = 9'b101000100;
assign F[45][62] = 9'b101000100;
assign F[45][63] = 9'b101101000;
assign F[45][64] = 9'b101101000;
assign F[45][65] = 9'b101101000;
assign F[46][37] = 9'b111110001;
assign F[46][38] = 9'b111110001;
assign F[46][39] = 9'b111110001;
assign F[46][40] = 9'b111110001;
assign F[46][41] = 9'b111110001;
assign F[46][42] = 9'b111110001;
assign F[46][43] = 9'b111110001;
assign F[46][44] = 9'b111110001;
assign F[46][45] = 9'b111110001;
assign F[46][46] = 9'b110101101;
assign F[46][47] = 9'b110001101;
assign F[46][48] = 9'b110001101;
assign F[46][49] = 9'b110001001;
assign F[46][50] = 9'b110001101;
assign F[46][51] = 9'b110101101;
assign F[46][52] = 9'b111110001;
assign F[46][53] = 9'b111110001;
assign F[46][54] = 9'b111110001;
assign F[46][55] = 9'b110101101;
assign F[46][56] = 9'b110001101;
assign F[46][57] = 9'b110001101;
assign F[46][58] = 9'b101101000;
assign F[46][59] = 9'b101101000;
assign F[46][60] = 9'b101101000;
assign F[46][61] = 9'b101000100;
assign F[46][62] = 9'b101001000;
assign F[46][63] = 9'b101101000;
assign F[46][64] = 9'b101101000;
assign F[46][65] = 9'b101101000;
assign F[47][37] = 9'b111110001;
assign F[47][38] = 9'b111110001;
assign F[47][39] = 9'b111110001;
assign F[47][40] = 9'b111110001;
assign F[47][41] = 9'b111110001;
assign F[47][42] = 9'b111110001;
assign F[47][43] = 9'b111110001;
assign F[47][44] = 9'b111110001;
assign F[47][45] = 9'b111110001;
assign F[47][46] = 9'b111110001;
assign F[47][47] = 9'b110101101;
assign F[47][48] = 9'b110101101;
assign F[47][49] = 9'b111110001;
assign F[47][50] = 9'b111110001;
assign F[47][51] = 9'b111110001;
assign F[47][52] = 9'b111110001;
assign F[47][53] = 9'b111110001;
assign F[47][54] = 9'b111110001;
assign F[47][55] = 9'b110001101;
assign F[47][56] = 9'b110001101;
assign F[47][57] = 9'b110001101;
assign F[47][58] = 9'b101101000;
assign F[47][59] = 9'b101101000;
assign F[47][60] = 9'b101101000;
assign F[47][61] = 9'b110001101;
assign F[47][62] = 9'b110001101;
assign F[47][63] = 9'b101101000;
assign F[47][64] = 9'b101101000;
assign F[47][65] = 9'b101101000;
assign F[48][37] = 9'b111101101;
assign F[48][38] = 9'b111110001;
assign F[48][39] = 9'b111110001;
assign F[48][40] = 9'b110001101;
assign F[48][41] = 9'b110101101;
assign F[48][42] = 9'b110101101;
assign F[48][43] = 9'b111110001;
assign F[48][44] = 9'b111110001;
assign F[48][45] = 9'b111110001;
assign F[48][46] = 9'b111110101;
assign F[48][47] = 9'b111110001;
assign F[48][48] = 9'b110101101;
assign F[48][49] = 9'b111110001;
assign F[48][50] = 9'b111110001;
assign F[48][51] = 9'b111110001;
assign F[48][52] = 9'b111110001;
assign F[48][53] = 9'b111110001;
assign F[48][54] = 9'b110101101;
assign F[48][55] = 9'b110001000;
assign F[48][56] = 9'b101101000;
assign F[48][57] = 9'b101101000;
assign F[48][58] = 9'b101101000;
assign F[48][59] = 9'b110001001;
assign F[48][60] = 9'b110001001;
assign F[48][61] = 9'b110001101;
assign F[48][62] = 9'b110001101;
assign F[48][63] = 9'b101101000;
assign F[48][64] = 9'b101101000;
assign F[48][65] = 9'b101101000;
assign F[49][37] = 9'b111110101;
assign F[49][38] = 9'b111110001;
assign F[49][39] = 9'b111110001;
assign F[49][40] = 9'b110101101;
assign F[49][41] = 9'b110101101;
assign F[49][42] = 9'b110101101;
assign F[49][43] = 9'b111110001;
assign F[49][44] = 9'b111110001;
assign F[49][45] = 9'b111110001;
assign F[49][46] = 9'b111110001;
assign F[49][47] = 9'b111110001;
assign F[49][48] = 9'b111110001;
assign F[49][49] = 9'b111110001;
assign F[49][50] = 9'b111110001;
assign F[49][51] = 9'b111110001;
assign F[49][52] = 9'b111110001;
assign F[49][53] = 9'b111110001;
assign F[49][54] = 9'b111110001;
assign F[49][55] = 9'b110110001;
assign F[49][56] = 9'b110001101;
assign F[49][57] = 9'b101101000;
assign F[49][58] = 9'b110001101;
assign F[49][59] = 9'b110001101;
assign F[49][60] = 9'b110001101;
assign F[49][61] = 9'b101101000;
assign F[49][62] = 9'b101101000;
assign F[49][63] = 9'b101101000;
assign F[50][37] = 9'b111110101;
assign F[50][38] = 9'b111110001;
assign F[50][39] = 9'b111110001;
assign F[50][40] = 9'b111110001;
assign F[50][41] = 9'b111110001;
assign F[50][42] = 9'b110101101;
assign F[50][43] = 9'b110101101;
assign F[50][44] = 9'b111110001;
assign F[50][45] = 9'b111110001;
assign F[50][46] = 9'b111110001;
assign F[50][47] = 9'b111110001;
assign F[50][48] = 9'b111110001;
assign F[50][49] = 9'b111110001;
assign F[50][50] = 9'b111110001;
assign F[50][51] = 9'b111110001;
assign F[50][52] = 9'b111110001;
assign F[50][53] = 9'b111110001;
assign F[50][54] = 9'b111110001;
assign F[50][55] = 9'b110101101;
assign F[50][56] = 9'b110101101;
assign F[50][57] = 9'b110101101;
assign F[50][58] = 9'b110001000;
assign F[50][59] = 9'b101101000;
assign F[50][60] = 9'b101101000;
assign F[50][61] = 9'b101101000;
assign F[50][62] = 9'b101101000;
assign F[50][63] = 9'b101101000;
assign F[51][37] = 9'b111110101;
assign F[51][38] = 9'b111110001;
assign F[51][39] = 9'b111110001;
assign F[51][40] = 9'b111110001;
assign F[51][41] = 9'b111110001;
assign F[51][42] = 9'b111110001;
assign F[51][43] = 9'b111110001;
assign F[51][44] = 9'b111110001;
assign F[51][45] = 9'b111110001;
assign F[51][46] = 9'b111110001;
assign F[51][47] = 9'b111110001;
assign F[51][48] = 9'b111110001;
assign F[51][49] = 9'b110101101;
assign F[51][50] = 9'b111110001;
assign F[51][51] = 9'b111110001;
assign F[51][52] = 9'b111110001;
assign F[51][53] = 9'b111110001;
assign F[51][54] = 9'b110101101;
assign F[51][55] = 9'b110101101;
assign F[51][56] = 9'b110101101;
assign F[51][57] = 9'b110101101;
assign F[51][58] = 9'b101101000;
assign F[51][59] = 9'b101101000;
assign F[51][60] = 9'b101101000;
assign F[51][61] = 9'b101101000;
assign F[51][62] = 9'b101101000;
assign F[52][34] = 9'b100000000;
assign F[52][35] = 9'b100000000;
assign F[52][36] = 9'b101101000;
assign F[52][37] = 9'b111110001;
assign F[52][38] = 9'b111110001;
assign F[52][39] = 9'b111110001;
assign F[52][40] = 9'b111110001;
assign F[52][41] = 9'b111110001;
assign F[52][42] = 9'b111110001;
assign F[52][43] = 9'b111110001;
assign F[52][44] = 9'b111110001;
assign F[52][45] = 9'b111110001;
assign F[52][46] = 9'b110101101;
assign F[52][47] = 9'b111110001;
assign F[52][48] = 9'b111101101;
assign F[52][49] = 9'b110101101;
assign F[52][50] = 9'b110101101;
assign F[52][51] = 9'b111110001;
assign F[52][52] = 9'b111110001;
assign F[52][53] = 9'b111110001;
assign F[52][54] = 9'b111110001;
assign F[52][55] = 9'b110101101;
assign F[52][56] = 9'b110101101;
assign F[52][57] = 9'b110101101;
assign F[52][58] = 9'b101101000;
assign F[52][59] = 9'b101101000;
assign F[52][60] = 9'b101101000;
assign F[52][61] = 9'b101101001;
assign F[52][62] = 9'b101101000;
assign F[53][32] = 9'b100000000;
assign F[53][33] = 9'b100000000;
assign F[53][34] = 9'b100000000;
assign F[53][35] = 9'b100100000;
assign F[53][36] = 9'b101000100;
assign F[53][37] = 9'b110001101;
assign F[53][38] = 9'b110110001;
assign F[53][39] = 9'b111110001;
assign F[53][40] = 9'b111110101;
assign F[53][41] = 9'b111110001;
assign F[53][42] = 9'b111110001;
assign F[53][43] = 9'b111110001;
assign F[53][44] = 9'b111110001;
assign F[53][45] = 9'b111110001;
assign F[53][46] = 9'b111110001;
assign F[53][47] = 9'b110101101;
assign F[53][48] = 9'b110001101;
assign F[53][49] = 9'b110101101;
assign F[53][50] = 9'b110101101;
assign F[53][51] = 9'b110101101;
assign F[53][52] = 9'b111110001;
assign F[53][53] = 9'b111110001;
assign F[53][54] = 9'b111110001;
assign F[53][55] = 9'b110101101;
assign F[53][56] = 9'b110001101;
assign F[53][57] = 9'b110001001;
assign F[53][58] = 9'b101101000;
assign F[53][59] = 9'b101101000;
assign F[53][60] = 9'b101101000;
assign F[53][61] = 9'b101101000;
assign F[53][62] = 9'b101101001;
assign F[54][32] = 9'b100000000;
assign F[54][33] = 9'b100000000;
assign F[54][34] = 9'b100100100;
assign F[54][35] = 9'b100000000;
assign F[54][36] = 9'b100100100;
assign F[54][37] = 9'b101000100;
assign F[54][38] = 9'b101101000;
assign F[54][39] = 9'b110001101;
assign F[54][40] = 9'b111110001;
assign F[54][41] = 9'b111110001;
assign F[54][42] = 9'b111110101;
assign F[54][43] = 9'b111110001;
assign F[54][44] = 9'b111110001;
assign F[54][45] = 9'b111110001;
assign F[54][46] = 9'b111110001;
assign F[54][47] = 9'b111110001;
assign F[54][48] = 9'b110101101;
assign F[54][49] = 9'b110101101;
assign F[54][50] = 9'b110101101;
assign F[54][51] = 9'b110001101;
assign F[54][52] = 9'b110001101;
assign F[54][53] = 9'b110001101;
assign F[54][54] = 9'b110001101;
assign F[54][55] = 9'b110001101;
assign F[54][56] = 9'b110001001;
assign F[54][57] = 9'b101101000;
assign F[54][58] = 9'b101101000;
assign F[54][59] = 9'b101101000;
assign F[54][60] = 9'b101101000;
assign F[55][32] = 9'b100000000;
assign F[55][33] = 9'b100000000;
assign F[55][34] = 9'b100100100;
assign F[55][35] = 9'b100000000;
assign F[55][36] = 9'b100000000;
assign F[55][37] = 9'b100000000;
assign F[55][38] = 9'b100100000;
assign F[55][39] = 9'b100100100;
assign F[55][40] = 9'b101000100;
assign F[55][41] = 9'b110001101;
assign F[55][42] = 9'b111110001;
assign F[55][43] = 9'b111110001;
assign F[55][44] = 9'b111110001;
assign F[55][45] = 9'b111110001;
assign F[55][46] = 9'b111110001;
assign F[55][47] = 9'b111110001;
assign F[55][48] = 9'b111110001;
assign F[55][49] = 9'b110101101;
assign F[55][50] = 9'b110101101;
assign F[55][51] = 9'b110101101;
assign F[55][52] = 9'b110001000;
assign F[55][53] = 9'b101101000;
assign F[55][54] = 9'b101101000;
assign F[55][55] = 9'b101101000;
assign F[55][56] = 9'b101101000;
assign F[55][57] = 9'b101101000;
assign F[55][58] = 9'b101101000;
assign F[55][59] = 9'b101101000;
assign F[55][60] = 9'b101101001;
assign F[55][61] = 9'b101101000;
assign F[56][32] = 9'b100000000;
assign F[56][33] = 9'b100000000;
assign F[56][34] = 9'b100100100;
assign F[56][35] = 9'b100000000;
assign F[56][36] = 9'b100000000;
assign F[56][37] = 9'b100000000;
assign F[56][38] = 9'b100000000;
assign F[56][39] = 9'b100000000;
assign F[56][40] = 9'b100000000;
assign F[56][41] = 9'b100000000;
assign F[56][42] = 9'b100100100;
assign F[56][43] = 9'b101101000;
assign F[56][44] = 9'b110101101;
assign F[56][45] = 9'b111110001;
assign F[56][46] = 9'b111110001;
assign F[56][47] = 9'b111110001;
assign F[56][48] = 9'b111110001;
assign F[56][49] = 9'b111110001;
assign F[56][50] = 9'b111110001;
assign F[56][51] = 9'b111110001;
assign F[56][52] = 9'b111110001;
assign F[56][53] = 9'b111110001;
assign F[56][54] = 9'b110101101;
assign F[56][55] = 9'b110101101;
assign F[56][56] = 9'b110101101;
assign F[56][57] = 9'b110101101;
assign F[56][58] = 9'b110101101;
assign F[56][59] = 9'b110101101;
assign F[56][60] = 9'b110101101;
assign F[56][61] = 9'b110001000;
assign F[56][62] = 9'b101000100;
assign F[56][63] = 9'b100000000;
assign F[57][32] = 9'b100000000;
assign F[57][33] = 9'b100000000;
assign F[57][34] = 9'b100100100;
assign F[57][35] = 9'b100100100;
assign F[57][36] = 9'b100000000;
assign F[57][37] = 9'b100000000;
assign F[57][38] = 9'b100000000;
assign F[57][39] = 9'b100000000;
assign F[57][40] = 9'b100000000;
assign F[57][41] = 9'b100000000;
assign F[57][42] = 9'b100000000;
assign F[57][43] = 9'b100000000;
assign F[57][44] = 9'b100100100;
assign F[57][45] = 9'b101000100;
assign F[57][46] = 9'b101101000;
assign F[57][47] = 9'b110001101;
assign F[57][48] = 9'b111110001;
assign F[57][49] = 9'b110101101;
assign F[57][50] = 9'b110101101;
assign F[57][51] = 9'b110101101;
assign F[57][52] = 9'b110101101;
assign F[57][53] = 9'b110101101;
assign F[57][54] = 9'b110101101;
assign F[57][55] = 9'b110101101;
assign F[57][56] = 9'b110101101;
assign F[57][57] = 9'b110101101;
assign F[57][58] = 9'b110101101;
assign F[57][59] = 9'b110101101;
assign F[57][60] = 9'b110101101;
assign F[57][61] = 9'b110110001;
assign F[57][62] = 9'b101101001;
assign F[57][63] = 9'b100000000;
assign F[57][64] = 9'b100000000;
assign F[57][65] = 9'b100000000;
assign F[58][31] = 9'b100000000;
assign F[58][32] = 9'b100100100;
assign F[58][33] = 9'b100100100;
assign F[58][34] = 9'b100100100;
assign F[58][35] = 9'b100100100;
assign F[58][36] = 9'b100000000;
assign F[58][37] = 9'b100000000;
assign F[58][38] = 9'b100000000;
assign F[58][39] = 9'b100000000;
assign F[58][40] = 9'b100000000;
assign F[58][41] = 9'b100000000;
assign F[58][42] = 9'b100000000;
assign F[58][43] = 9'b100000000;
assign F[58][44] = 9'b100000000;
assign F[58][45] = 9'b100000000;
assign F[58][46] = 9'b100100000;
assign F[58][47] = 9'b101000100;
assign F[58][48] = 9'b101101000;
assign F[58][49] = 9'b101101000;
assign F[58][50] = 9'b110001101;
assign F[58][51] = 9'b110101101;
assign F[58][52] = 9'b110101101;
assign F[58][53] = 9'b110101101;
assign F[58][54] = 9'b110101101;
assign F[58][55] = 9'b110101101;
assign F[58][56] = 9'b110101101;
assign F[58][57] = 9'b110101101;
assign F[58][58] = 9'b110101101;
assign F[58][59] = 9'b110101101;
assign F[58][60] = 9'b110101101;
assign F[58][61] = 9'b110001101;
assign F[58][62] = 9'b101001000;
assign F[58][63] = 9'b100000000;
assign F[58][64] = 9'b100000000;
assign F[58][65] = 9'b100000000;
assign F[58][66] = 9'b100000000;
assign F[59][29] = 9'b100000000;
assign F[59][30] = 9'b100000000;
assign F[59][31] = 9'b100000000;
assign F[59][32] = 9'b100100100;
assign F[59][33] = 9'b100100100;
assign F[59][34] = 9'b100100100;
assign F[59][35] = 9'b100100100;
assign F[59][36] = 9'b100000000;
assign F[59][37] = 9'b100000000;
assign F[59][38] = 9'b100000000;
assign F[59][39] = 9'b100000000;
assign F[59][40] = 9'b100000000;
assign F[59][41] = 9'b100000100;
assign F[59][42] = 9'b100100100;
assign F[59][43] = 9'b100100100;
assign F[59][44] = 9'b100000000;
assign F[59][45] = 9'b100000000;
assign F[59][46] = 9'b100000000;
assign F[59][47] = 9'b100000000;
assign F[59][48] = 9'b100100000;
assign F[59][49] = 9'b100100100;
assign F[59][50] = 9'b101000100;
assign F[59][51] = 9'b101101000;
assign F[59][52] = 9'b110001001;
assign F[59][53] = 9'b110001101;
assign F[59][54] = 9'b110101101;
assign F[59][55] = 9'b110101101;
assign F[59][56] = 9'b110101101;
assign F[59][57] = 9'b110101101;
assign F[59][58] = 9'b110101101;
assign F[59][59] = 9'b110101101;
assign F[59][60] = 9'b110101101;
assign F[59][61] = 9'b110001000;
assign F[59][62] = 9'b101000100;
assign F[59][63] = 9'b100000000;
assign F[59][64] = 9'b100000000;
assign F[59][65] = 9'b100000000;
assign F[59][66] = 9'b100000000;
assign F[59][67] = 9'b100000000;
assign F[59][68] = 9'b100000000;
assign F[60][28] = 9'b100000000;
assign F[60][29] = 9'b100000000;
assign F[60][30] = 9'b100000000;
assign F[60][31] = 9'b100100100;
assign F[60][32] = 9'b100000000;
assign F[60][33] = 9'b100000000;
assign F[60][34] = 9'b100000000;
assign F[60][35] = 9'b100000000;
assign F[60][36] = 9'b100000000;
assign F[60][37] = 9'b100000000;
assign F[60][38] = 9'b100000000;
assign F[60][39] = 9'b100000000;
assign F[60][40] = 9'b100000000;
assign F[60][41] = 9'b100000000;
assign F[60][42] = 9'b100000000;
assign F[60][43] = 9'b100000000;
assign F[60][44] = 9'b100000000;
assign F[60][45] = 9'b100000000;
assign F[60][46] = 9'b100000000;
assign F[60][47] = 9'b100000000;
assign F[60][48] = 9'b100000000;
assign F[60][49] = 9'b100000000;
assign F[60][50] = 9'b100000000;
assign F[60][51] = 9'b100100000;
assign F[60][52] = 9'b101000100;
assign F[60][53] = 9'b101101000;
assign F[60][54] = 9'b110001101;
assign F[60][55] = 9'b110001101;
assign F[60][56] = 9'b110001101;
assign F[60][57] = 9'b110001101;
assign F[60][58] = 9'b110001101;
assign F[60][59] = 9'b110001101;
assign F[60][60] = 9'b110001101;
assign F[60][61] = 9'b110001000;
assign F[60][62] = 9'b101000100;
assign F[60][63] = 9'b100000000;
assign F[60][64] = 9'b100000000;
assign F[60][65] = 9'b100000000;
assign F[60][66] = 9'b100000000;
assign F[60][67] = 9'b100000000;
assign F[60][68] = 9'b100000000;
assign F[60][69] = 9'b100000000;
assign F[61][27] = 9'b100000000;
assign F[61][28] = 9'b100000000;
assign F[61][29] = 9'b100100100;
assign F[61][30] = 9'b100100100;
assign F[61][31] = 9'b100000000;
assign F[61][32] = 9'b100000000;
assign F[61][33] = 9'b100000000;
assign F[61][34] = 9'b100000000;
assign F[61][35] = 9'b100000000;
assign F[61][36] = 9'b100000000;
assign F[61][37] = 9'b100000000;
assign F[61][38] = 9'b100000000;
assign F[61][39] = 9'b100000000;
assign F[61][40] = 9'b100000000;
assign F[61][41] = 9'b100000000;
assign F[61][42] = 9'b100000000;
assign F[61][43] = 9'b100000000;
assign F[61][44] = 9'b100000000;
assign F[61][45] = 9'b100000000;
assign F[61][46] = 9'b100000000;
assign F[61][47] = 9'b100000000;
assign F[61][48] = 9'b100000000;
assign F[61][49] = 9'b100000000;
assign F[61][50] = 9'b100000000;
assign F[61][51] = 9'b100000000;
assign F[61][52] = 9'b100000000;
assign F[61][53] = 9'b100100100;
assign F[61][54] = 9'b101001000;
assign F[61][55] = 9'b101000100;
assign F[61][56] = 9'b101101000;
assign F[61][57] = 9'b101101000;
assign F[61][58] = 9'b101101000;
assign F[61][59] = 9'b101101000;
assign F[61][60] = 9'b101101000;
assign F[61][61] = 9'b101101000;
assign F[61][62] = 9'b101000100;
assign F[61][63] = 9'b100000000;
assign F[61][64] = 9'b100000000;
assign F[61][65] = 9'b100000000;
assign F[61][66] = 9'b100100100;
assign F[61][67] = 9'b100100100;
assign F[61][68] = 9'b100000000;
assign F[61][69] = 9'b100000000;
assign F[61][70] = 9'b100000000;
assign F[62][26] = 9'b100000000;
assign F[62][27] = 9'b100100100;
assign F[62][28] = 9'b101101101;
assign F[62][29] = 9'b101001001;
assign F[62][30] = 9'b101001000;
assign F[62][31] = 9'b100000000;
assign F[62][32] = 9'b100000000;
assign F[62][33] = 9'b100000000;
assign F[62][34] = 9'b100000000;
assign F[62][35] = 9'b100000000;
assign F[62][36] = 9'b100000000;
assign F[62][37] = 9'b100000000;
assign F[62][38] = 9'b100000000;
assign F[62][39] = 9'b100000000;
assign F[62][40] = 9'b100000000;
assign F[62][41] = 9'b100000000;
assign F[62][42] = 9'b100000000;
assign F[62][43] = 9'b100000000;
assign F[62][44] = 9'b100000000;
assign F[62][45] = 9'b100000000;
assign F[62][46] = 9'b100000000;
assign F[62][47] = 9'b100000000;
assign F[62][48] = 9'b100000000;
assign F[62][49] = 9'b100000000;
assign F[62][50] = 9'b100000000;
assign F[62][51] = 9'b100000000;
assign F[62][52] = 9'b100000000;
assign F[62][53] = 9'b100000000;
assign F[62][54] = 9'b100000000;
assign F[62][55] = 9'b100000000;
assign F[62][56] = 9'b100100100;
assign F[62][57] = 9'b101101000;
assign F[62][58] = 9'b101101000;
assign F[62][59] = 9'b101101000;
assign F[62][60] = 9'b101101000;
assign F[62][61] = 9'b101101000;
assign F[62][62] = 9'b101000100;
assign F[62][63] = 9'b100000000;
assign F[62][64] = 9'b100000000;
assign F[62][65] = 9'b100000000;
assign F[62][66] = 9'b100000000;
assign F[62][67] = 9'b100000000;
assign F[62][68] = 9'b100000000;
assign F[62][69] = 9'b100100100;
assign F[62][70] = 9'b100000000;
assign F[62][71] = 9'b100000000;
assign F[63][24] = 9'b100000000;
assign F[63][25] = 9'b100000000;
assign F[63][26] = 9'b100000000;
assign F[63][27] = 9'b100100100;
assign F[63][28] = 9'b101101101;
assign F[63][29] = 9'b101001001;
assign F[63][30] = 9'b100100100;
assign F[63][31] = 9'b100000000;
assign F[63][32] = 9'b100000000;
assign F[63][33] = 9'b100000000;
assign F[63][34] = 9'b100000000;
assign F[63][35] = 9'b100000000;
assign F[63][36] = 9'b100000000;
assign F[63][37] = 9'b100000000;
assign F[63][38] = 9'b100000000;
assign F[63][39] = 9'b100000000;
assign F[63][40] = 9'b100000000;
assign F[63][41] = 9'b100000000;
assign F[63][42] = 9'b100000000;
assign F[63][43] = 9'b100000000;
assign F[63][44] = 9'b100000000;
assign F[63][45] = 9'b100000000;
assign F[63][46] = 9'b100000000;
assign F[63][47] = 9'b100000000;
assign F[63][48] = 9'b100000000;
assign F[63][49] = 9'b100000000;
assign F[63][50] = 9'b100000000;
assign F[63][51] = 9'b100000000;
assign F[63][52] = 9'b100000000;
assign F[63][53] = 9'b100000000;
assign F[63][54] = 9'b100000000;
assign F[63][55] = 9'b100000000;
assign F[63][56] = 9'b100000000;
assign F[63][57] = 9'b100000000;
assign F[63][58] = 9'b101001000;
assign F[63][59] = 9'b110001101;
assign F[63][60] = 9'b110101101;
assign F[63][61] = 9'b110001000;
assign F[63][62] = 9'b101000100;
assign F[63][63] = 9'b100000000;
assign F[63][64] = 9'b100000000;
assign F[63][65] = 9'b100000000;
assign F[63][66] = 9'b100000000;
assign F[63][67] = 9'b100000000;
assign F[63][68] = 9'b100000000;
assign F[63][69] = 9'b100000000;
assign F[63][70] = 9'b100000000;
assign F[63][71] = 9'b100000000;
assign F[63][72] = 9'b100000000;
assign F[63][73] = 9'b100000000;
assign F[64][23] = 9'b100000000;
assign F[64][24] = 9'b100000000;
assign F[64][25] = 9'b100000000;
assign F[64][26] = 9'b101001001;
assign F[64][27] = 9'b101001001;
assign F[64][28] = 9'b101001001;
assign F[64][29] = 9'b100100100;
assign F[64][30] = 9'b100000000;
assign F[64][31] = 9'b100000000;
assign F[64][32] = 9'b100000000;
assign F[64][33] = 9'b100000000;
assign F[64][34] = 9'b100000000;
assign F[64][35] = 9'b100000000;
assign F[64][36] = 9'b100000000;
assign F[64][37] = 9'b100000000;
assign F[64][38] = 9'b100000000;
assign F[64][39] = 9'b100000000;
assign F[64][40] = 9'b100000000;
assign F[64][41] = 9'b100000000;
assign F[64][42] = 9'b100000000;
assign F[64][43] = 9'b100000000;
assign F[64][44] = 9'b100000000;
assign F[64][45] = 9'b100000000;
assign F[64][46] = 9'b100000000;
assign F[64][47] = 9'b100000000;
assign F[64][48] = 9'b100000000;
assign F[64][49] = 9'b100000000;
assign F[64][50] = 9'b100000000;
assign F[64][51] = 9'b100000000;
assign F[64][52] = 9'b100000000;
assign F[64][53] = 9'b100000000;
assign F[64][54] = 9'b100000000;
assign F[64][55] = 9'b100000000;
assign F[64][56] = 9'b100000000;
assign F[64][57] = 9'b100000000;
assign F[64][58] = 9'b100000000;
assign F[64][59] = 9'b101000100;
assign F[64][60] = 9'b111110001;
assign F[64][61] = 9'b110001000;
assign F[64][62] = 9'b101000100;
assign F[64][63] = 9'b100100000;
assign F[64][64] = 9'b100000000;
assign F[64][65] = 9'b100000000;
assign F[64][66] = 9'b100000000;
assign F[64][67] = 9'b100000000;
assign F[64][68] = 9'b100000000;
assign F[64][69] = 9'b100000000;
assign F[64][70] = 9'b100000000;
assign F[64][71] = 9'b100000000;
assign F[64][72] = 9'b100000000;
assign F[64][73] = 9'b100000000;
assign F[64][74] = 9'b100000000;
assign F[65][21] = 9'b100000000;
assign F[65][22] = 9'b100000000;
assign F[65][23] = 9'b101001000;
assign F[65][24] = 9'b101001001;
assign F[65][25] = 9'b101001000;
assign F[65][26] = 9'b100100100;
assign F[65][27] = 9'b100100100;
assign F[65][28] = 9'b100100100;
assign F[65][29] = 9'b100000000;
assign F[65][30] = 9'b100000000;
assign F[65][31] = 9'b100000000;
assign F[65][32] = 9'b100000000;
assign F[65][33] = 9'b100000000;
assign F[65][34] = 9'b100000000;
assign F[65][35] = 9'b100000000;
assign F[65][36] = 9'b100000000;
assign F[65][37] = 9'b100000000;
assign F[65][38] = 9'b100000000;
assign F[65][39] = 9'b100000000;
assign F[65][40] = 9'b100000000;
assign F[65][41] = 9'b100000000;
assign F[65][42] = 9'b100000000;
assign F[65][43] = 9'b100000000;
assign F[65][44] = 9'b100000000;
assign F[65][45] = 9'b100000000;
assign F[65][46] = 9'b100000000;
assign F[65][47] = 9'b100000000;
assign F[65][48] = 9'b100000000;
assign F[65][49] = 9'b100000000;
assign F[65][50] = 9'b100000000;
assign F[65][51] = 9'b100000000;
assign F[65][52] = 9'b100000000;
assign F[65][53] = 9'b100000000;
assign F[65][54] = 9'b100000000;
assign F[65][55] = 9'b100000000;
assign F[65][56] = 9'b100000000;
assign F[65][57] = 9'b100000000;
assign F[65][58] = 9'b100000000;
assign F[65][59] = 9'b100100100;
assign F[65][60] = 9'b110001101;
assign F[65][61] = 9'b101101000;
assign F[65][62] = 9'b101001000;
assign F[65][63] = 9'b100100000;
assign F[65][64] = 9'b100000000;
assign F[65][65] = 9'b100000000;
assign F[65][66] = 9'b100000000;
assign F[65][67] = 9'b100000000;
assign F[65][68] = 9'b100000000;
assign F[65][69] = 9'b100000000;
assign F[65][70] = 9'b100000000;
assign F[65][71] = 9'b100000000;
assign F[65][72] = 9'b100000000;
assign F[65][73] = 9'b100000000;
assign F[65][74] = 9'b100000000;
assign F[65][75] = 9'b100000000;
assign F[65][76] = 9'b100000000;
assign F[65][77] = 9'b100000000;
assign F[66][20] = 9'b100000000;
assign F[66][21] = 9'b100100100;
assign F[66][22] = 9'b101001001;
assign F[66][23] = 9'b101101101;
assign F[66][24] = 9'b101001001;
assign F[66][25] = 9'b100100100;
assign F[66][26] = 9'b100000000;
assign F[66][27] = 9'b100000000;
assign F[66][28] = 9'b100000000;
assign F[66][29] = 9'b100000000;
assign F[66][30] = 9'b100000000;
assign F[66][31] = 9'b100000000;
assign F[66][32] = 9'b100000000;
assign F[66][33] = 9'b100000000;
assign F[66][34] = 9'b100000000;
assign F[66][35] = 9'b100000000;
assign F[66][36] = 9'b100000000;
assign F[66][37] = 9'b100000000;
assign F[66][38] = 9'b100000000;
assign F[66][39] = 9'b100000000;
assign F[66][40] = 9'b100000000;
assign F[66][41] = 9'b100000000;
assign F[66][42] = 9'b100000000;
assign F[66][43] = 9'b100000000;
assign F[66][44] = 9'b100000000;
assign F[66][45] = 9'b100000000;
assign F[66][46] = 9'b100000000;
assign F[66][47] = 9'b100000000;
assign F[66][48] = 9'b100000000;
assign F[66][49] = 9'b100000000;
assign F[66][50] = 9'b100000000;
assign F[66][51] = 9'b100000000;
assign F[66][52] = 9'b100000000;
assign F[66][53] = 9'b100000000;
assign F[66][54] = 9'b100000000;
assign F[66][55] = 9'b100000000;
assign F[66][56] = 9'b100000000;
assign F[66][57] = 9'b100000000;
assign F[66][58] = 9'b100000000;
assign F[66][59] = 9'b100100100;
assign F[66][60] = 9'b101101000;
assign F[66][61] = 9'b101101000;
assign F[66][62] = 9'b101101000;
assign F[66][63] = 9'b100100000;
assign F[66][64] = 9'b100000000;
assign F[66][65] = 9'b100000000;
assign F[66][66] = 9'b100000000;
assign F[66][67] = 9'b100000000;
assign F[66][68] = 9'b100000000;
assign F[66][69] = 9'b100000000;
assign F[66][70] = 9'b100000000;
assign F[66][71] = 9'b100000000;
assign F[66][72] = 9'b100000000;
assign F[66][73] = 9'b100000000;
assign F[66][74] = 9'b100000000;
assign F[66][75] = 9'b100000000;
assign F[66][76] = 9'b100000000;
assign F[66][77] = 9'b100000000;
assign F[66][78] = 9'b100000000;
assign F[67][19] = 9'b100000000;
assign F[67][20] = 9'b100000000;
assign F[67][21] = 9'b101001001;
assign F[67][22] = 9'b101101101;
assign F[67][23] = 9'b101001000;
assign F[67][24] = 9'b100100100;
assign F[67][25] = 9'b100000000;
assign F[67][26] = 9'b100000000;
assign F[67][27] = 9'b100000000;
assign F[67][28] = 9'b100000000;
assign F[67][29] = 9'b100000000;
assign F[67][30] = 9'b100000000;
assign F[67][31] = 9'b100000000;
assign F[67][32] = 9'b100000000;
assign F[67][33] = 9'b100000000;
assign F[67][34] = 9'b100000000;
assign F[67][35] = 9'b100000000;
assign F[67][36] = 9'b100000000;
assign F[67][37] = 9'b100000000;
assign F[67][38] = 9'b100000000;
assign F[67][39] = 9'b100000000;
assign F[67][40] = 9'b100000000;
assign F[67][41] = 9'b100000000;
assign F[67][42] = 9'b100000000;
assign F[67][43] = 9'b100000000;
assign F[67][44] = 9'b100000000;
assign F[67][45] = 9'b100000000;
assign F[67][46] = 9'b100000000;
assign F[67][47] = 9'b100000000;
assign F[67][48] = 9'b100000000;
assign F[67][49] = 9'b100000000;
assign F[67][50] = 9'b100000000;
assign F[67][51] = 9'b100000000;
assign F[67][52] = 9'b100000000;
assign F[67][53] = 9'b100000000;
assign F[67][54] = 9'b100000000;
assign F[67][55] = 9'b100000000;
assign F[67][56] = 9'b100000000;
assign F[67][57] = 9'b100000000;
assign F[67][58] = 9'b100000000;
assign F[67][59] = 9'b100000000;
assign F[67][60] = 9'b100100100;
assign F[67][61] = 9'b101101000;
assign F[67][62] = 9'b101101000;
assign F[67][63] = 9'b100100000;
assign F[67][64] = 9'b100000000;
assign F[67][65] = 9'b100000000;
assign F[67][66] = 9'b100000000;
assign F[67][67] = 9'b100000000;
assign F[67][68] = 9'b100000000;
assign F[67][69] = 9'b100000000;
assign F[67][70] = 9'b100000000;
assign F[67][71] = 9'b100000000;
assign F[67][72] = 9'b100000000;
assign F[67][73] = 9'b100000000;
assign F[67][74] = 9'b100000000;
assign F[67][75] = 9'b100000000;
assign F[67][76] = 9'b100000000;
assign F[67][77] = 9'b100000000;
assign F[67][78] = 9'b100000000;
assign F[67][79] = 9'b100000000;
assign F[67][80] = 9'b100000000;
assign F[68][18] = 9'b100000000;
assign F[68][19] = 9'b100000000;
assign F[68][20] = 9'b101001000;
assign F[68][21] = 9'b101001000;
assign F[68][22] = 9'b100100100;
assign F[68][23] = 9'b100000000;
assign F[68][24] = 9'b100000000;
assign F[68][25] = 9'b100000000;
assign F[68][26] = 9'b100000000;
assign F[68][27] = 9'b100000000;
assign F[68][28] = 9'b100000000;
assign F[68][29] = 9'b100000000;
assign F[68][30] = 9'b100000000;
assign F[68][31] = 9'b100000000;
assign F[68][32] = 9'b100000000;
assign F[68][33] = 9'b100000000;
assign F[68][34] = 9'b100000000;
assign F[68][35] = 9'b100000000;
assign F[68][36] = 9'b100000000;
assign F[68][37] = 9'b100000000;
assign F[68][38] = 9'b100000000;
assign F[68][39] = 9'b100000000;
assign F[68][40] = 9'b100000000;
assign F[68][41] = 9'b100000000;
assign F[68][42] = 9'b100000000;
assign F[68][43] = 9'b100000000;
assign F[68][44] = 9'b100000000;
assign F[68][45] = 9'b100000000;
assign F[68][46] = 9'b100000000;
assign F[68][47] = 9'b100000000;
assign F[68][48] = 9'b100000000;
assign F[68][49] = 9'b100000000;
assign F[68][50] = 9'b100000000;
assign F[68][51] = 9'b100000000;
assign F[68][52] = 9'b100000000;
assign F[68][53] = 9'b100000000;
assign F[68][54] = 9'b100000000;
assign F[68][55] = 9'b100000000;
assign F[68][56] = 9'b100000000;
assign F[68][57] = 9'b100000000;
assign F[68][58] = 9'b100000000;
assign F[68][59] = 9'b100000000;
assign F[68][60] = 9'b100000000;
assign F[68][61] = 9'b101001000;
assign F[68][62] = 9'b101001000;
assign F[68][63] = 9'b100100000;
assign F[68][64] = 9'b100000000;
assign F[68][65] = 9'b100000000;
assign F[68][66] = 9'b100000000;
assign F[68][67] = 9'b100000000;
assign F[68][68] = 9'b100000000;
assign F[68][69] = 9'b100000000;
assign F[68][70] = 9'b100000000;
assign F[68][71] = 9'b100000000;
assign F[68][72] = 9'b100000000;
assign F[68][73] = 9'b100000000;
assign F[68][74] = 9'b100000000;
assign F[68][75] = 9'b100000000;
assign F[68][76] = 9'b100000000;
assign F[68][77] = 9'b100000000;
assign F[68][78] = 9'b100000000;
assign F[68][79] = 9'b100000000;
assign F[68][80] = 9'b100000000;
assign F[69][17] = 9'b100000000;
assign F[69][18] = 9'b100100100;
assign F[69][19] = 9'b101001001;
assign F[69][20] = 9'b100100100;
assign F[69][21] = 9'b100100100;
assign F[69][22] = 9'b100000000;
assign F[69][23] = 9'b100000000;
assign F[69][24] = 9'b100000000;
assign F[69][25] = 9'b100000000;
assign F[69][26] = 9'b100000000;
assign F[69][27] = 9'b100000000;
assign F[69][28] = 9'b100000000;
assign F[69][29] = 9'b100000000;
assign F[69][30] = 9'b100000000;
assign F[69][31] = 9'b100000000;
assign F[69][32] = 9'b100000000;
assign F[69][33] = 9'b100000000;
assign F[69][34] = 9'b100000000;
assign F[69][35] = 9'b100000000;
assign F[69][36] = 9'b100000000;
assign F[69][37] = 9'b100000000;
assign F[69][38] = 9'b100000000;
assign F[69][39] = 9'b100000000;
assign F[69][40] = 9'b100000000;
assign F[69][41] = 9'b100000000;
assign F[69][42] = 9'b100000000;
assign F[69][43] = 9'b100000000;
assign F[69][44] = 9'b100000000;
assign F[69][45] = 9'b100000000;
assign F[69][46] = 9'b100000000;
assign F[69][47] = 9'b100000000;
assign F[69][48] = 9'b100000000;
assign F[69][49] = 9'b100000000;
assign F[69][50] = 9'b100000000;
assign F[69][51] = 9'b100000000;
assign F[69][52] = 9'b100000000;
assign F[69][53] = 9'b100000000;
assign F[69][54] = 9'b100000000;
assign F[69][55] = 9'b100000000;
assign F[69][56] = 9'b100000000;
assign F[69][57] = 9'b100000000;
assign F[69][58] = 9'b100000000;
assign F[69][59] = 9'b100000000;
assign F[69][60] = 9'b100000000;
assign F[69][61] = 9'b100100100;
assign F[69][62] = 9'b101000100;
assign F[69][63] = 9'b100100100;
assign F[69][64] = 9'b100000000;
assign F[69][65] = 9'b100000000;
assign F[69][66] = 9'b100000000;
assign F[69][67] = 9'b100000000;
assign F[69][68] = 9'b100000000;
assign F[69][69] = 9'b100000000;
assign F[69][70] = 9'b100000000;
assign F[69][71] = 9'b100000000;
assign F[69][72] = 9'b100000000;
assign F[69][73] = 9'b100000000;
assign F[69][74] = 9'b100000000;
assign F[69][75] = 9'b100000000;
assign F[69][76] = 9'b100000000;
assign F[69][77] = 9'b100000000;
assign F[69][78] = 9'b100000000;
assign F[69][79] = 9'b100000000;
assign F[69][80] = 9'b100000000;
assign F[70][14] = 9'b100000000;
assign F[70][15] = 9'b100000000;
assign F[70][16] = 9'b100000000;
assign F[70][17] = 9'b100100100;
assign F[70][18] = 9'b100100100;
assign F[70][19] = 9'b100100100;
assign F[70][20] = 9'b100100100;
assign F[70][21] = 9'b100000000;
assign F[70][22] = 9'b100000000;
assign F[70][23] = 9'b100000000;
assign F[70][24] = 9'b100000000;
assign F[70][25] = 9'b100000000;
assign F[70][26] = 9'b100000000;
assign F[70][27] = 9'b100000000;
assign F[70][28] = 9'b100000000;
assign F[70][29] = 9'b100000000;
assign F[70][30] = 9'b100000000;
assign F[70][31] = 9'b100000000;
assign F[70][32] = 9'b100000000;
assign F[70][33] = 9'b100000000;
assign F[70][34] = 9'b100000000;
assign F[70][35] = 9'b100000000;
assign F[70][36] = 9'b100000000;
assign F[70][37] = 9'b100000000;
assign F[70][38] = 9'b100000000;
assign F[70][39] = 9'b100000000;
assign F[70][40] = 9'b100000000;
assign F[70][41] = 9'b100000000;
assign F[70][42] = 9'b100000000;
assign F[70][43] = 9'b100000000;
assign F[70][44] = 9'b100000000;
assign F[70][45] = 9'b100000000;
assign F[70][46] = 9'b100000000;
assign F[70][47] = 9'b100000000;
assign F[70][48] = 9'b100000000;
assign F[70][49] = 9'b100000000;
assign F[70][50] = 9'b100000000;
assign F[70][51] = 9'b100000000;
assign F[70][52] = 9'b100000000;
assign F[70][53] = 9'b100000000;
assign F[70][54] = 9'b100000000;
assign F[70][55] = 9'b100000000;
assign F[70][56] = 9'b100000000;
assign F[70][57] = 9'b100000000;
assign F[70][58] = 9'b100000000;
assign F[70][59] = 9'b100000000;
assign F[70][60] = 9'b100000000;
assign F[70][61] = 9'b100000000;
assign F[70][62] = 9'b100100100;
assign F[70][63] = 9'b101001000;
assign F[70][64] = 9'b100000000;
assign F[70][65] = 9'b100000000;
assign F[70][66] = 9'b100000000;
assign F[70][67] = 9'b100000000;
assign F[70][68] = 9'b100000000;
assign F[70][69] = 9'b100000000;
assign F[70][70] = 9'b100000000;
assign F[70][71] = 9'b100000000;
assign F[70][72] = 9'b100000000;
assign F[70][73] = 9'b100000000;
assign F[70][74] = 9'b100000000;
assign F[70][75] = 9'b100000000;
assign F[70][76] = 9'b100000000;
assign F[70][77] = 9'b100000000;
assign F[70][78] = 9'b100000000;
assign F[70][79] = 9'b100000000;
assign F[70][80] = 9'b100000000;
assign F[70][81] = 9'b100000000;
assign F[70][82] = 9'b100000000;
assign F[71][12] = 9'b100000000;
assign F[71][13] = 9'b100000000;
assign F[71][14] = 9'b100000000;
assign F[71][15] = 9'b100000000;
assign F[71][16] = 9'b100100100;
assign F[71][17] = 9'b100100100;
assign F[71][18] = 9'b100100100;
assign F[71][19] = 9'b100100100;
assign F[71][20] = 9'b100100100;
assign F[71][21] = 9'b100000000;
assign F[71][22] = 9'b100000000;
assign F[71][23] = 9'b100000000;
assign F[71][24] = 9'b100000000;
assign F[71][25] = 9'b100000000;
assign F[71][26] = 9'b100000000;
assign F[71][27] = 9'b100000000;
assign F[71][28] = 9'b100000000;
assign F[71][29] = 9'b100000000;
assign F[71][30] = 9'b100000000;
assign F[71][31] = 9'b100000000;
assign F[71][32] = 9'b100000000;
assign F[71][33] = 9'b100000000;
assign F[71][34] = 9'b100000000;
assign F[71][35] = 9'b100000000;
assign F[71][36] = 9'b100000000;
assign F[71][37] = 9'b100000000;
assign F[71][38] = 9'b100000000;
assign F[71][39] = 9'b100000000;
assign F[71][40] = 9'b100000000;
assign F[71][41] = 9'b100000000;
assign F[71][42] = 9'b100000000;
assign F[71][43] = 9'b100000000;
assign F[71][44] = 9'b100000000;
assign F[71][45] = 9'b100000000;
assign F[71][46] = 9'b100000000;
assign F[71][47] = 9'b100000000;
assign F[71][48] = 9'b100000000;
assign F[71][49] = 9'b100000000;
assign F[71][50] = 9'b100000000;
assign F[71][51] = 9'b100000000;
assign F[71][52] = 9'b100000000;
assign F[71][53] = 9'b100000000;
assign F[71][54] = 9'b100000000;
assign F[71][55] = 9'b100000000;
assign F[71][56] = 9'b100000000;
assign F[71][57] = 9'b100000000;
assign F[71][58] = 9'b100000000;
assign F[71][59] = 9'b100000000;
assign F[71][60] = 9'b100000000;
assign F[71][61] = 9'b100000000;
assign F[71][62] = 9'b100000000;
assign F[71][63] = 9'b100000000;
assign F[71][64] = 9'b100000000;
assign F[71][65] = 9'b100000000;
assign F[71][66] = 9'b100000000;
assign F[71][67] = 9'b100000000;
assign F[71][68] = 9'b100000000;
assign F[71][69] = 9'b100000000;
assign F[71][70] = 9'b100000000;
assign F[71][71] = 9'b100000000;
assign F[71][72] = 9'b100000000;
assign F[71][73] = 9'b100100100;
assign F[71][74] = 9'b101001000;
assign F[71][75] = 9'b101101101;
assign F[71][76] = 9'b101101101;
assign F[71][77] = 9'b101101101;
assign F[71][78] = 9'b101101101;
assign F[71][79] = 9'b100100100;
assign F[71][80] = 9'b100000000;
assign F[71][81] = 9'b100000000;
assign F[71][82] = 9'b100000000;
assign F[72][12] = 9'b100000000;
assign F[72][13] = 9'b100000000;
assign F[72][14] = 9'b100100100;
assign F[72][15] = 9'b100100100;
assign F[72][16] = 9'b100100100;
assign F[72][17] = 9'b100100100;
assign F[72][18] = 9'b100100100;
assign F[72][19] = 9'b100100100;
assign F[72][20] = 9'b100100100;
assign F[72][21] = 9'b100100100;
assign F[72][22] = 9'b100000000;
assign F[72][23] = 9'b100000000;
assign F[72][24] = 9'b100000000;
assign F[72][25] = 9'b100000000;
assign F[72][26] = 9'b100000000;
assign F[72][27] = 9'b100000000;
assign F[72][28] = 9'b100000000;
assign F[72][29] = 9'b100000000;
assign F[72][30] = 9'b100000000;
assign F[72][31] = 9'b100000000;
assign F[72][32] = 9'b100000000;
assign F[72][33] = 9'b100000000;
assign F[72][34] = 9'b100000000;
assign F[72][35] = 9'b100000000;
assign F[72][36] = 9'b100000000;
assign F[72][37] = 9'b100000000;
assign F[72][38] = 9'b100000000;
assign F[72][39] = 9'b100000000;
assign F[72][40] = 9'b100000000;
assign F[72][41] = 9'b100000000;
assign F[72][42] = 9'b100000000;
assign F[72][43] = 9'b100000000;
assign F[72][44] = 9'b100000000;
assign F[72][45] = 9'b100000000;
assign F[72][46] = 9'b100000000;
assign F[72][47] = 9'b100000000;
assign F[72][48] = 9'b100000000;
assign F[72][49] = 9'b100000000;
assign F[72][50] = 9'b100000000;
assign F[72][51] = 9'b100000000;
assign F[72][52] = 9'b100000000;
assign F[72][53] = 9'b100000000;
assign F[72][54] = 9'b100000000;
assign F[72][55] = 9'b100000000;
assign F[72][56] = 9'b100000000;
assign F[72][57] = 9'b100000000;
assign F[72][58] = 9'b100000000;
assign F[72][59] = 9'b100000000;
assign F[72][60] = 9'b100000000;
assign F[72][61] = 9'b100000000;
assign F[72][62] = 9'b100000000;
assign F[72][63] = 9'b100000000;
assign F[72][64] = 9'b100000000;
assign F[72][65] = 9'b100000000;
assign F[72][66] = 9'b100000000;
assign F[72][67] = 9'b100000000;
assign F[72][68] = 9'b100000000;
assign F[72][69] = 9'b100000000;
assign F[72][70] = 9'b100000000;
assign F[72][71] = 9'b100000000;
assign F[72][72] = 9'b100000000;
assign F[72][73] = 9'b100000000;
assign F[72][74] = 9'b100100100;
assign F[72][75] = 9'b101001001;
assign F[72][76] = 9'b101101101;
assign F[72][77] = 9'b110010010;
assign F[72][78] = 9'b110010001;
assign F[72][79] = 9'b101001001;
assign F[72][80] = 9'b100100100;
assign F[72][81] = 9'b100000000;
assign F[72][82] = 9'b100000000;
assign F[73][11] = 9'b100000000;
assign F[73][12] = 9'b100000000;
assign F[73][13] = 9'b100000000;
assign F[73][14] = 9'b100100100;
assign F[73][15] = 9'b100100100;
assign F[73][16] = 9'b100100100;
assign F[73][17] = 9'b100100100;
assign F[73][18] = 9'b100100100;
assign F[73][19] = 9'b100100100;
assign F[73][20] = 9'b100100100;
assign F[73][21] = 9'b100100100;
assign F[73][22] = 9'b100100100;
assign F[73][23] = 9'b100000000;
assign F[73][24] = 9'b100000000;
assign F[73][25] = 9'b100000000;
assign F[73][26] = 9'b100000000;
assign F[73][27] = 9'b100000000;
assign F[73][28] = 9'b100000000;
assign F[73][29] = 9'b100000000;
assign F[73][30] = 9'b100000000;
assign F[73][31] = 9'b100000000;
assign F[73][32] = 9'b100000000;
assign F[73][33] = 9'b100000000;
assign F[73][34] = 9'b100000000;
assign F[73][35] = 9'b100000000;
assign F[73][36] = 9'b100000000;
assign F[73][37] = 9'b100000000;
assign F[73][38] = 9'b100000000;
assign F[73][39] = 9'b100000000;
assign F[73][40] = 9'b100000000;
assign F[73][41] = 9'b100000000;
assign F[73][42] = 9'b100000000;
assign F[73][43] = 9'b100000000;
assign F[73][44] = 9'b100000000;
assign F[73][45] = 9'b100000000;
assign F[73][46] = 9'b100000000;
assign F[73][47] = 9'b100000000;
assign F[73][48] = 9'b100000000;
assign F[73][49] = 9'b100000000;
assign F[73][50] = 9'b100000000;
assign F[73][51] = 9'b100000000;
assign F[73][52] = 9'b100000000;
assign F[73][53] = 9'b100000000;
assign F[73][54] = 9'b100000000;
assign F[73][55] = 9'b100000000;
assign F[73][56] = 9'b100000000;
assign F[73][57] = 9'b100000000;
assign F[73][58] = 9'b100000000;
assign F[73][59] = 9'b100000000;
assign F[73][60] = 9'b100000000;
assign F[73][61] = 9'b100000000;
assign F[73][62] = 9'b100000000;
assign F[73][63] = 9'b100000000;
assign F[73][64] = 9'b100000000;
assign F[73][65] = 9'b100000000;
assign F[73][66] = 9'b100000000;
assign F[73][67] = 9'b100000000;
assign F[73][68] = 9'b100000000;
assign F[73][69] = 9'b100000000;
assign F[73][70] = 9'b100000000;
assign F[73][71] = 9'b100000000;
assign F[73][72] = 9'b100000000;
assign F[73][73] = 9'b100000000;
assign F[73][74] = 9'b100000000;
assign F[73][75] = 9'b100100100;
assign F[73][76] = 9'b101001000;
assign F[73][77] = 9'b101001001;
assign F[73][78] = 9'b101101101;
assign F[73][79] = 9'b101001001;
assign F[73][80] = 9'b101001000;
assign F[73][81] = 9'b100000000;
assign F[73][82] = 9'b100000000;
assign F[73][83] = 9'b100000000;
assign F[74][10] = 9'b100000000;
assign F[74][11] = 9'b100000000;
assign F[74][12] = 9'b100100100;
assign F[74][13] = 9'b100100100;
assign F[74][14] = 9'b100100100;
assign F[74][15] = 9'b100100100;
assign F[74][16] = 9'b100100100;
assign F[74][17] = 9'b100100100;
assign F[74][18] = 9'b100100100;
assign F[74][19] = 9'b100100100;
assign F[74][20] = 9'b100100100;
assign F[74][21] = 9'b100100100;
assign F[74][22] = 9'b100100100;
assign F[74][23] = 9'b100100100;
assign F[74][24] = 9'b100100100;
assign F[74][25] = 9'b100100100;
assign F[74][26] = 9'b100000000;
assign F[74][27] = 9'b100000000;
assign F[74][28] = 9'b100000000;
assign F[74][29] = 9'b100000000;
assign F[74][30] = 9'b100000000;
assign F[74][31] = 9'b100000000;
assign F[74][32] = 9'b100000000;
assign F[74][33] = 9'b100000000;
assign F[74][34] = 9'b100000000;
assign F[74][35] = 9'b100000000;
assign F[74][36] = 9'b100000000;
assign F[74][37] = 9'b100000000;
assign F[74][38] = 9'b100000000;
assign F[74][39] = 9'b100000000;
assign F[74][40] = 9'b100000000;
assign F[74][41] = 9'b100000000;
assign F[74][42] = 9'b100000000;
assign F[74][43] = 9'b100000000;
assign F[74][44] = 9'b100000000;
assign F[74][45] = 9'b100000000;
assign F[74][46] = 9'b100000000;
assign F[74][47] = 9'b100000000;
assign F[74][48] = 9'b100000000;
assign F[74][49] = 9'b100000000;
assign F[74][50] = 9'b100000000;
assign F[74][51] = 9'b100000000;
assign F[74][52] = 9'b100000000;
assign F[74][53] = 9'b100000000;
assign F[74][54] = 9'b100000000;
assign F[74][55] = 9'b100000000;
assign F[74][56] = 9'b100000000;
assign F[74][57] = 9'b100000000;
assign F[74][58] = 9'b100000000;
assign F[74][59] = 9'b100000000;
assign F[74][60] = 9'b100000000;
assign F[74][61] = 9'b100000000;
assign F[74][62] = 9'b100000000;
assign F[74][63] = 9'b100000000;
assign F[74][64] = 9'b100000000;
assign F[74][65] = 9'b100000000;
assign F[74][66] = 9'b100100100;
assign F[74][67] = 9'b100000000;
assign F[74][68] = 9'b100000000;
assign F[74][69] = 9'b100000000;
assign F[74][70] = 9'b100000000;
assign F[74][71] = 9'b100000000;
assign F[74][72] = 9'b100000000;
assign F[74][73] = 9'b100000000;
assign F[74][74] = 9'b100000000;
assign F[74][75] = 9'b100000000;
assign F[74][76] = 9'b100000000;
assign F[74][77] = 9'b100000000;
assign F[74][78] = 9'b100100100;
assign F[74][79] = 9'b100100100;
assign F[74][80] = 9'b100100100;
assign F[74][81] = 9'b100100100;
assign F[74][82] = 9'b100000000;
assign F[74][83] = 9'b100000000;
assign F[75][9] = 9'b100000000;
assign F[75][10] = 9'b100000000;
assign F[75][11] = 9'b100100100;
assign F[75][12] = 9'b100100100;
assign F[75][13] = 9'b100100100;
assign F[75][14] = 9'b100100100;
assign F[75][15] = 9'b100100100;
assign F[75][16] = 9'b100100100;
assign F[75][17] = 9'b100100100;
assign F[75][18] = 9'b100100100;
assign F[75][19] = 9'b100100100;
assign F[75][20] = 9'b100100100;
assign F[75][21] = 9'b100100100;
assign F[75][22] = 9'b100100100;
assign F[75][23] = 9'b100000000;
assign F[75][24] = 9'b100100100;
assign F[75][25] = 9'b100100100;
assign F[75][26] = 9'b100100100;
assign F[75][27] = 9'b100000000;
assign F[75][28] = 9'b100000000;
assign F[75][29] = 9'b100000000;
assign F[75][30] = 9'b100000000;
assign F[75][31] = 9'b100000000;
assign F[75][32] = 9'b100000000;
assign F[75][33] = 9'b100000000;
assign F[75][34] = 9'b100000000;
assign F[75][35] = 9'b100000000;
assign F[75][36] = 9'b100000000;
assign F[75][37] = 9'b100000000;
assign F[75][38] = 9'b100000000;
assign F[75][39] = 9'b100000000;
assign F[75][40] = 9'b100000000;
assign F[75][41] = 9'b100000000;
assign F[75][42] = 9'b100000000;
assign F[75][43] = 9'b100000000;
assign F[75][44] = 9'b100000000;
assign F[75][45] = 9'b100000000;
assign F[75][46] = 9'b100000000;
assign F[75][47] = 9'b100000000;
assign F[75][48] = 9'b100000000;
assign F[75][49] = 9'b100000000;
assign F[75][50] = 9'b100000000;
assign F[75][51] = 9'b100000000;
assign F[75][52] = 9'b100000000;
assign F[75][53] = 9'b100000000;
assign F[75][54] = 9'b100000000;
assign F[75][55] = 9'b100000000;
assign F[75][56] = 9'b100000000;
assign F[75][57] = 9'b100000000;
assign F[75][58] = 9'b100000000;
assign F[75][59] = 9'b100000000;
assign F[75][60] = 9'b100000000;
assign F[75][61] = 9'b100000000;
assign F[75][62] = 9'b100000000;
assign F[75][63] = 9'b100000000;
assign F[75][64] = 9'b100000000;
assign F[75][65] = 9'b100000000;
assign F[75][66] = 9'b101001000;
assign F[75][67] = 9'b100000000;
assign F[75][68] = 9'b100000000;
assign F[75][69] = 9'b100000000;
assign F[75][70] = 9'b100000000;
assign F[75][71] = 9'b100000000;
assign F[75][72] = 9'b100000000;
assign F[75][73] = 9'b100000000;
assign F[75][74] = 9'b100000000;
assign F[75][75] = 9'b100000000;
assign F[75][76] = 9'b100000000;
assign F[75][77] = 9'b100000000;
assign F[75][78] = 9'b100000000;
assign F[75][79] = 9'b100000000;
assign F[75][80] = 9'b100000000;
assign F[75][81] = 9'b100000000;
assign F[75][82] = 9'b100000000;
assign F[75][83] = 9'b100000000;
assign F[76][9] = 9'b100000000;
assign F[76][10] = 9'b100000000;
assign F[76][11] = 9'b100000000;
assign F[76][12] = 9'b100100100;
assign F[76][13] = 9'b100100100;
assign F[76][14] = 9'b100100100;
assign F[76][15] = 9'b100100100;
assign F[76][16] = 9'b100100100;
assign F[76][17] = 9'b100100100;
assign F[76][18] = 9'b100100100;
assign F[76][19] = 9'b100100100;
assign F[76][20] = 9'b100100100;
assign F[76][21] = 9'b100100100;
assign F[76][22] = 9'b100100100;
assign F[76][23] = 9'b100000000;
assign F[76][24] = 9'b100100100;
assign F[76][25] = 9'b100100100;
assign F[76][26] = 9'b100000000;
assign F[76][27] = 9'b100000000;
assign F[76][28] = 9'b100000000;
assign F[76][29] = 9'b100000000;
assign F[76][30] = 9'b100000000;
assign F[76][31] = 9'b100000000;
assign F[76][32] = 9'b100000000;
assign F[76][33] = 9'b100000000;
assign F[76][34] = 9'b100000000;
assign F[76][35] = 9'b100000000;
assign F[76][36] = 9'b100000000;
assign F[76][37] = 9'b100000000;
assign F[76][38] = 9'b100000000;
assign F[76][39] = 9'b100000000;
assign F[76][40] = 9'b100000000;
assign F[76][41] = 9'b100000000;
assign F[76][42] = 9'b100000000;
assign F[76][43] = 9'b100000000;
assign F[76][44] = 9'b100000000;
assign F[76][45] = 9'b100000000;
assign F[76][46] = 9'b100000000;
assign F[76][47] = 9'b100000000;
assign F[76][48] = 9'b100000000;
assign F[76][49] = 9'b100000000;
assign F[76][50] = 9'b100000000;
assign F[76][51] = 9'b100000000;
assign F[76][52] = 9'b100000000;
assign F[76][53] = 9'b100000000;
assign F[76][54] = 9'b100000000;
assign F[76][55] = 9'b100000000;
assign F[76][56] = 9'b100000000;
assign F[76][57] = 9'b100000000;
assign F[76][58] = 9'b100000000;
assign F[76][59] = 9'b100000000;
assign F[76][60] = 9'b100000000;
assign F[76][61] = 9'b100000000;
assign F[76][62] = 9'b100000000;
assign F[76][63] = 9'b100000000;
assign F[76][64] = 9'b100000000;
assign F[76][65] = 9'b100000000;
assign F[76][66] = 9'b100000000;
assign F[76][67] = 9'b100000000;
assign F[76][68] = 9'b100000000;
assign F[76][69] = 9'b100000000;
assign F[76][70] = 9'b100000000;
assign F[76][71] = 9'b100000000;
assign F[76][72] = 9'b100000000;
assign F[76][73] = 9'b100000000;
assign F[76][74] = 9'b100000000;
assign F[76][75] = 9'b100000000;
assign F[76][76] = 9'b100000000;
assign F[76][77] = 9'b100000000;
assign F[76][78] = 9'b100000000;
assign F[76][79] = 9'b100000000;
assign F[76][80] = 9'b100000000;
assign F[76][81] = 9'b100000000;
assign F[76][82] = 9'b100000000;
assign F[76][83] = 9'b100000000;
assign F[77][9] = 9'b100000000;
assign F[77][10] = 9'b100000000;
assign F[77][11] = 9'b100000000;
assign F[77][12] = 9'b100100100;
assign F[77][13] = 9'b100100100;
assign F[77][14] = 9'b100100100;
assign F[77][15] = 9'b100100100;
assign F[77][16] = 9'b100100100;
assign F[77][17] = 9'b100100100;
assign F[77][18] = 9'b101001000;
assign F[77][19] = 9'b101001001;
assign F[77][20] = 9'b101001001;
assign F[77][21] = 9'b100100100;
assign F[77][22] = 9'b100100100;
assign F[77][23] = 9'b100000000;
assign F[77][24] = 9'b100100100;
assign F[77][25] = 9'b100100100;
assign F[77][26] = 9'b100100100;
assign F[77][27] = 9'b100100100;
assign F[77][28] = 9'b100000000;
assign F[77][29] = 9'b100000000;
assign F[77][30] = 9'b100000000;
assign F[77][31] = 9'b100000000;
assign F[77][32] = 9'b100000000;
assign F[77][33] = 9'b100000000;
assign F[77][34] = 9'b100000000;
assign F[77][35] = 9'b100000000;
assign F[77][36] = 9'b100000000;
assign F[77][37] = 9'b100000000;
assign F[77][38] = 9'b100000000;
assign F[77][39] = 9'b100000000;
assign F[77][40] = 9'b100000000;
assign F[77][41] = 9'b100000000;
assign F[77][42] = 9'b100000000;
assign F[77][43] = 9'b100000000;
assign F[77][44] = 9'b100000000;
assign F[77][45] = 9'b100000000;
assign F[77][46] = 9'b100000000;
assign F[77][47] = 9'b100000000;
assign F[77][48] = 9'b100000000;
assign F[77][49] = 9'b100000000;
assign F[77][50] = 9'b100000000;
assign F[77][51] = 9'b100000000;
assign F[77][52] = 9'b100000000;
assign F[77][53] = 9'b100000000;
assign F[77][54] = 9'b100000000;
assign F[77][55] = 9'b100000000;
assign F[77][56] = 9'b100000000;
assign F[77][57] = 9'b100000000;
assign F[77][58] = 9'b100000000;
assign F[77][59] = 9'b100000000;
assign F[77][60] = 9'b100000000;
assign F[77][61] = 9'b100000000;
assign F[77][62] = 9'b100000000;
assign F[77][63] = 9'b100000000;
assign F[77][64] = 9'b100000000;
assign F[77][65] = 9'b100000000;
assign F[77][66] = 9'b100000000;
assign F[77][67] = 9'b100000000;
assign F[77][68] = 9'b100000000;
assign F[77][69] = 9'b100000000;
assign F[77][70] = 9'b100000000;
assign F[77][71] = 9'b100000000;
assign F[77][72] = 9'b100000000;
assign F[77][73] = 9'b100000000;
assign F[77][74] = 9'b100000000;
assign F[77][75] = 9'b100000000;
assign F[77][76] = 9'b100000000;
assign F[77][77] = 9'b100000000;
assign F[77][78] = 9'b100000000;
assign F[77][79] = 9'b100000000;
assign F[77][80] = 9'b100000000;
assign F[77][81] = 9'b100100100;
assign F[77][82] = 9'b100100100;
assign F[77][83] = 9'b100000000;
assign F[78][9] = 9'b100000000;
assign F[78][10] = 9'b100000000;
assign F[78][11] = 9'b101001001;
assign F[78][12] = 9'b101001001;
assign F[78][13] = 9'b101001001;
assign F[78][14] = 9'b101001001;
assign F[78][15] = 9'b101001001;
assign F[78][16] = 9'b101001001;
assign F[78][17] = 9'b101001001;
assign F[78][18] = 9'b101101101;
assign F[78][19] = 9'b110010001;
assign F[78][20] = 9'b101101101;
assign F[78][21] = 9'b100100100;
assign F[78][22] = 9'b100000000;
assign F[78][23] = 9'b100100100;
assign F[78][24] = 9'b100100100;
assign F[78][25] = 9'b100100100;
assign F[78][26] = 9'b100100100;
assign F[78][27] = 9'b100100100;
assign F[78][28] = 9'b100000000;
assign F[78][29] = 9'b100000000;
assign F[78][30] = 9'b100000000;
assign F[78][31] = 9'b100000000;
assign F[78][32] = 9'b100000000;
assign F[78][33] = 9'b100000000;
assign F[78][34] = 9'b100000000;
assign F[78][35] = 9'b100000000;
assign F[78][36] = 9'b100000000;
assign F[78][37] = 9'b100000000;
assign F[78][38] = 9'b100000000;
assign F[78][39] = 9'b100000000;
assign F[78][40] = 9'b100000000;
assign F[78][41] = 9'b100000000;
assign F[78][42] = 9'b100000000;
assign F[78][43] = 9'b100000000;
assign F[78][44] = 9'b100000000;
assign F[78][45] = 9'b100000000;
assign F[78][46] = 9'b100000000;
assign F[78][47] = 9'b100000000;
assign F[78][48] = 9'b100000000;
assign F[78][49] = 9'b100000000;
assign F[78][50] = 9'b100000000;
assign F[78][51] = 9'b100000000;
assign F[78][52] = 9'b100000000;
assign F[78][53] = 9'b100000000;
assign F[78][54] = 9'b100000000;
assign F[78][55] = 9'b100000000;
assign F[78][56] = 9'b100000000;
assign F[78][57] = 9'b100000000;
assign F[78][58] = 9'b100000000;
assign F[78][59] = 9'b100000000;
assign F[78][60] = 9'b100000000;
assign F[78][61] = 9'b100000000;
assign F[78][62] = 9'b100000000;
assign F[78][63] = 9'b100000000;
assign F[78][64] = 9'b100000000;
assign F[78][65] = 9'b100000000;
assign F[78][66] = 9'b100000000;
assign F[78][67] = 9'b100000000;
assign F[78][68] = 9'b100000000;
assign F[78][69] = 9'b100000000;
assign F[78][70] = 9'b100000000;
assign F[78][71] = 9'b100000000;
assign F[78][72] = 9'b100000000;
assign F[78][73] = 9'b100000000;
assign F[78][74] = 9'b100000000;
assign F[78][75] = 9'b100000000;
assign F[78][76] = 9'b100000000;
assign F[78][77] = 9'b100000000;
assign F[78][78] = 9'b100000000;
assign F[78][79] = 9'b100000000;
assign F[78][80] = 9'b100000000;
assign F[78][81] = 9'b101101101;
assign F[78][82] = 9'b101001000;
assign F[78][83] = 9'b100000000;
assign F[79][8] = 9'b100000000;
assign F[79][9] = 9'b100000000;
assign F[79][10] = 9'b100100100;
assign F[79][11] = 9'b110010001;
assign F[79][12] = 9'b101101101;
assign F[79][13] = 9'b101101101;
assign F[79][14] = 9'b101101101;
assign F[79][15] = 9'b101101101;
assign F[79][16] = 9'b101101101;
assign F[79][17] = 9'b101101101;
assign F[79][18] = 9'b110010001;
assign F[79][19] = 9'b110010001;
assign F[79][20] = 9'b101101101;
assign F[79][21] = 9'b100100100;
assign F[79][22] = 9'b100000000;
assign F[79][23] = 9'b100100100;
assign F[79][24] = 9'b100100100;
assign F[79][25] = 9'b100100100;
assign F[79][26] = 9'b100100100;
assign F[79][27] = 9'b100100100;
assign F[79][28] = 9'b100100100;
assign F[79][29] = 9'b100100100;
assign F[79][30] = 9'b100000000;
assign F[79][31] = 9'b100000000;
assign F[79][32] = 9'b100000000;
assign F[79][33] = 9'b100000000;
assign F[79][34] = 9'b100000000;
assign F[79][35] = 9'b100000000;
assign F[79][36] = 9'b100000000;
assign F[79][37] = 9'b100000000;
assign F[79][38] = 9'b100000000;
assign F[79][39] = 9'b100000000;
assign F[79][40] = 9'b100000000;
assign F[79][41] = 9'b100000000;
assign F[79][42] = 9'b100000000;
assign F[79][43] = 9'b100000000;
assign F[79][44] = 9'b100000000;
assign F[79][45] = 9'b100000000;
assign F[79][46] = 9'b100000000;
assign F[79][47] = 9'b100000000;
assign F[79][48] = 9'b100000000;
assign F[79][49] = 9'b100000000;
assign F[79][50] = 9'b100000000;
assign F[79][51] = 9'b100000000;
assign F[79][52] = 9'b100000000;
assign F[79][53] = 9'b100000000;
assign F[79][54] = 9'b100000000;
assign F[79][55] = 9'b100000000;
assign F[79][56] = 9'b100000000;
assign F[79][57] = 9'b100000000;
assign F[79][58] = 9'b100000000;
assign F[79][59] = 9'b100000000;
assign F[79][60] = 9'b100000000;
assign F[79][61] = 9'b100000000;
assign F[79][62] = 9'b100000000;
assign F[79][63] = 9'b100000000;
assign F[79][64] = 9'b100000000;
assign F[79][65] = 9'b100000000;
assign F[79][66] = 9'b100000000;
assign F[79][67] = 9'b100000000;
assign F[79][68] = 9'b100000000;
assign F[79][69] = 9'b100000000;
assign F[79][70] = 9'b100000000;
assign F[79][71] = 9'b100000000;
assign F[79][72] = 9'b100000000;
assign F[79][73] = 9'b100000000;
assign F[79][74] = 9'b100000000;
assign F[79][75] = 9'b100000000;
assign F[79][76] = 9'b100000000;
assign F[79][77] = 9'b100000000;
assign F[79][78] = 9'b100000000;
assign F[79][79] = 9'b100000000;
assign F[79][80] = 9'b100000000;
assign F[79][81] = 9'b101101101;
assign F[79][82] = 9'b100100100;
assign F[79][83] = 9'b100000000;
assign F[80][7] = 9'b100000000;
assign F[80][8] = 9'b100000000;
assign F[80][9] = 9'b100100100;
assign F[80][10] = 9'b101001000;
assign F[80][11] = 9'b101101101;
assign F[80][12] = 9'b101101101;
assign F[80][13] = 9'b101101101;
assign F[80][14] = 9'b101101101;
assign F[80][15] = 9'b101001001;
assign F[80][16] = 9'b101001001;
assign F[80][17] = 9'b101001001;
assign F[80][18] = 9'b101101101;
assign F[80][19] = 9'b101101101;
assign F[80][20] = 9'b101001001;
assign F[80][21] = 9'b100100100;
assign F[80][22] = 9'b100000000;
assign F[80][23] = 9'b100100100;
assign F[80][24] = 9'b100100100;
assign F[80][25] = 9'b100100100;
assign F[80][26] = 9'b100100100;
assign F[80][27] = 9'b100100100;
assign F[80][28] = 9'b100100100;
assign F[80][29] = 9'b100100100;
assign F[80][30] = 9'b100000000;
assign F[80][31] = 9'b100000000;
assign F[80][32] = 9'b100000000;
assign F[80][33] = 9'b100000000;
assign F[80][34] = 9'b100000000;
assign F[80][35] = 9'b100000000;
assign F[80][36] = 9'b100000000;
assign F[80][37] = 9'b100000000;
assign F[80][38] = 9'b100000000;
assign F[80][39] = 9'b100000000;
assign F[80][40] = 9'b100000000;
assign F[80][41] = 9'b100000000;
assign F[80][42] = 9'b100000000;
assign F[80][43] = 9'b100000000;
assign F[80][44] = 9'b100000000;
assign F[80][45] = 9'b100000000;
assign F[80][46] = 9'b100000000;
assign F[80][47] = 9'b100000000;
assign F[80][48] = 9'b100000000;
assign F[80][49] = 9'b100100100;
assign F[80][50] = 9'b100100100;
assign F[80][51] = 9'b100000000;
assign F[80][52] = 9'b100000000;
assign F[80][53] = 9'b100000000;
assign F[80][54] = 9'b100000000;
assign F[80][55] = 9'b100000000;
assign F[80][56] = 9'b100000000;
assign F[80][57] = 9'b100000000;
assign F[80][58] = 9'b100000000;
assign F[80][59] = 9'b100000000;
assign F[80][60] = 9'b100000000;
assign F[80][61] = 9'b100000000;
assign F[80][62] = 9'b100000000;
assign F[80][63] = 9'b100000000;
assign F[80][64] = 9'b100000000;
assign F[80][65] = 9'b100000000;
assign F[80][66] = 9'b100000000;
assign F[80][67] = 9'b100000000;
assign F[80][68] = 9'b100000000;
assign F[80][69] = 9'b100000000;
assign F[80][70] = 9'b100000000;
assign F[80][71] = 9'b100000000;
assign F[80][72] = 9'b100000000;
assign F[80][73] = 9'b100000000;
assign F[80][74] = 9'b100000000;
assign F[80][75] = 9'b100000000;
assign F[80][76] = 9'b100000000;
assign F[80][77] = 9'b100000000;
assign F[80][78] = 9'b100000000;
assign F[80][79] = 9'b100000000;
assign F[80][80] = 9'b100000000;
assign F[80][81] = 9'b100100100;
assign F[80][82] = 9'b100000000;
assign F[80][83] = 9'b100000000;
assign F[81][8] = 9'b100000000;
assign F[81][9] = 9'b100100100;
assign F[81][10] = 9'b100100100;
assign F[81][11] = 9'b100100100;
assign F[81][12] = 9'b100100100;
assign F[81][13] = 9'b100100100;
assign F[81][14] = 9'b100100100;
assign F[81][15] = 9'b100100100;
assign F[81][16] = 9'b100100100;
assign F[81][17] = 9'b100100100;
assign F[81][18] = 9'b101001000;
assign F[81][19] = 9'b101001001;
assign F[81][20] = 9'b100100100;
assign F[81][21] = 9'b100100100;
assign F[81][22] = 9'b100100100;
assign F[81][23] = 9'b100100100;
assign F[81][24] = 9'b100100100;
assign F[81][25] = 9'b100100100;
assign F[81][26] = 9'b100100100;
assign F[81][27] = 9'b100100100;
assign F[81][28] = 9'b100100100;
assign F[81][29] = 9'b100100100;
assign F[81][30] = 9'b100100100;
assign F[81][31] = 9'b100100100;
assign F[81][32] = 9'b100000000;
assign F[81][33] = 9'b100000000;
assign F[81][34] = 9'b100000000;
assign F[81][35] = 9'b100000000;
assign F[81][36] = 9'b100000000;
assign F[81][37] = 9'b100000000;
assign F[81][38] = 9'b100000000;
assign F[81][39] = 9'b100000000;
assign F[81][40] = 9'b100000000;
assign F[81][41] = 9'b100000000;
assign F[81][42] = 9'b100000000;
assign F[81][43] = 9'b100000000;
assign F[81][44] = 9'b100000000;
assign F[81][45] = 9'b100000000;
assign F[81][46] = 9'b100000000;
assign F[81][47] = 9'b100000000;
assign F[81][48] = 9'b100100100;
assign F[81][49] = 9'b110010001;
assign F[81][50] = 9'b101001001;
assign F[81][51] = 9'b100000000;
assign F[81][52] = 9'b100000000;
assign F[81][53] = 9'b100000000;
assign F[81][54] = 9'b100000000;
assign F[81][55] = 9'b100000000;
assign F[81][56] = 9'b100000000;
assign F[81][57] = 9'b100000000;
assign F[81][58] = 9'b100000000;
assign F[81][59] = 9'b100000000;
assign F[81][60] = 9'b100000000;
assign F[81][61] = 9'b100000000;
assign F[81][62] = 9'b100000000;
assign F[81][63] = 9'b100000000;
assign F[81][64] = 9'b100000000;
assign F[81][65] = 9'b100000000;
assign F[81][66] = 9'b100000000;
assign F[81][67] = 9'b100000000;
assign F[81][68] = 9'b100000000;
assign F[81][69] = 9'b100000000;
assign F[81][70] = 9'b100000000;
assign F[81][71] = 9'b100000000;
assign F[81][72] = 9'b100000000;
assign F[81][73] = 9'b100000000;
assign F[81][74] = 9'b100000000;
assign F[81][75] = 9'b100000000;
assign F[81][76] = 9'b100000000;
assign F[81][77] = 9'b100000000;
assign F[81][78] = 9'b100000000;
assign F[81][79] = 9'b100000000;
assign F[81][80] = 9'b100000000;
assign F[81][81] = 9'b100000000;
assign F[81][82] = 9'b100000000;
assign F[81][83] = 9'b100000000;
assign F[81][84] = 9'b100000000;
assign F[82][8] = 9'b100000000;
assign F[82][9] = 9'b100000000;
assign F[82][10] = 9'b100100100;
assign F[82][11] = 9'b100100100;
assign F[82][12] = 9'b100100100;
assign F[82][13] = 9'b100100100;
assign F[82][14] = 9'b100100100;
assign F[82][15] = 9'b100100100;
assign F[82][16] = 9'b100100100;
assign F[82][17] = 9'b100100100;
assign F[82][18] = 9'b100100100;
assign F[82][19] = 9'b100000000;
assign F[82][20] = 9'b100100100;
assign F[82][21] = 9'b100100100;
assign F[82][22] = 9'b100100100;
assign F[82][23] = 9'b100100100;
assign F[82][24] = 9'b100100100;
assign F[82][25] = 9'b100100100;
assign F[82][26] = 9'b100100100;
assign F[82][27] = 9'b100100100;
assign F[82][28] = 9'b100100100;
assign F[82][29] = 9'b100100100;
assign F[82][30] = 9'b100100100;
assign F[82][31] = 9'b100000000;
assign F[82][32] = 9'b100000000;
assign F[82][33] = 9'b100000000;
assign F[82][34] = 9'b100000000;
assign F[82][35] = 9'b100000000;
assign F[82][36] = 9'b100000000;
assign F[82][37] = 9'b100000000;
assign F[82][38] = 9'b100000000;
assign F[82][39] = 9'b100000000;
assign F[82][40] = 9'b100000000;
assign F[82][41] = 9'b100000000;
assign F[82][42] = 9'b100000000;
assign F[82][43] = 9'b100000000;
assign F[82][44] = 9'b100000000;
assign F[82][45] = 9'b100000000;
assign F[82][46] = 9'b100000000;
assign F[82][47] = 9'b101001001;
assign F[82][48] = 9'b101110001;
assign F[82][49] = 9'b101101101;
assign F[82][50] = 9'b101001001;
assign F[82][51] = 9'b100100100;
assign F[82][52] = 9'b100000000;
assign F[82][53] = 9'b100000000;
assign F[82][54] = 9'b100000000;
assign F[82][55] = 9'b100000000;
assign F[82][56] = 9'b100000000;
assign F[82][57] = 9'b100000000;
assign F[82][58] = 9'b100000000;
assign F[82][59] = 9'b100000000;
assign F[82][60] = 9'b100000000;
assign F[82][61] = 9'b100000000;
assign F[82][62] = 9'b100000000;
assign F[82][63] = 9'b100000000;
assign F[82][64] = 9'b100000000;
assign F[82][65] = 9'b100000000;
assign F[82][66] = 9'b100000000;
assign F[82][67] = 9'b100000000;
assign F[82][68] = 9'b100000000;
assign F[82][69] = 9'b100000000;
assign F[82][70] = 9'b100000000;
assign F[82][71] = 9'b100000000;
assign F[82][72] = 9'b100000000;
assign F[82][73] = 9'b100000000;
assign F[82][74] = 9'b100000000;
assign F[82][75] = 9'b100000000;
assign F[82][76] = 9'b100000000;
assign F[82][77] = 9'b100000000;
assign F[82][78] = 9'b100000000;
assign F[82][79] = 9'b100000000;
assign F[82][80] = 9'b100000000;
assign F[82][81] = 9'b100000000;
assign F[82][82] = 9'b100000000;
assign F[82][83] = 9'b100000000;
assign F[82][84] = 9'b100000000;
assign F[82][85] = 9'b100000000;
assign F[83][8] = 9'b100000000;
assign F[83][9] = 9'b100000000;
assign F[83][10] = 9'b100100100;
assign F[83][11] = 9'b100100100;
assign F[83][12] = 9'b100100100;
assign F[83][13] = 9'b100100100;
assign F[83][14] = 9'b100100100;
assign F[83][15] = 9'b100100100;
assign F[83][16] = 9'b100100100;
assign F[83][17] = 9'b100100100;
assign F[83][18] = 9'b100100100;
assign F[83][19] = 9'b100100100;
assign F[83][20] = 9'b100100100;
assign F[83][21] = 9'b100100100;
assign F[83][22] = 9'b100100100;
assign F[83][23] = 9'b100100100;
assign F[83][24] = 9'b100100100;
assign F[83][25] = 9'b100000000;
assign F[83][26] = 9'b100100100;
assign F[83][27] = 9'b100100100;
assign F[83][28] = 9'b100100100;
assign F[83][29] = 9'b100100100;
assign F[83][30] = 9'b100100100;
assign F[83][31] = 9'b100000000;
assign F[83][32] = 9'b100000000;
assign F[83][33] = 9'b100000000;
assign F[83][34] = 9'b100000000;
assign F[83][35] = 9'b100000000;
assign F[83][36] = 9'b100000000;
assign F[83][37] = 9'b100000000;
assign F[83][38] = 9'b100000000;
assign F[83][39] = 9'b100000000;
assign F[83][40] = 9'b100000000;
assign F[83][41] = 9'b100000000;
assign F[83][42] = 9'b100000000;
assign F[83][43] = 9'b100000000;
assign F[83][44] = 9'b100000000;
assign F[83][45] = 9'b100000000;
assign F[83][46] = 9'b100000000;
assign F[83][47] = 9'b101001001;
assign F[83][48] = 9'b101101101;
assign F[83][49] = 9'b101101101;
assign F[83][50] = 9'b101101101;
assign F[83][51] = 9'b101101001;
assign F[83][52] = 9'b101101001;
assign F[83][53] = 9'b101000100;
assign F[83][54] = 9'b100000000;
assign F[83][55] = 9'b100000000;
assign F[83][56] = 9'b100000000;
assign F[83][57] = 9'b100000000;
assign F[83][58] = 9'b100000000;
assign F[83][59] = 9'b100000000;
assign F[83][60] = 9'b100000000;
assign F[83][61] = 9'b100000000;
assign F[83][62] = 9'b100000000;
assign F[83][63] = 9'b100000000;
assign F[83][64] = 9'b100000000;
assign F[83][65] = 9'b100000000;
assign F[83][66] = 9'b100000000;
assign F[83][67] = 9'b100000000;
assign F[83][68] = 9'b100000000;
assign F[83][69] = 9'b100000000;
assign F[83][70] = 9'b100000000;
assign F[83][71] = 9'b100000000;
assign F[83][72] = 9'b100000000;
assign F[83][73] = 9'b100000000;
assign F[83][74] = 9'b100000000;
assign F[83][75] = 9'b100000000;
assign F[83][76] = 9'b100000000;
assign F[83][77] = 9'b100000000;
assign F[83][78] = 9'b100000000;
assign F[83][79] = 9'b100000000;
assign F[83][80] = 9'b100000000;
assign F[83][81] = 9'b100000000;
assign F[83][82] = 9'b100000000;
assign F[83][83] = 9'b100000000;
assign F[83][84] = 9'b100000000;
assign F[83][85] = 9'b100000000;
assign F[84][7] = 9'b100000000;
assign F[84][8] = 9'b100000000;
assign F[84][9] = 9'b100000000;
assign F[84][10] = 9'b100100100;
assign F[84][11] = 9'b100100100;
assign F[84][12] = 9'b100100100;
assign F[84][13] = 9'b100100100;
assign F[84][14] = 9'b100100100;
assign F[84][15] = 9'b100100100;
assign F[84][16] = 9'b100100100;
assign F[84][17] = 9'b100100100;
assign F[84][18] = 9'b100100100;
assign F[84][19] = 9'b100100100;
assign F[84][20] = 9'b100100100;
assign F[84][21] = 9'b100100100;
assign F[84][22] = 9'b100100100;
assign F[84][23] = 9'b100100100;
assign F[84][24] = 9'b100100100;
assign F[84][25] = 9'b100100100;
assign F[84][26] = 9'b100100100;
assign F[84][27] = 9'b100100100;
assign F[84][28] = 9'b100100100;
assign F[84][29] = 9'b100100100;
assign F[84][30] = 9'b100100100;
assign F[84][31] = 9'b100100100;
assign F[84][32] = 9'b100000000;
assign F[84][33] = 9'b100000000;
assign F[84][34] = 9'b100000000;
assign F[84][35] = 9'b100000000;
assign F[84][36] = 9'b100000000;
assign F[84][37] = 9'b100000000;
assign F[84][38] = 9'b100000000;
assign F[84][39] = 9'b100000000;
assign F[84][40] = 9'b100000000;
assign F[84][41] = 9'b100000000;
assign F[84][42] = 9'b100000000;
assign F[84][43] = 9'b100000000;
assign F[84][44] = 9'b100000000;
assign F[84][45] = 9'b100000000;
assign F[84][46] = 9'b100000000;
assign F[84][47] = 9'b100100100;
assign F[84][48] = 9'b101001001;
assign F[84][49] = 9'b101101001;
assign F[84][50] = 9'b101101001;
assign F[84][51] = 9'b110001001;
assign F[84][52] = 9'b110001001;
assign F[84][53] = 9'b101000100;
assign F[84][54] = 9'b100000000;
assign F[84][55] = 9'b100000000;
assign F[84][56] = 9'b100000000;
assign F[84][57] = 9'b100000000;
assign F[84][58] = 9'b100000000;
assign F[84][59] = 9'b100000000;
assign F[84][60] = 9'b100000000;
assign F[84][61] = 9'b100000000;
assign F[84][62] = 9'b100000000;
assign F[84][63] = 9'b100000000;
assign F[84][64] = 9'b100000000;
assign F[84][65] = 9'b100000000;
assign F[84][66] = 9'b100000000;
assign F[84][67] = 9'b100000000;
assign F[84][68] = 9'b100000000;
assign F[84][69] = 9'b100000000;
assign F[84][70] = 9'b100000000;
assign F[84][71] = 9'b100000000;
assign F[84][72] = 9'b100000000;
assign F[84][73] = 9'b100000000;
assign F[84][74] = 9'b100000000;
assign F[84][75] = 9'b100000000;
assign F[84][76] = 9'b100000000;
assign F[84][77] = 9'b100000000;
assign F[84][78] = 9'b100000000;
assign F[84][79] = 9'b100000000;
assign F[84][80] = 9'b100000000;
assign F[84][81] = 9'b100000000;
assign F[84][82] = 9'b100100100;
assign F[84][83] = 9'b100000000;
assign F[84][84] = 9'b100000000;
assign F[84][85] = 9'b100000000;
assign F[85][8] = 9'b100000000;
assign F[85][9] = 9'b100000000;
assign F[85][10] = 9'b100000000;
assign F[85][11] = 9'b101001001;
assign F[85][12] = 9'b101001001;
assign F[85][13] = 9'b101001001;
assign F[85][14] = 9'b101001001;
assign F[85][15] = 9'b101001001;
assign F[85][16] = 9'b101001001;
assign F[85][17] = 9'b101001001;
assign F[85][18] = 9'b101001001;
assign F[85][19] = 9'b101001000;
assign F[85][20] = 9'b100100100;
assign F[85][21] = 9'b100100100;
assign F[85][22] = 9'b100100100;
assign F[85][23] = 9'b100100100;
assign F[85][24] = 9'b100100100;
assign F[85][25] = 9'b100100100;
assign F[85][26] = 9'b100100100;
assign F[85][27] = 9'b100100100;
assign F[85][28] = 9'b100000000;
assign F[85][29] = 9'b100000000;
assign F[85][30] = 9'b100100100;
assign F[85][31] = 9'b100100100;
assign F[85][32] = 9'b100100100;
assign F[85][33] = 9'b100000000;
assign F[85][34] = 9'b100000000;
assign F[85][35] = 9'b100000000;
assign F[85][36] = 9'b100000000;
assign F[85][37] = 9'b100000000;
assign F[85][38] = 9'b100000000;
assign F[85][39] = 9'b100000000;
assign F[85][40] = 9'b100000000;
assign F[85][41] = 9'b100000000;
assign F[85][42] = 9'b100000000;
assign F[85][43] = 9'b100000000;
assign F[85][44] = 9'b100000000;
assign F[85][45] = 9'b100000000;
assign F[85][46] = 9'b100000000;
assign F[85][47] = 9'b100100100;
assign F[85][48] = 9'b101001000;
assign F[85][49] = 9'b101001001;
assign F[85][50] = 9'b101000100;
assign F[85][51] = 9'b101000100;
assign F[85][52] = 9'b101000100;
assign F[85][53] = 9'b100100100;
assign F[85][54] = 9'b100000000;
assign F[85][55] = 9'b100000000;
assign F[85][56] = 9'b100000000;
assign F[85][57] = 9'b100000000;
assign F[85][58] = 9'b100000000;
assign F[85][59] = 9'b100000000;
assign F[85][60] = 9'b100000000;
assign F[85][61] = 9'b100000000;
assign F[85][62] = 9'b100000000;
assign F[85][63] = 9'b100000000;
assign F[85][64] = 9'b100000000;
assign F[85][65] = 9'b100000000;
assign F[85][66] = 9'b100000000;
assign F[85][67] = 9'b100000000;
assign F[85][68] = 9'b100000000;
assign F[85][69] = 9'b100000000;
assign F[85][70] = 9'b100000000;
assign F[85][71] = 9'b100000000;
assign F[85][72] = 9'b100000000;
assign F[85][73] = 9'b100000000;
assign F[85][74] = 9'b100000000;
assign F[85][75] = 9'b100000000;
assign F[85][76] = 9'b100000000;
assign F[85][77] = 9'b100000000;
assign F[85][78] = 9'b100000000;
assign F[85][79] = 9'b100000000;
assign F[85][80] = 9'b100000000;
assign F[85][81] = 9'b100000000;
assign F[85][82] = 9'b100000000;
assign F[85][83] = 9'b100000000;
assign F[85][84] = 9'b100000000;
assign F[85][85] = 9'b100000000;
assign F[85][86] = 9'b100000000;
assign F[86][9] = 9'b100000000;
assign F[86][10] = 9'b100000000;
assign F[86][11] = 9'b110010001;
assign F[86][12] = 9'b101101101;
assign F[86][13] = 9'b101101101;
assign F[86][14] = 9'b101101101;
assign F[86][15] = 9'b101101101;
assign F[86][16] = 9'b101101101;
assign F[86][17] = 9'b101101101;
assign F[86][18] = 9'b101101101;
assign F[86][19] = 9'b101101101;
assign F[86][20] = 9'b100100100;
assign F[86][21] = 9'b100100100;
assign F[86][22] = 9'b100100100;
assign F[86][23] = 9'b100100100;
assign F[86][24] = 9'b100100100;
assign F[86][25] = 9'b100100100;
assign F[86][26] = 9'b100100100;
assign F[86][27] = 9'b100100100;
assign F[86][28] = 9'b100000000;
assign F[86][29] = 9'b100000000;
assign F[86][30] = 9'b100100100;
assign F[86][31] = 9'b100100100;
assign F[86][32] = 9'b100100100;
assign F[86][33] = 9'b100000000;
assign F[86][34] = 9'b100000000;
assign F[86][35] = 9'b100000000;
assign F[86][36] = 9'b100000000;
assign F[86][37] = 9'b100000000;
assign F[86][38] = 9'b100000000;
assign F[86][39] = 9'b100000000;
assign F[86][40] = 9'b100000000;
assign F[86][41] = 9'b100000000;
assign F[86][42] = 9'b100000000;
assign F[86][43] = 9'b100000000;
assign F[86][44] = 9'b100000000;
assign F[86][45] = 9'b100000000;
assign F[86][46] = 9'b100000000;
assign F[86][47] = 9'b100000100;
assign F[86][48] = 9'b100100100;
assign F[86][49] = 9'b100100100;
assign F[86][50] = 9'b100000000;
assign F[86][51] = 9'b100000000;
assign F[86][52] = 9'b100000000;
assign F[86][53] = 9'b100000000;
assign F[86][54] = 9'b100000000;
assign F[86][55] = 9'b100000000;
assign F[86][56] = 9'b100000000;
assign F[86][57] = 9'b100000000;
assign F[86][58] = 9'b100000000;
assign F[86][59] = 9'b100000000;
assign F[86][60] = 9'b100000000;
assign F[86][61] = 9'b100000000;
assign F[86][62] = 9'b100000000;
assign F[86][63] = 9'b100000000;
assign F[86][64] = 9'b100000000;
assign F[86][65] = 9'b100000000;
assign F[86][66] = 9'b100000000;
assign F[86][67] = 9'b100000000;
assign F[86][68] = 9'b100000000;
assign F[86][69] = 9'b100000000;
assign F[86][70] = 9'b100000000;
assign F[86][71] = 9'b100000000;
assign F[86][72] = 9'b100000000;
assign F[86][73] = 9'b100000000;
assign F[86][74] = 9'b100000000;
assign F[86][75] = 9'b100000000;
assign F[86][76] = 9'b100000000;
assign F[86][77] = 9'b100000000;
assign F[86][78] = 9'b100000000;
assign F[86][79] = 9'b100000000;
assign F[86][80] = 9'b100000000;
assign F[86][81] = 9'b100000000;
assign F[86][82] = 9'b100000000;
assign F[86][83] = 9'b100100100;
assign F[86][84] = 9'b100100100;
assign F[86][85] = 9'b100000000;
assign F[86][86] = 9'b100000000;
assign F[87][9] = 9'b100000000;
assign F[87][10] = 9'b100000000;
assign F[87][11] = 9'b101101101;
assign F[87][12] = 9'b101001001;
assign F[87][13] = 9'b101001001;
assign F[87][14] = 9'b101001001;
assign F[87][15] = 9'b101001001;
assign F[87][16] = 9'b101001001;
assign F[87][17] = 9'b101001001;
assign F[87][18] = 9'b101001001;
assign F[87][19] = 9'b101001001;
assign F[87][20] = 9'b100100100;
assign F[87][21] = 9'b100100100;
assign F[87][22] = 9'b100100100;
assign F[87][23] = 9'b100100100;
assign F[87][24] = 9'b100100100;
assign F[87][25] = 9'b100100100;
assign F[87][26] = 9'b100100100;
assign F[87][27] = 9'b100100100;
assign F[87][28] = 9'b100000000;
assign F[87][29] = 9'b100000000;
assign F[87][30] = 9'b100000000;
assign F[87][31] = 9'b100000000;
assign F[87][32] = 9'b100000000;
assign F[87][33] = 9'b100100100;
assign F[87][34] = 9'b100100100;
assign F[87][35] = 9'b100000000;
assign F[87][36] = 9'b100000000;
assign F[87][37] = 9'b100000000;
assign F[87][38] = 9'b100000000;
assign F[87][39] = 9'b100000000;
assign F[87][40] = 9'b100000000;
assign F[87][41] = 9'b100000000;
assign F[87][42] = 9'b100000000;
assign F[87][43] = 9'b100000000;
assign F[87][44] = 9'b100000000;
assign F[87][45] = 9'b100000000;
assign F[87][46] = 9'b100000000;
assign F[87][47] = 9'b100000000;
assign F[87][48] = 9'b100000000;
assign F[87][49] = 9'b100000000;
assign F[87][50] = 9'b100000000;
assign F[87][51] = 9'b100000000;
assign F[87][52] = 9'b100000000;
assign F[87][53] = 9'b100000000;
assign F[87][54] = 9'b100000000;
assign F[87][55] = 9'b100000000;
assign F[87][56] = 9'b100000000;
assign F[87][57] = 9'b100000000;
assign F[87][58] = 9'b100000000;
assign F[87][59] = 9'b100000000;
assign F[87][60] = 9'b100000000;
assign F[87][61] = 9'b100000000;
assign F[87][62] = 9'b100000000;
assign F[87][63] = 9'b100000000;
assign F[87][64] = 9'b100000000;
assign F[87][65] = 9'b100000000;
assign F[87][66] = 9'b100000000;
assign F[87][67] = 9'b100000000;
assign F[87][68] = 9'b100000000;
assign F[87][69] = 9'b100000000;
assign F[87][70] = 9'b100000000;
assign F[87][71] = 9'b100000000;
assign F[87][72] = 9'b100000000;
assign F[87][73] = 9'b100000000;
assign F[87][74] = 9'b100000000;
assign F[87][75] = 9'b100000000;
assign F[87][76] = 9'b100000000;
assign F[87][77] = 9'b100000000;
assign F[87][78] = 9'b100000000;
assign F[87][79] = 9'b100000000;
assign F[87][80] = 9'b100000000;
assign F[87][81] = 9'b100000000;
assign F[87][82] = 9'b100000000;
assign F[87][83] = 9'b100100100;
assign F[87][84] = 9'b100100100;
assign F[87][85] = 9'b100000000;
assign F[87][86] = 9'b100000000;
assign F[88][9] = 9'b100000000;
assign F[88][10] = 9'b100000000;
assign F[88][11] = 9'b100100100;
assign F[88][12] = 9'b100100100;
assign F[88][13] = 9'b100100100;
assign F[88][14] = 9'b100000000;
assign F[88][15] = 9'b100100100;
assign F[88][16] = 9'b100100100;
assign F[88][17] = 9'b100100100;
assign F[88][18] = 9'b100100100;
assign F[88][19] = 9'b100100100;
assign F[88][20] = 9'b100100100;
assign F[88][21] = 9'b100100100;
assign F[88][22] = 9'b100100100;
assign F[88][23] = 9'b100000000;
assign F[88][24] = 9'b100100100;
assign F[88][25] = 9'b100100100;
assign F[88][26] = 9'b100000000;
assign F[88][27] = 9'b100000000;
assign F[88][28] = 9'b100000000;
assign F[88][29] = 9'b100000000;
assign F[88][30] = 9'b100000000;
assign F[88][31] = 9'b100000000;
assign F[88][32] = 9'b100000000;
assign F[88][33] = 9'b100000000;
assign F[88][34] = 9'b100000000;
assign F[88][35] = 9'b100000000;
assign F[88][36] = 9'b100000000;
assign F[88][37] = 9'b100000000;
assign F[88][38] = 9'b100000000;
assign F[88][39] = 9'b100000000;
assign F[88][40] = 9'b100000000;
assign F[88][41] = 9'b100000000;
assign F[88][42] = 9'b100000000;
assign F[88][43] = 9'b100000000;
assign F[88][44] = 9'b100000000;
assign F[88][45] = 9'b100000000;
assign F[88][46] = 9'b100000000;
assign F[88][47] = 9'b100000000;
assign F[88][48] = 9'b100000000;
assign F[88][49] = 9'b100000000;
assign F[88][50] = 9'b100000000;
assign F[88][51] = 9'b100000000;
assign F[88][52] = 9'b100000000;
assign F[88][53] = 9'b100000000;
assign F[88][54] = 9'b100000000;
assign F[88][55] = 9'b100000000;
assign F[88][56] = 9'b100000000;
assign F[88][57] = 9'b100000000;
assign F[88][58] = 9'b100000000;
assign F[88][59] = 9'b100000000;
assign F[88][60] = 9'b100000000;
assign F[88][61] = 9'b100000000;
assign F[88][62] = 9'b100000000;
assign F[88][63] = 9'b100000000;
assign F[88][64] = 9'b100000000;
assign F[88][65] = 9'b100000000;
assign F[88][66] = 9'b100000000;
assign F[88][67] = 9'b100000000;
assign F[88][68] = 9'b100000000;
assign F[88][69] = 9'b100000000;
assign F[88][70] = 9'b100000000;
assign F[88][71] = 9'b100000000;
assign F[88][72] = 9'b100000000;
assign F[88][73] = 9'b100000000;
assign F[88][74] = 9'b100000000;
assign F[88][75] = 9'b100000000;
assign F[88][76] = 9'b100000000;
assign F[88][77] = 9'b100000000;
assign F[88][78] = 9'b100000000;
assign F[88][79] = 9'b100000000;
assign F[88][80] = 9'b100000000;
assign F[88][81] = 9'b100000000;
assign F[88][82] = 9'b100000000;
assign F[88][83] = 9'b100000000;
assign F[88][84] = 9'b100100100;
assign F[88][85] = 9'b100000000;
assign F[88][86] = 9'b100000000;
//Total de Lineas = 3655
endmodule*/

