`timescale 1ns / 1ps
module prueba_4 (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (micromatriz[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= micromatriz[vcount- posy][hcount- posx][7:5];
				green <= micromatriz[vcount- posy][hcount- posx][4:2];
            blue 	<= micromatriz[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 100;
parameter RESOLUCION_Y = 100;
wire [8:0] micromatriz[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign micromatriz[0][0] = 9'b111111111;
assign micromatriz[0][1] = 9'b111111111;
assign micromatriz[0][2] = 9'b111111111;
assign micromatriz[0][3] = 9'b111111111;
assign micromatriz[0][4] = 9'b111111111;
assign micromatriz[0][5] = 9'b111111111;
assign micromatriz[0][6] = 9'b111111111;
assign micromatriz[0][7] = 9'b111111111;
assign micromatriz[0][8] = 9'b111111111;
assign micromatriz[0][9] = 9'b111111111;
assign micromatriz[0][10] = 9'b111111111;
assign micromatriz[0][11] = 9'b111111111;
assign micromatriz[0][12] = 9'b111111111;
assign micromatriz[0][13] = 9'b111111111;
assign micromatriz[0][14] = 9'b111111111;
assign micromatriz[0][15] = 9'b111111111;
assign micromatriz[0][16] = 9'b111111111;
assign micromatriz[0][17] = 9'b111111111;
assign micromatriz[0][18] = 9'b111111111;
assign micromatriz[0][19] = 9'b111111111;
assign micromatriz[0][20] = 9'b111111111;
assign micromatriz[0][21] = 9'b111111111;
assign micromatriz[0][22] = 9'b111111111;
assign micromatriz[0][23] = 9'b111111111;
assign micromatriz[0][24] = 9'b111111111;
assign micromatriz[0][25] = 9'b111111111;
assign micromatriz[0][26] = 9'b111111111;
assign micromatriz[0][27] = 9'b111111111;
assign micromatriz[0][28] = 9'b111111111;
assign micromatriz[0][29] = 9'b111111111;
assign micromatriz[0][30] = 9'b111111111;
assign micromatriz[0][31] = 9'b111111111;
assign micromatriz[0][32] = 9'b111111111;
assign micromatriz[0][33] = 9'b111111111;
assign micromatriz[0][34] = 9'b111111111;
assign micromatriz[0][35] = 9'b111111111;
assign micromatriz[0][36] = 9'b111111111;
assign micromatriz[0][37] = 9'b111111111;
assign micromatriz[0][38] = 9'b111111111;
assign micromatriz[0][39] = 9'b111111111;
assign micromatriz[0][40] = 9'b111111111;
assign micromatriz[0][41] = 9'b111111111;
assign micromatriz[0][42] = 9'b111111111;
assign micromatriz[0][43] = 9'b111111111;
assign micromatriz[0][44] = 9'b111111111;
assign micromatriz[0][45] = 9'b111111111;
assign micromatriz[0][46] = 9'b111111111;
assign micromatriz[0][47] = 9'b111111111;
assign micromatriz[0][48] = 9'b111111111;
assign micromatriz[0][49] = 9'b111111111;
assign micromatriz[0][50] = 9'b111111111;
assign micromatriz[0][51] = 9'b111111111;
assign micromatriz[0][52] = 9'b111111111;
assign micromatriz[0][53] = 9'b111111111;
assign micromatriz[0][54] = 9'b111111111;
assign micromatriz[0][55] = 9'b111111111;
assign micromatriz[0][56] = 9'b111111111;
assign micromatriz[0][57] = 9'b111111111;
assign micromatriz[0][58] = 9'b111111111;
assign micromatriz[0][59] = 9'b111111111;
assign micromatriz[0][60] = 9'b111111111;
assign micromatriz[0][61] = 9'b111111111;
assign micromatriz[0][62] = 9'b111111111;
assign micromatriz[0][63] = 9'b111111111;
assign micromatriz[0][64] = 9'b111111111;
assign micromatriz[0][65] = 9'b111111111;
assign micromatriz[0][66] = 9'b111111111;
assign micromatriz[0][67] = 9'b111111111;
assign micromatriz[0][68] = 9'b111111111;
assign micromatriz[0][69] = 9'b111111111;
assign micromatriz[0][70] = 9'b111111111;
assign micromatriz[0][71] = 9'b111111111;
assign micromatriz[0][72] = 9'b111111111;
assign micromatriz[0][73] = 9'b111111111;
assign micromatriz[0][74] = 9'b111111111;
assign micromatriz[0][75] = 9'b111111111;
assign micromatriz[0][76] = 9'b111111111;
assign micromatriz[0][77] = 9'b111111111;
assign micromatriz[0][78] = 9'b111111111;
assign micromatriz[0][79] = 9'b111111111;
assign micromatriz[0][80] = 9'b111111111;
assign micromatriz[0][81] = 9'b111111111;
assign micromatriz[0][82] = 9'b111111111;
assign micromatriz[0][83] = 9'b111111111;
assign micromatriz[0][84] = 9'b111111111;
assign micromatriz[0][85] = 9'b111111111;
assign micromatriz[0][86] = 9'b111111111;
assign micromatriz[0][87] = 9'b111111111;
assign micromatriz[0][88] = 9'b111111111;
assign micromatriz[0][89] = 9'b111111111;
assign micromatriz[0][90] = 9'b111111111;
assign micromatriz[0][91] = 9'b111111111;
assign micromatriz[0][92] = 9'b111111111;
assign micromatriz[0][93] = 9'b111111111;
assign micromatriz[0][94] = 9'b111111111;
assign micromatriz[0][95] = 9'b111111111;
assign micromatriz[0][96] = 9'b111111111;
assign micromatriz[0][97] = 9'b111111111;
assign micromatriz[0][98] = 9'b111111111;
assign micromatriz[0][99] = 9'b111111111;
assign micromatriz[1][0] = 9'b111111111;
assign micromatriz[1][1] = 9'b111111111;
assign micromatriz[1][2] = 9'b111111111;
assign micromatriz[1][3] = 9'b111111111;
assign micromatriz[1][4] = 9'b111111111;
assign micromatriz[1][5] = 9'b111111111;
assign micromatriz[1][6] = 9'b111111111;
assign micromatriz[1][7] = 9'b111111111;
assign micromatriz[1][8] = 9'b111111111;
assign micromatriz[1][9] = 9'b111111111;
assign micromatriz[1][10] = 9'b111111111;
assign micromatriz[1][11] = 9'b111111111;
assign micromatriz[1][12] = 9'b111111111;
assign micromatriz[1][13] = 9'b111111111;
assign micromatriz[1][14] = 9'b111111111;
assign micromatriz[1][15] = 9'b111111111;
assign micromatriz[1][16] = 9'b111111111;
assign micromatriz[1][17] = 9'b111111111;
assign micromatriz[1][18] = 9'b111111111;
assign micromatriz[1][19] = 9'b111111111;
assign micromatriz[1][20] = 9'b111111111;
assign micromatriz[1][21] = 9'b111111111;
assign micromatriz[1][22] = 9'b111111111;
assign micromatriz[1][23] = 9'b111111111;
assign micromatriz[1][24] = 9'b111111111;
assign micromatriz[1][25] = 9'b111111111;
assign micromatriz[1][26] = 9'b111111111;
assign micromatriz[1][27] = 9'b111111111;
assign micromatriz[1][28] = 9'b111111111;
assign micromatriz[1][29] = 9'b111111111;
assign micromatriz[1][30] = 9'b111111111;
assign micromatriz[1][31] = 9'b111111111;
assign micromatriz[1][32] = 9'b111111111;
assign micromatriz[1][33] = 9'b111111111;
assign micromatriz[1][34] = 9'b111111111;
assign micromatriz[1][35] = 9'b111111111;
assign micromatriz[1][36] = 9'b111111111;
assign micromatriz[1][37] = 9'b111111111;
assign micromatriz[1][38] = 9'b111111111;
assign micromatriz[1][39] = 9'b111111111;
assign micromatriz[1][40] = 9'b111111111;
assign micromatriz[1][41] = 9'b111111111;
assign micromatriz[1][42] = 9'b111111111;
assign micromatriz[1][43] = 9'b111111111;
assign micromatriz[1][44] = 9'b111111111;
assign micromatriz[1][45] = 9'b111111111;
assign micromatriz[1][46] = 9'b111111111;
assign micromatriz[1][47] = 9'b111111111;
assign micromatriz[1][48] = 9'b111111111;
assign micromatriz[1][49] = 9'b111111111;
assign micromatriz[1][50] = 9'b111111111;
assign micromatriz[1][51] = 9'b111111111;
assign micromatriz[1][52] = 9'b111111111;
assign micromatriz[1][53] = 9'b111111111;
assign micromatriz[1][54] = 9'b111111111;
assign micromatriz[1][55] = 9'b111111111;
assign micromatriz[1][56] = 9'b111111111;
assign micromatriz[1][57] = 9'b111111111;
assign micromatriz[1][58] = 9'b111111111;
assign micromatriz[1][59] = 9'b111111111;
assign micromatriz[1][60] = 9'b111111111;
assign micromatriz[1][61] = 9'b111111111;
assign micromatriz[1][62] = 9'b111111111;
assign micromatriz[1][63] = 9'b111111111;
assign micromatriz[1][64] = 9'b111111111;
assign micromatriz[1][65] = 9'b111111111;
assign micromatriz[1][66] = 9'b111111111;
assign micromatriz[1][67] = 9'b111111111;
assign micromatriz[1][68] = 9'b111111111;
assign micromatriz[1][69] = 9'b111111111;
assign micromatriz[1][70] = 9'b111111111;
assign micromatriz[1][71] = 9'b111111111;
assign micromatriz[1][72] = 9'b111111111;
assign micromatriz[1][73] = 9'b111111111;
assign micromatriz[1][74] = 9'b111111111;
assign micromatriz[1][75] = 9'b111111111;
assign micromatriz[1][76] = 9'b111111111;
assign micromatriz[1][77] = 9'b111111111;
assign micromatriz[1][78] = 9'b111111111;
assign micromatriz[1][79] = 9'b111111111;
assign micromatriz[1][80] = 9'b111111111;
assign micromatriz[1][81] = 9'b111111111;
assign micromatriz[1][82] = 9'b111111111;
assign micromatriz[1][83] = 9'b111111111;
assign micromatriz[1][84] = 9'b111111111;
assign micromatriz[1][85] = 9'b111111111;
assign micromatriz[1][86] = 9'b111111111;
assign micromatriz[1][87] = 9'b111111111;
assign micromatriz[1][88] = 9'b111111111;
assign micromatriz[1][89] = 9'b111111111;
assign micromatriz[1][90] = 9'b111111111;
assign micromatriz[1][91] = 9'b111111111;
assign micromatriz[1][92] = 9'b111111111;
assign micromatriz[1][93] = 9'b111111111;
assign micromatriz[1][94] = 9'b111111111;
assign micromatriz[1][95] = 9'b111111111;
assign micromatriz[1][96] = 9'b111111111;
assign micromatriz[1][97] = 9'b111111111;
assign micromatriz[1][98] = 9'b111111111;
assign micromatriz[1][99] = 9'b111111111;
assign micromatriz[2][0] = 9'b111111111;
assign micromatriz[2][1] = 9'b111111111;
assign micromatriz[2][2] = 9'b111111111;
assign micromatriz[2][3] = 9'b111111111;
assign micromatriz[2][4] = 9'b111111111;
assign micromatriz[2][5] = 9'b111111111;
assign micromatriz[2][6] = 9'b111111111;
assign micromatriz[2][7] = 9'b111111111;
assign micromatriz[2][8] = 9'b111111111;
assign micromatriz[2][9] = 9'b111111111;
assign micromatriz[2][10] = 9'b111111111;
assign micromatriz[2][11] = 9'b111111111;
assign micromatriz[2][12] = 9'b111111111;
assign micromatriz[2][13] = 9'b111111111;
assign micromatriz[2][14] = 9'b111111111;
assign micromatriz[2][15] = 9'b111111111;
assign micromatriz[2][16] = 9'b111111111;
assign micromatriz[2][17] = 9'b111111111;
assign micromatriz[2][18] = 9'b111111111;
assign micromatriz[2][19] = 9'b111111111;
assign micromatriz[2][20] = 9'b111111111;
assign micromatriz[2][21] = 9'b111111111;
assign micromatriz[2][22] = 9'b111111111;
assign micromatriz[2][23] = 9'b111111111;
assign micromatriz[2][24] = 9'b111111111;
assign micromatriz[2][25] = 9'b111111111;
assign micromatriz[2][26] = 9'b111111111;
assign micromatriz[2][27] = 9'b111111111;
assign micromatriz[2][28] = 9'b111111111;
assign micromatriz[2][29] = 9'b111111111;
assign micromatriz[2][30] = 9'b111111111;
assign micromatriz[2][31] = 9'b111111111;
assign micromatriz[2][32] = 9'b111111111;
assign micromatriz[2][33] = 9'b111111111;
assign micromatriz[2][34] = 9'b111111111;
assign micromatriz[2][35] = 9'b111111111;
assign micromatriz[2][36] = 9'b111111111;
assign micromatriz[2][37] = 9'b111111111;
assign micromatriz[2][38] = 9'b111111111;
assign micromatriz[2][39] = 9'b111111111;
assign micromatriz[2][40] = 9'b111111111;
assign micromatriz[2][41] = 9'b111111111;
assign micromatriz[2][42] = 9'b111111111;
assign micromatriz[2][43] = 9'b111111111;
assign micromatriz[2][44] = 9'b111111111;
assign micromatriz[2][45] = 9'b111111111;
assign micromatriz[2][46] = 9'b111111111;
assign micromatriz[2][47] = 9'b111111111;
assign micromatriz[2][48] = 9'b111111111;
assign micromatriz[2][49] = 9'b111111111;
assign micromatriz[2][50] = 9'b111111111;
assign micromatriz[2][51] = 9'b111111111;
assign micromatriz[2][52] = 9'b111111111;
assign micromatriz[2][53] = 9'b111111111;
assign micromatriz[2][54] = 9'b111111111;
assign micromatriz[2][55] = 9'b111111111;
assign micromatriz[2][56] = 9'b111111111;
assign micromatriz[2][57] = 9'b111111111;
assign micromatriz[2][58] = 9'b111111111;
assign micromatriz[2][59] = 9'b111111111;
assign micromatriz[2][60] = 9'b111111111;
assign micromatriz[2][61] = 9'b111111111;
assign micromatriz[2][62] = 9'b111111111;
assign micromatriz[2][63] = 9'b111111111;
assign micromatriz[2][64] = 9'b111111111;
assign micromatriz[2][65] = 9'b111111111;
assign micromatriz[2][66] = 9'b111111111;
assign micromatriz[2][67] = 9'b111111111;
assign micromatriz[2][68] = 9'b111111111;
assign micromatriz[2][69] = 9'b111111111;
assign micromatriz[2][70] = 9'b111111111;
assign micromatriz[2][71] = 9'b111111111;
assign micromatriz[2][72] = 9'b111111111;
assign micromatriz[2][73] = 9'b111111111;
assign micromatriz[2][74] = 9'b111111111;
assign micromatriz[2][75] = 9'b111111111;
assign micromatriz[2][76] = 9'b111111111;
assign micromatriz[2][77] = 9'b111111111;
assign micromatriz[2][78] = 9'b111111111;
assign micromatriz[2][79] = 9'b111111111;
assign micromatriz[2][80] = 9'b111111111;
assign micromatriz[2][81] = 9'b111111111;
assign micromatriz[2][82] = 9'b111111111;
assign micromatriz[2][83] = 9'b111111111;
assign micromatriz[2][84] = 9'b111111111;
assign micromatriz[2][85] = 9'b111111111;
assign micromatriz[2][86] = 9'b111111111;
assign micromatriz[2][87] = 9'b111111111;
assign micromatriz[2][88] = 9'b111111111;
assign micromatriz[2][89] = 9'b111111111;
assign micromatriz[2][90] = 9'b111111111;
assign micromatriz[2][91] = 9'b111111111;
assign micromatriz[2][92] = 9'b111111111;
assign micromatriz[2][93] = 9'b111111111;
assign micromatriz[2][94] = 9'b111111111;
assign micromatriz[2][95] = 9'b111111111;
assign micromatriz[2][96] = 9'b111111111;
assign micromatriz[2][97] = 9'b111111111;
assign micromatriz[2][98] = 9'b111111111;
assign micromatriz[2][99] = 9'b111111111;
assign micromatriz[3][0] = 9'b111111111;
assign micromatriz[3][1] = 9'b111111111;
assign micromatriz[3][2] = 9'b111111111;
assign micromatriz[3][3] = 9'b111111111;
assign micromatriz[3][4] = 9'b111111111;
assign micromatriz[3][5] = 9'b111111111;
assign micromatriz[3][6] = 9'b111111111;
assign micromatriz[3][7] = 9'b111111111;
assign micromatriz[3][8] = 9'b111111111;
assign micromatriz[3][9] = 9'b111111111;
assign micromatriz[3][10] = 9'b111111111;
assign micromatriz[3][11] = 9'b111111111;
assign micromatriz[3][12] = 9'b111111111;
assign micromatriz[3][13] = 9'b111111111;
assign micromatriz[3][14] = 9'b111111111;
assign micromatriz[3][15] = 9'b111111111;
assign micromatriz[3][16] = 9'b111111111;
assign micromatriz[3][17] = 9'b111111111;
assign micromatriz[3][18] = 9'b111111111;
assign micromatriz[3][19] = 9'b111111111;
assign micromatriz[3][20] = 9'b111111111;
assign micromatriz[3][21] = 9'b111111111;
assign micromatriz[3][22] = 9'b111111111;
assign micromatriz[3][23] = 9'b111111111;
assign micromatriz[3][24] = 9'b111111111;
assign micromatriz[3][25] = 9'b111111111;
assign micromatriz[3][26] = 9'b111111111;
assign micromatriz[3][27] = 9'b111111111;
assign micromatriz[3][28] = 9'b111111111;
assign micromatriz[3][29] = 9'b111111111;
assign micromatriz[3][30] = 9'b111111111;
assign micromatriz[3][31] = 9'b111111111;
assign micromatriz[3][32] = 9'b111111111;
assign micromatriz[3][33] = 9'b111111111;
assign micromatriz[3][34] = 9'b111111111;
assign micromatriz[3][35] = 9'b111111111;
assign micromatriz[3][36] = 9'b111111111;
assign micromatriz[3][37] = 9'b111111111;
assign micromatriz[3][38] = 9'b111111111;
assign micromatriz[3][39] = 9'b111111111;
assign micromatriz[3][40] = 9'b111111111;
assign micromatriz[3][41] = 9'b111111111;
assign micromatriz[3][42] = 9'b111111111;
assign micromatriz[3][43] = 9'b111111111;
assign micromatriz[3][44] = 9'b111111111;
assign micromatriz[3][45] = 9'b111111111;
assign micromatriz[3][46] = 9'b111111111;
assign micromatriz[3][47] = 9'b111111111;
assign micromatriz[3][48] = 9'b111111111;
assign micromatriz[3][49] = 9'b111111111;
assign micromatriz[3][50] = 9'b111111111;
assign micromatriz[3][51] = 9'b111111111;
assign micromatriz[3][52] = 9'b111111111;
assign micromatriz[3][53] = 9'b111111111;
assign micromatriz[3][54] = 9'b111111111;
assign micromatriz[3][55] = 9'b111111111;
assign micromatriz[3][56] = 9'b111111111;
assign micromatriz[3][57] = 9'b111111111;
assign micromatriz[3][58] = 9'b111111111;
assign micromatriz[3][59] = 9'b111111111;
assign micromatriz[3][60] = 9'b111111111;
assign micromatriz[3][61] = 9'b111111111;
assign micromatriz[3][62] = 9'b111111111;
assign micromatriz[3][63] = 9'b111111111;
assign micromatriz[3][64] = 9'b111111111;
assign micromatriz[3][65] = 9'b111111111;
assign micromatriz[3][66] = 9'b111111111;
assign micromatriz[3][67] = 9'b111111111;
assign micromatriz[3][68] = 9'b111111111;
assign micromatriz[3][69] = 9'b111111111;
assign micromatriz[3][70] = 9'b111111111;
assign micromatriz[3][71] = 9'b111111111;
assign micromatriz[3][72] = 9'b111111111;
assign micromatriz[3][73] = 9'b111111111;
assign micromatriz[3][74] = 9'b111111111;
assign micromatriz[3][75] = 9'b111111111;
assign micromatriz[3][76] = 9'b111111111;
assign micromatriz[3][77] = 9'b111111111;
assign micromatriz[3][78] = 9'b111111111;
assign micromatriz[3][79] = 9'b111111111;
assign micromatriz[3][80] = 9'b111111111;
assign micromatriz[3][81] = 9'b111111111;
assign micromatriz[3][82] = 9'b111111111;
assign micromatriz[3][83] = 9'b111111111;
assign micromatriz[3][84] = 9'b111111111;
assign micromatriz[3][85] = 9'b111111111;
assign micromatriz[3][86] = 9'b111111111;
assign micromatriz[3][87] = 9'b111111111;
assign micromatriz[3][88] = 9'b111111111;
assign micromatriz[3][89] = 9'b111111111;
assign micromatriz[3][90] = 9'b111111111;
assign micromatriz[3][91] = 9'b111111111;
assign micromatriz[3][92] = 9'b111111111;
assign micromatriz[3][93] = 9'b111111111;
assign micromatriz[3][94] = 9'b111111111;
assign micromatriz[3][95] = 9'b111111111;
assign micromatriz[3][96] = 9'b111111111;
assign micromatriz[3][97] = 9'b111111111;
assign micromatriz[3][98] = 9'b111111111;
assign micromatriz[3][99] = 9'b111111111;
assign micromatriz[4][0] = 9'b111111111;
assign micromatriz[4][1] = 9'b111111111;
assign micromatriz[4][2] = 9'b111111111;
assign micromatriz[4][3] = 9'b111111111;
assign micromatriz[4][4] = 9'b111111111;
assign micromatriz[4][5] = 9'b111111111;
assign micromatriz[4][6] = 9'b111111111;
assign micromatriz[4][7] = 9'b111111111;
assign micromatriz[4][8] = 9'b111111111;
assign micromatriz[4][9] = 9'b111111111;
assign micromatriz[4][10] = 9'b111111111;
assign micromatriz[4][11] = 9'b111111111;
assign micromatriz[4][12] = 9'b111111111;
assign micromatriz[4][13] = 9'b111111111;
assign micromatriz[4][14] = 9'b111111111;
assign micromatriz[4][15] = 9'b111111111;
assign micromatriz[4][16] = 9'b111111111;
assign micromatriz[4][17] = 9'b111111111;
assign micromatriz[4][18] = 9'b111111111;
assign micromatriz[4][19] = 9'b111111111;
assign micromatriz[4][20] = 9'b111111111;
assign micromatriz[4][21] = 9'b111111111;
assign micromatriz[4][22] = 9'b111111111;
assign micromatriz[4][23] = 9'b111111111;
assign micromatriz[4][24] = 9'b111111111;
assign micromatriz[4][25] = 9'b111111111;
assign micromatriz[4][26] = 9'b111111111;
assign micromatriz[4][27] = 9'b111111111;
assign micromatriz[4][28] = 9'b111111111;
assign micromatriz[4][29] = 9'b111111111;
assign micromatriz[4][30] = 9'b111111111;
assign micromatriz[4][31] = 9'b111111111;
assign micromatriz[4][32] = 9'b111111111;
assign micromatriz[4][33] = 9'b111111111;
assign micromatriz[4][34] = 9'b111111111;
assign micromatriz[4][35] = 9'b111111111;
assign micromatriz[4][36] = 9'b111111111;
assign micromatriz[4][37] = 9'b111111111;
assign micromatriz[4][38] = 9'b111111111;
assign micromatriz[4][39] = 9'b111111111;
assign micromatriz[4][40] = 9'b111111111;
assign micromatriz[4][41] = 9'b111111111;
assign micromatriz[4][42] = 9'b111111111;
assign micromatriz[4][43] = 9'b111111111;
assign micromatriz[4][44] = 9'b111111111;
assign micromatriz[4][45] = 9'b111111111;
assign micromatriz[4][46] = 9'b111111111;
assign micromatriz[4][47] = 9'b111111111;
assign micromatriz[4][48] = 9'b111111111;
assign micromatriz[4][49] = 9'b111111111;
assign micromatriz[4][50] = 9'b111111111;
assign micromatriz[4][51] = 9'b111111111;
assign micromatriz[4][52] = 9'b111111111;
assign micromatriz[4][53] = 9'b111111111;
assign micromatriz[4][54] = 9'b111111111;
assign micromatriz[4][55] = 9'b111111111;
assign micromatriz[4][56] = 9'b111111111;
assign micromatriz[4][57] = 9'b111111111;
assign micromatriz[4][58] = 9'b111111111;
assign micromatriz[4][59] = 9'b111111111;
assign micromatriz[4][60] = 9'b111111111;
assign micromatriz[4][61] = 9'b111111111;
assign micromatriz[4][62] = 9'b111111111;
assign micromatriz[4][63] = 9'b111111111;
assign micromatriz[4][64] = 9'b111111111;
assign micromatriz[4][65] = 9'b111111111;
assign micromatriz[4][66] = 9'b111111111;
assign micromatriz[4][67] = 9'b111111111;
assign micromatriz[4][68] = 9'b111111111;
assign micromatriz[4][69] = 9'b111111111;
assign micromatriz[4][70] = 9'b111111111;
assign micromatriz[4][71] = 9'b111111111;
assign micromatriz[4][72] = 9'b111111111;
assign micromatriz[4][73] = 9'b111111111;
assign micromatriz[4][74] = 9'b111111111;
assign micromatriz[4][75] = 9'b111111111;
assign micromatriz[4][76] = 9'b111111111;
assign micromatriz[4][77] = 9'b111111111;
assign micromatriz[4][78] = 9'b111111111;
assign micromatriz[4][79] = 9'b111111111;
assign micromatriz[4][80] = 9'b111111111;
assign micromatriz[4][81] = 9'b111111111;
assign micromatriz[4][82] = 9'b111111111;
assign micromatriz[4][83] = 9'b111111111;
assign micromatriz[4][84] = 9'b111111111;
assign micromatriz[4][85] = 9'b111111111;
assign micromatriz[4][86] = 9'b111111111;
assign micromatriz[4][87] = 9'b111111111;
assign micromatriz[4][88] = 9'b111111111;
assign micromatriz[4][89] = 9'b111111111;
assign micromatriz[4][90] = 9'b111111111;
assign micromatriz[4][91] = 9'b111111111;
assign micromatriz[4][92] = 9'b111111111;
assign micromatriz[4][93] = 9'b111111111;
assign micromatriz[4][94] = 9'b111111111;
assign micromatriz[4][95] = 9'b111111111;
assign micromatriz[4][96] = 9'b111111111;
assign micromatriz[4][97] = 9'b111111111;
assign micromatriz[4][98] = 9'b111111111;
assign micromatriz[4][99] = 9'b111111111;
assign micromatriz[5][0] = 9'b111111111;
assign micromatriz[5][1] = 9'b111111111;
assign micromatriz[5][2] = 9'b111111111;
assign micromatriz[5][3] = 9'b111111111;
assign micromatriz[5][4] = 9'b111111111;
assign micromatriz[5][5] = 9'b111111111;
assign micromatriz[5][6] = 9'b111111111;
assign micromatriz[5][7] = 9'b111111111;
assign micromatriz[5][8] = 9'b111111111;
assign micromatriz[5][9] = 9'b111111111;
assign micromatriz[5][10] = 9'b111111111;
assign micromatriz[5][11] = 9'b111111111;
assign micromatriz[5][12] = 9'b111111111;
assign micromatriz[5][13] = 9'b111111111;
assign micromatriz[5][14] = 9'b111111111;
assign micromatriz[5][15] = 9'b111111111;
assign micromatriz[5][16] = 9'b111111111;
assign micromatriz[5][17] = 9'b111111111;
assign micromatriz[5][18] = 9'b111111111;
assign micromatriz[5][19] = 9'b111111111;
assign micromatriz[5][20] = 9'b111111111;
assign micromatriz[5][21] = 9'b111111111;
assign micromatriz[5][22] = 9'b111111111;
assign micromatriz[5][23] = 9'b111111111;
assign micromatriz[5][24] = 9'b111111111;
assign micromatriz[5][25] = 9'b111111111;
assign micromatriz[5][26] = 9'b111111111;
assign micromatriz[5][27] = 9'b111111111;
assign micromatriz[5][28] = 9'b111111111;
assign micromatriz[5][29] = 9'b111111111;
assign micromatriz[5][30] = 9'b111111111;
assign micromatriz[5][31] = 9'b111111111;
assign micromatriz[5][32] = 9'b111111111;
assign micromatriz[5][33] = 9'b111111111;
assign micromatriz[5][34] = 9'b111111111;
assign micromatriz[5][35] = 9'b111111111;
assign micromatriz[5][36] = 9'b111111111;
assign micromatriz[5][37] = 9'b111111111;
assign micromatriz[5][38] = 9'b111111111;
assign micromatriz[5][39] = 9'b111111111;
assign micromatriz[5][40] = 9'b111111111;
assign micromatriz[5][41] = 9'b111111111;
assign micromatriz[5][42] = 9'b111111111;
assign micromatriz[5][43] = 9'b111111111;
assign micromatriz[5][44] = 9'b111111111;
assign micromatriz[5][45] = 9'b111111111;
assign micromatriz[5][46] = 9'b111111111;
assign micromatriz[5][47] = 9'b111111111;
assign micromatriz[5][48] = 9'b111111111;
assign micromatriz[5][49] = 9'b111111111;
assign micromatriz[5][50] = 9'b111111111;
assign micromatriz[5][51] = 9'b111111111;
assign micromatriz[5][52] = 9'b111111111;
assign micromatriz[5][53] = 9'b111111111;
assign micromatriz[5][54] = 9'b111111111;
assign micromatriz[5][55] = 9'b111111111;
assign micromatriz[5][56] = 9'b111111111;
assign micromatriz[5][57] = 9'b111111111;
assign micromatriz[5][58] = 9'b111111111;
assign micromatriz[5][59] = 9'b111111111;
assign micromatriz[5][60] = 9'b111111111;
assign micromatriz[5][61] = 9'b111111111;
assign micromatriz[5][62] = 9'b111111111;
assign micromatriz[5][63] = 9'b111111111;
assign micromatriz[5][64] = 9'b111111111;
assign micromatriz[5][65] = 9'b111111111;
assign micromatriz[5][66] = 9'b111111111;
assign micromatriz[5][67] = 9'b111111111;
assign micromatriz[5][68] = 9'b111111111;
assign micromatriz[5][69] = 9'b111111111;
assign micromatriz[5][70] = 9'b111111111;
assign micromatriz[5][71] = 9'b111111111;
assign micromatriz[5][72] = 9'b111111111;
assign micromatriz[5][73] = 9'b111111111;
assign micromatriz[5][74] = 9'b111111111;
assign micromatriz[5][75] = 9'b111111111;
assign micromatriz[5][76] = 9'b111111111;
assign micromatriz[5][77] = 9'b111111111;
assign micromatriz[5][78] = 9'b111111111;
assign micromatriz[5][79] = 9'b111111111;
assign micromatriz[5][80] = 9'b111111111;
assign micromatriz[5][81] = 9'b111111111;
assign micromatriz[5][82] = 9'b111111111;
assign micromatriz[5][83] = 9'b111111111;
assign micromatriz[5][84] = 9'b111111111;
assign micromatriz[5][85] = 9'b111111111;
assign micromatriz[5][86] = 9'b111111111;
assign micromatriz[5][87] = 9'b111111111;
assign micromatriz[5][88] = 9'b111111111;
assign micromatriz[5][89] = 9'b111111111;
assign micromatriz[5][90] = 9'b111111111;
assign micromatriz[5][91] = 9'b111111111;
assign micromatriz[5][92] = 9'b111111111;
assign micromatriz[5][93] = 9'b111111111;
assign micromatriz[5][94] = 9'b111111111;
assign micromatriz[5][95] = 9'b111111111;
assign micromatriz[5][96] = 9'b111111111;
assign micromatriz[5][97] = 9'b111111111;
assign micromatriz[5][98] = 9'b111111111;
assign micromatriz[5][99] = 9'b111111111;
assign micromatriz[6][0] = 9'b111111111;
assign micromatriz[6][1] = 9'b111111111;
assign micromatriz[6][2] = 9'b111111111;
assign micromatriz[6][3] = 9'b111111111;
assign micromatriz[6][4] = 9'b111111111;
assign micromatriz[6][5] = 9'b111111111;
assign micromatriz[6][6] = 9'b111111111;
assign micromatriz[6][7] = 9'b111111111;
assign micromatriz[6][8] = 9'b111111111;
assign micromatriz[6][9] = 9'b111111111;
assign micromatriz[6][10] = 9'b111111111;
assign micromatriz[6][11] = 9'b111111111;
assign micromatriz[6][12] = 9'b111111111;
assign micromatriz[6][13] = 9'b111111111;
assign micromatriz[6][14] = 9'b111111111;
assign micromatriz[6][15] = 9'b111111111;
assign micromatriz[6][16] = 9'b111111111;
assign micromatriz[6][17] = 9'b111111111;
assign micromatriz[6][18] = 9'b111111111;
assign micromatriz[6][19] = 9'b111111111;
assign micromatriz[6][20] = 9'b111111111;
assign micromatriz[6][21] = 9'b111111111;
assign micromatriz[6][22] = 9'b111111111;
assign micromatriz[6][23] = 9'b111111111;
assign micromatriz[6][24] = 9'b111111111;
assign micromatriz[6][25] = 9'b111111111;
assign micromatriz[6][26] = 9'b111111111;
assign micromatriz[6][27] = 9'b111111111;
assign micromatriz[6][28] = 9'b111111111;
assign micromatriz[6][29] = 9'b111111111;
assign micromatriz[6][30] = 9'b111111111;
assign micromatriz[6][31] = 9'b111111111;
assign micromatriz[6][32] = 9'b111111111;
assign micromatriz[6][33] = 9'b111111111;
assign micromatriz[6][34] = 9'b111111111;
assign micromatriz[6][35] = 9'b111111111;
assign micromatriz[6][36] = 9'b111111111;
assign micromatriz[6][37] = 9'b111111111;
assign micromatriz[6][38] = 9'b111111111;
assign micromatriz[6][39] = 9'b111111111;
assign micromatriz[6][40] = 9'b111111111;
assign micromatriz[6][41] = 9'b111111111;
assign micromatriz[6][42] = 9'b111111111;
assign micromatriz[6][43] = 9'b111111111;
assign micromatriz[6][44] = 9'b111111111;
assign micromatriz[6][45] = 9'b111111111;
assign micromatriz[6][46] = 9'b111111111;
assign micromatriz[6][47] = 9'b111111111;
assign micromatriz[6][48] = 9'b111111111;
assign micromatriz[6][49] = 9'b111111111;
assign micromatriz[6][50] = 9'b111111111;
assign micromatriz[6][51] = 9'b111111111;
assign micromatriz[6][52] = 9'b111111111;
assign micromatriz[6][53] = 9'b111111111;
assign micromatriz[6][54] = 9'b111111111;
assign micromatriz[6][55] = 9'b111111111;
assign micromatriz[6][56] = 9'b111111111;
assign micromatriz[6][57] = 9'b111111111;
assign micromatriz[6][58] = 9'b111111111;
assign micromatriz[6][59] = 9'b111111111;
assign micromatriz[6][60] = 9'b111111111;
assign micromatriz[6][61] = 9'b111111111;
assign micromatriz[6][62] = 9'b111111111;
assign micromatriz[6][63] = 9'b111111111;
assign micromatriz[6][64] = 9'b111111111;
assign micromatriz[6][65] = 9'b111111111;
assign micromatriz[6][66] = 9'b111111111;
assign micromatriz[6][67] = 9'b111111111;
assign micromatriz[6][68] = 9'b111111111;
assign micromatriz[6][69] = 9'b111111111;
assign micromatriz[6][70] = 9'b111111111;
assign micromatriz[6][71] = 9'b111111111;
assign micromatriz[6][72] = 9'b111111111;
assign micromatriz[6][73] = 9'b111111111;
assign micromatriz[6][74] = 9'b111111111;
assign micromatriz[6][75] = 9'b111111111;
assign micromatriz[6][76] = 9'b111111111;
assign micromatriz[6][77] = 9'b111111111;
assign micromatriz[6][78] = 9'b111111111;
assign micromatriz[6][79] = 9'b111111111;
assign micromatriz[6][80] = 9'b111111111;
assign micromatriz[6][81] = 9'b111111111;
assign micromatriz[6][82] = 9'b111111111;
assign micromatriz[6][83] = 9'b111111111;
assign micromatriz[6][84] = 9'b111111111;
assign micromatriz[6][85] = 9'b111111111;
assign micromatriz[6][86] = 9'b111111111;
assign micromatriz[6][87] = 9'b111111111;
assign micromatriz[6][88] = 9'b111111111;
assign micromatriz[6][89] = 9'b111111111;
assign micromatriz[6][90] = 9'b111111111;
assign micromatriz[6][91] = 9'b111111111;
assign micromatriz[6][92] = 9'b111111111;
assign micromatriz[6][93] = 9'b111111111;
assign micromatriz[6][94] = 9'b111111111;
assign micromatriz[6][95] = 9'b111111111;
assign micromatriz[6][96] = 9'b111111111;
assign micromatriz[6][97] = 9'b111111111;
assign micromatriz[6][98] = 9'b111111111;
assign micromatriz[6][99] = 9'b111111111;
assign micromatriz[7][0] = 9'b111111111;
assign micromatriz[7][1] = 9'b111111111;
assign micromatriz[7][2] = 9'b111111111;
assign micromatriz[7][3] = 9'b111111111;
assign micromatriz[7][4] = 9'b111111111;
assign micromatriz[7][5] = 9'b111111111;
assign micromatriz[7][6] = 9'b111111111;
assign micromatriz[7][7] = 9'b111111111;
assign micromatriz[7][8] = 9'b111111111;
assign micromatriz[7][9] = 9'b111111111;
assign micromatriz[7][10] = 9'b111111111;
assign micromatriz[7][11] = 9'b111111111;
assign micromatriz[7][12] = 9'b111111111;
assign micromatriz[7][13] = 9'b111111111;
assign micromatriz[7][14] = 9'b111111111;
assign micromatriz[7][15] = 9'b111111111;
assign micromatriz[7][16] = 9'b111111111;
assign micromatriz[7][17] = 9'b111111111;
assign micromatriz[7][18] = 9'b111111111;
assign micromatriz[7][19] = 9'b111111111;
assign micromatriz[7][20] = 9'b111111111;
assign micromatriz[7][21] = 9'b111111111;
assign micromatriz[7][22] = 9'b111111111;
assign micromatriz[7][23] = 9'b111111111;
assign micromatriz[7][24] = 9'b111111111;
assign micromatriz[7][25] = 9'b111111111;
assign micromatriz[7][26] = 9'b111111111;
assign micromatriz[7][27] = 9'b111111111;
assign micromatriz[7][28] = 9'b111111111;
assign micromatriz[7][29] = 9'b111111111;
assign micromatriz[7][30] = 9'b111111111;
assign micromatriz[7][31] = 9'b111111111;
assign micromatriz[7][32] = 9'b111111111;
assign micromatriz[7][33] = 9'b111111111;
assign micromatriz[7][34] = 9'b111111111;
assign micromatriz[7][35] = 9'b111111111;
assign micromatriz[7][36] = 9'b111111111;
assign micromatriz[7][37] = 9'b111111111;
assign micromatriz[7][38] = 9'b111111111;
assign micromatriz[7][39] = 9'b111111111;
assign micromatriz[7][40] = 9'b111111111;
assign micromatriz[7][41] = 9'b111111111;
assign micromatriz[7][42] = 9'b111111111;
assign micromatriz[7][43] = 9'b111111111;
assign micromatriz[7][44] = 9'b111111111;
assign micromatriz[7][45] = 9'b111111111;
assign micromatriz[7][46] = 9'b111111111;
assign micromatriz[7][47] = 9'b111111111;
assign micromatriz[7][48] = 9'b111111111;
assign micromatriz[7][49] = 9'b111111111;
assign micromatriz[7][50] = 9'b111111111;
assign micromatriz[7][51] = 9'b111111111;
assign micromatriz[7][52] = 9'b111111111;
assign micromatriz[7][53] = 9'b111111111;
assign micromatriz[7][54] = 9'b111111111;
assign micromatriz[7][55] = 9'b111111111;
assign micromatriz[7][56] = 9'b111111111;
assign micromatriz[7][57] = 9'b111111111;
assign micromatriz[7][58] = 9'b111111111;
assign micromatriz[7][59] = 9'b111111111;
assign micromatriz[7][60] = 9'b111111111;
assign micromatriz[7][61] = 9'b111111111;
assign micromatriz[7][62] = 9'b111111111;
assign micromatriz[7][63] = 9'b111111111;
assign micromatriz[7][64] = 9'b111111111;
assign micromatriz[7][65] = 9'b111111111;
assign micromatriz[7][66] = 9'b111111111;
assign micromatriz[7][67] = 9'b111111111;
assign micromatriz[7][68] = 9'b111111111;
assign micromatriz[7][69] = 9'b111111111;
assign micromatriz[7][70] = 9'b111111111;
assign micromatriz[7][71] = 9'b111111111;
assign micromatriz[7][72] = 9'b111111111;
assign micromatriz[7][73] = 9'b111111111;
assign micromatriz[7][74] = 9'b111111111;
assign micromatriz[7][75] = 9'b111111111;
assign micromatriz[7][76] = 9'b111111111;
assign micromatriz[7][77] = 9'b111111111;
assign micromatriz[7][78] = 9'b111111111;
assign micromatriz[7][79] = 9'b111111111;
assign micromatriz[7][80] = 9'b111111111;
assign micromatriz[7][81] = 9'b111111111;
assign micromatriz[7][82] = 9'b111111111;
assign micromatriz[7][83] = 9'b111111111;
assign micromatriz[7][84] = 9'b111111111;
assign micromatriz[7][85] = 9'b111111111;
assign micromatriz[7][86] = 9'b111111111;
assign micromatriz[7][87] = 9'b111111111;
assign micromatriz[7][88] = 9'b111111111;
assign micromatriz[7][89] = 9'b111111111;
assign micromatriz[7][90] = 9'b111111111;
assign micromatriz[7][91] = 9'b111111111;
assign micromatriz[7][92] = 9'b111111111;
assign micromatriz[7][93] = 9'b111111111;
assign micromatriz[7][94] = 9'b111111111;
assign micromatriz[7][95] = 9'b111111111;
assign micromatriz[7][96] = 9'b111111111;
assign micromatriz[7][97] = 9'b111111111;
assign micromatriz[7][98] = 9'b111111111;
assign micromatriz[7][99] = 9'b111111111;
assign micromatriz[8][0] = 9'b111111111;
assign micromatriz[8][1] = 9'b111111111;
assign micromatriz[8][2] = 9'b111111111;
assign micromatriz[8][3] = 9'b111111111;
assign micromatriz[8][4] = 9'b111111111;
assign micromatriz[8][5] = 9'b111111111;
assign micromatriz[8][6] = 9'b111111111;
assign micromatriz[8][7] = 9'b111111111;
assign micromatriz[8][8] = 9'b111111111;
assign micromatriz[8][9] = 9'b111111111;
assign micromatriz[8][10] = 9'b111111111;
assign micromatriz[8][11] = 9'b111111111;
assign micromatriz[8][12] = 9'b111111111;
assign micromatriz[8][13] = 9'b111111111;
assign micromatriz[8][14] = 9'b111111111;
assign micromatriz[8][15] = 9'b111111111;
assign micromatriz[8][16] = 9'b111111111;
assign micromatriz[8][17] = 9'b111111111;
assign micromatriz[8][18] = 9'b111111111;
assign micromatriz[8][19] = 9'b111111111;
assign micromatriz[8][20] = 9'b111111111;
assign micromatriz[8][21] = 9'b111111111;
assign micromatriz[8][22] = 9'b111111111;
assign micromatriz[8][23] = 9'b111111111;
assign micromatriz[8][24] = 9'b111111111;
assign micromatriz[8][25] = 9'b111111111;
assign micromatriz[8][26] = 9'b111111111;
assign micromatriz[8][27] = 9'b111111111;
assign micromatriz[8][28] = 9'b111111111;
assign micromatriz[8][29] = 9'b111111111;
assign micromatriz[8][30] = 9'b111111111;
assign micromatriz[8][31] = 9'b111111111;
assign micromatriz[8][32] = 9'b111111111;
assign micromatriz[8][33] = 9'b111111111;
assign micromatriz[8][34] = 9'b111111111;
assign micromatriz[8][35] = 9'b111111111;
assign micromatriz[8][36] = 9'b111111111;
assign micromatriz[8][37] = 9'b111111111;
assign micromatriz[8][38] = 9'b111111111;
assign micromatriz[8][39] = 9'b111111111;
assign micromatriz[8][40] = 9'b111111111;
assign micromatriz[8][41] = 9'b111111111;
assign micromatriz[8][42] = 9'b111111111;
assign micromatriz[8][43] = 9'b111111111;
assign micromatriz[8][44] = 9'b111111111;
assign micromatriz[8][45] = 9'b111111111;
assign micromatriz[8][46] = 9'b111111111;
assign micromatriz[8][47] = 9'b111111111;
assign micromatriz[8][48] = 9'b111111111;
assign micromatriz[8][49] = 9'b111111111;
assign micromatriz[8][50] = 9'b111111111;
assign micromatriz[8][51] = 9'b111111111;
assign micromatriz[8][52] = 9'b111111111;
assign micromatriz[8][53] = 9'b111111111;
assign micromatriz[8][54] = 9'b111111111;
assign micromatriz[8][55] = 9'b111111111;
assign micromatriz[8][56] = 9'b111111111;
assign micromatriz[8][57] = 9'b111111111;
assign micromatriz[8][58] = 9'b111111111;
assign micromatriz[8][59] = 9'b111111111;
assign micromatriz[8][60] = 9'b111111111;
assign micromatriz[8][61] = 9'b111111111;
assign micromatriz[8][62] = 9'b111111111;
assign micromatriz[8][63] = 9'b111111111;
assign micromatriz[8][64] = 9'b111111111;
assign micromatriz[8][65] = 9'b111111111;
assign micromatriz[8][66] = 9'b111111111;
assign micromatriz[8][67] = 9'b111111111;
assign micromatriz[8][68] = 9'b111111111;
assign micromatriz[8][69] = 9'b111111111;
assign micromatriz[8][70] = 9'b111111111;
assign micromatriz[8][71] = 9'b111111111;
assign micromatriz[8][72] = 9'b111111111;
assign micromatriz[8][73] = 9'b111111111;
assign micromatriz[8][74] = 9'b111111111;
assign micromatriz[8][75] = 9'b111111111;
assign micromatriz[8][76] = 9'b111111111;
assign micromatriz[8][77] = 9'b111111111;
assign micromatriz[8][78] = 9'b111111111;
assign micromatriz[8][79] = 9'b111111111;
assign micromatriz[8][80] = 9'b111111111;
assign micromatriz[8][81] = 9'b111111111;
assign micromatriz[8][82] = 9'b111111111;
assign micromatriz[8][83] = 9'b111111111;
assign micromatriz[8][84] = 9'b111111111;
assign micromatriz[8][85] = 9'b111111111;
assign micromatriz[8][86] = 9'b111111111;
assign micromatriz[8][87] = 9'b111111111;
assign micromatriz[8][88] = 9'b111111111;
assign micromatriz[8][89] = 9'b111111111;
assign micromatriz[8][90] = 9'b111111111;
assign micromatriz[8][91] = 9'b111111111;
assign micromatriz[8][92] = 9'b111111111;
assign micromatriz[8][93] = 9'b111111111;
assign micromatriz[8][94] = 9'b111111111;
assign micromatriz[8][95] = 9'b111111111;
assign micromatriz[8][96] = 9'b111111111;
assign micromatriz[8][97] = 9'b111111111;
assign micromatriz[8][98] = 9'b111111111;
assign micromatriz[8][99] = 9'b111111111;
assign micromatriz[9][0] = 9'b111111111;
assign micromatriz[9][1] = 9'b111111111;
assign micromatriz[9][2] = 9'b111111111;
assign micromatriz[9][3] = 9'b111111111;
assign micromatriz[9][4] = 9'b111111111;
assign micromatriz[9][5] = 9'b111111111;
assign micromatriz[9][6] = 9'b111111111;
assign micromatriz[9][7] = 9'b111111111;
assign micromatriz[9][8] = 9'b111111111;
assign micromatriz[9][9] = 9'b111111111;
assign micromatriz[9][10] = 9'b111111111;
assign micromatriz[9][11] = 9'b111111111;
assign micromatriz[9][12] = 9'b111111111;
assign micromatriz[9][13] = 9'b111111111;
assign micromatriz[9][14] = 9'b111111111;
assign micromatriz[9][15] = 9'b111111111;
assign micromatriz[9][16] = 9'b111111111;
assign micromatriz[9][17] = 9'b111111111;
assign micromatriz[9][18] = 9'b111111111;
assign micromatriz[9][19] = 9'b111111111;
assign micromatriz[9][20] = 9'b111111111;
assign micromatriz[9][21] = 9'b111111111;
assign micromatriz[9][22] = 9'b111111111;
assign micromatriz[9][23] = 9'b111111111;
assign micromatriz[9][24] = 9'b111111111;
assign micromatriz[9][25] = 9'b111111111;
assign micromatriz[9][26] = 9'b111111111;
assign micromatriz[9][27] = 9'b111111111;
assign micromatriz[9][28] = 9'b111111111;
assign micromatriz[9][29] = 9'b111111111;
assign micromatriz[9][30] = 9'b111111111;
assign micromatriz[9][31] = 9'b111111111;
assign micromatriz[9][32] = 9'b111111111;
assign micromatriz[9][33] = 9'b111111111;
assign micromatriz[9][34] = 9'b111111111;
assign micromatriz[9][35] = 9'b111111111;
assign micromatriz[9][36] = 9'b111111111;
assign micromatriz[9][37] = 9'b111111111;
assign micromatriz[9][38] = 9'b111111111;
assign micromatriz[9][39] = 9'b111111111;
assign micromatriz[9][40] = 9'b111111111;
assign micromatriz[9][41] = 9'b111111111;
assign micromatriz[9][42] = 9'b111111111;
assign micromatriz[9][43] = 9'b111111111;
assign micromatriz[9][44] = 9'b111111111;
assign micromatriz[9][45] = 9'b111111111;
assign micromatriz[9][46] = 9'b111111111;
assign micromatriz[9][47] = 9'b111111111;
assign micromatriz[9][48] = 9'b111111111;
assign micromatriz[9][49] = 9'b111111111;
assign micromatriz[9][50] = 9'b111111111;
assign micromatriz[9][51] = 9'b111111111;
assign micromatriz[9][52] = 9'b111111111;
assign micromatriz[9][53] = 9'b111111111;
assign micromatriz[9][54] = 9'b111111111;
assign micromatriz[9][55] = 9'b111111111;
assign micromatriz[9][56] = 9'b111111111;
assign micromatriz[9][57] = 9'b111111111;
assign micromatriz[9][58] = 9'b111111111;
assign micromatriz[9][59] = 9'b111111111;
assign micromatriz[9][60] = 9'b111111111;
assign micromatriz[9][61] = 9'b111111111;
assign micromatriz[9][62] = 9'b111111111;
assign micromatriz[9][63] = 9'b111111111;
assign micromatriz[9][64] = 9'b111111111;
assign micromatriz[9][65] = 9'b111111111;
assign micromatriz[9][66] = 9'b111111111;
assign micromatriz[9][67] = 9'b111111111;
assign micromatriz[9][68] = 9'b111111111;
assign micromatriz[9][69] = 9'b111111111;
assign micromatriz[9][70] = 9'b111111111;
assign micromatriz[9][71] = 9'b111111111;
assign micromatriz[9][72] = 9'b111111111;
assign micromatriz[9][73] = 9'b111111111;
assign micromatriz[9][74] = 9'b111111111;
assign micromatriz[9][75] = 9'b111111111;
assign micromatriz[9][76] = 9'b111111111;
assign micromatriz[9][77] = 9'b111111111;
assign micromatriz[9][78] = 9'b111111111;
assign micromatriz[9][79] = 9'b111111111;
assign micromatriz[9][80] = 9'b111111111;
assign micromatriz[9][81] = 9'b111111111;
assign micromatriz[9][82] = 9'b111111111;
assign micromatriz[9][83] = 9'b111111111;
assign micromatriz[9][84] = 9'b111111111;
assign micromatriz[9][85] = 9'b111111111;
assign micromatriz[9][86] = 9'b111111111;
assign micromatriz[9][87] = 9'b111111111;
assign micromatriz[9][88] = 9'b111111111;
assign micromatriz[9][89] = 9'b111111111;
assign micromatriz[9][90] = 9'b111111111;
assign micromatriz[9][91] = 9'b111111111;
assign micromatriz[9][92] = 9'b111111111;
assign micromatriz[9][93] = 9'b111111111;
assign micromatriz[9][94] = 9'b111111111;
assign micromatriz[9][95] = 9'b111111111;
assign micromatriz[9][96] = 9'b111111111;
assign micromatriz[9][97] = 9'b111111111;
assign micromatriz[9][98] = 9'b111111111;
assign micromatriz[9][99] = 9'b111111111;
assign micromatriz[10][0] = 9'b111111111;
assign micromatriz[10][1] = 9'b111111111;
assign micromatriz[10][2] = 9'b111111111;
assign micromatriz[10][3] = 9'b111111111;
assign micromatriz[10][4] = 9'b111111111;
assign micromatriz[10][5] = 9'b111111111;
assign micromatriz[10][6] = 9'b111111111;
assign micromatriz[10][7] = 9'b111111111;
assign micromatriz[10][8] = 9'b111111111;
assign micromatriz[10][9] = 9'b111111111;
assign micromatriz[10][10] = 9'b111111111;
assign micromatriz[10][11] = 9'b111111111;
assign micromatriz[10][12] = 9'b111111111;
assign micromatriz[10][13] = 9'b111111111;
assign micromatriz[10][14] = 9'b111111111;
assign micromatriz[10][15] = 9'b111111111;
assign micromatriz[10][16] = 9'b111111111;
assign micromatriz[10][17] = 9'b111111111;
assign micromatriz[10][18] = 9'b111111111;
assign micromatriz[10][19] = 9'b111111111;
assign micromatriz[10][20] = 9'b111111111;
assign micromatriz[10][21] = 9'b111111111;
assign micromatriz[10][22] = 9'b111111111;
assign micromatriz[10][23] = 9'b111111111;
assign micromatriz[10][24] = 9'b111111111;
assign micromatriz[10][25] = 9'b111111111;
assign micromatriz[10][26] = 9'b111111111;
assign micromatriz[10][27] = 9'b111111111;
assign micromatriz[10][28] = 9'b111111111;
assign micromatriz[10][29] = 9'b111111111;
assign micromatriz[10][30] = 9'b111111111;
assign micromatriz[10][31] = 9'b111111111;
assign micromatriz[10][32] = 9'b111111111;
assign micromatriz[10][33] = 9'b111111111;
assign micromatriz[10][34] = 9'b111111111;
assign micromatriz[10][35] = 9'b111111111;
assign micromatriz[10][36] = 9'b111111111;
assign micromatriz[10][37] = 9'b111111111;
assign micromatriz[10][38] = 9'b111111111;
assign micromatriz[10][39] = 9'b111111111;
assign micromatriz[10][40] = 9'b111111111;
assign micromatriz[10][41] = 9'b111111111;
assign micromatriz[10][42] = 9'b111111111;
assign micromatriz[10][43] = 9'b111111111;
assign micromatriz[10][44] = 9'b111111111;
assign micromatriz[10][45] = 9'b111111111;
assign micromatriz[10][46] = 9'b111111111;
assign micromatriz[10][47] = 9'b111111111;
assign micromatriz[10][48] = 9'b111111111;
assign micromatriz[10][49] = 9'b111111111;
assign micromatriz[10][50] = 9'b111111111;
assign micromatriz[10][51] = 9'b111111111;
assign micromatriz[10][52] = 9'b111111111;
assign micromatriz[10][53] = 9'b111111111;
assign micromatriz[10][54] = 9'b111111111;
assign micromatriz[10][55] = 9'b111111111;
assign micromatriz[10][56] = 9'b111111111;
assign micromatriz[10][57] = 9'b111111111;
assign micromatriz[10][58] = 9'b111111111;
assign micromatriz[10][59] = 9'b111111111;
assign micromatriz[10][60] = 9'b111111111;
assign micromatriz[10][61] = 9'b111111111;
assign micromatriz[10][62] = 9'b111111111;
assign micromatriz[10][63] = 9'b111111111;
assign micromatriz[10][64] = 9'b111111111;
assign micromatriz[10][65] = 9'b111111111;
assign micromatriz[10][66] = 9'b111111111;
assign micromatriz[10][67] = 9'b111111111;
assign micromatriz[10][68] = 9'b111111111;
assign micromatriz[10][69] = 9'b111111111;
assign micromatriz[10][70] = 9'b111111111;
assign micromatriz[10][71] = 9'b111111111;
assign micromatriz[10][72] = 9'b111111111;
assign micromatriz[10][73] = 9'b111111111;
assign micromatriz[10][74] = 9'b111111111;
assign micromatriz[10][75] = 9'b111111111;
assign micromatriz[10][76] = 9'b111111111;
assign micromatriz[10][77] = 9'b111111111;
assign micromatriz[10][78] = 9'b111111111;
assign micromatriz[10][79] = 9'b111111111;
assign micromatriz[10][80] = 9'b111111111;
assign micromatriz[10][81] = 9'b111111111;
assign micromatriz[10][82] = 9'b111111111;
assign micromatriz[10][83] = 9'b111111111;
assign micromatriz[10][84] = 9'b111111111;
assign micromatriz[10][85] = 9'b111111111;
assign micromatriz[10][86] = 9'b111111111;
assign micromatriz[10][87] = 9'b111111111;
assign micromatriz[10][88] = 9'b111111111;
assign micromatriz[10][89] = 9'b111111111;
assign micromatriz[10][90] = 9'b111111111;
assign micromatriz[10][91] = 9'b111111111;
assign micromatriz[10][92] = 9'b111111111;
assign micromatriz[10][93] = 9'b111111111;
assign micromatriz[10][94] = 9'b111111111;
assign micromatriz[10][95] = 9'b111111111;
assign micromatriz[10][96] = 9'b111111111;
assign micromatriz[10][97] = 9'b111111111;
assign micromatriz[10][98] = 9'b111111111;
assign micromatriz[10][99] = 9'b111111111;
assign micromatriz[11][0] = 9'b111111111;
assign micromatriz[11][1] = 9'b111111111;
assign micromatriz[11][2] = 9'b111111111;
assign micromatriz[11][3] = 9'b111111111;
assign micromatriz[11][4] = 9'b111111111;
assign micromatriz[11][5] = 9'b111111111;
assign micromatriz[11][6] = 9'b111111111;
assign micromatriz[11][7] = 9'b111111111;
assign micromatriz[11][8] = 9'b111111111;
assign micromatriz[11][9] = 9'b111111111;
assign micromatriz[11][10] = 9'b111111111;
assign micromatriz[11][11] = 9'b111111111;
assign micromatriz[11][12] = 9'b111111111;
assign micromatriz[11][13] = 9'b111111111;
assign micromatriz[11][14] = 9'b111111111;
assign micromatriz[11][15] = 9'b111111111;
assign micromatriz[11][16] = 9'b111111111;
assign micromatriz[11][17] = 9'b111111111;
assign micromatriz[11][18] = 9'b111111111;
assign micromatriz[11][19] = 9'b111111111;
assign micromatriz[11][20] = 9'b111111111;
assign micromatriz[11][21] = 9'b111111111;
assign micromatriz[11][22] = 9'b111111111;
assign micromatriz[11][23] = 9'b111111111;
assign micromatriz[11][24] = 9'b111111111;
assign micromatriz[11][25] = 9'b111111111;
assign micromatriz[11][26] = 9'b111111111;
assign micromatriz[11][27] = 9'b111111111;
assign micromatriz[11][28] = 9'b111111111;
assign micromatriz[11][29] = 9'b111111111;
assign micromatriz[11][30] = 9'b111111111;
assign micromatriz[11][31] = 9'b111111111;
assign micromatriz[11][32] = 9'b111111111;
assign micromatriz[11][33] = 9'b111111111;
assign micromatriz[11][34] = 9'b111111111;
assign micromatriz[11][35] = 9'b111111111;
assign micromatriz[11][36] = 9'b111111111;
assign micromatriz[11][37] = 9'b111111111;
assign micromatriz[11][38] = 9'b111111111;
assign micromatriz[11][39] = 9'b111111111;
assign micromatriz[11][40] = 9'b111111111;
assign micromatriz[11][41] = 9'b111111111;
assign micromatriz[11][42] = 9'b111111111;
assign micromatriz[11][43] = 9'b111111111;
assign micromatriz[11][44] = 9'b111111111;
assign micromatriz[11][45] = 9'b111111111;
assign micromatriz[11][46] = 9'b111111111;
assign micromatriz[11][47] = 9'b111111111;
assign micromatriz[11][48] = 9'b111111111;
assign micromatriz[11][49] = 9'b111111111;
assign micromatriz[11][50] = 9'b111111111;
assign micromatriz[11][51] = 9'b111111111;
assign micromatriz[11][52] = 9'b111111111;
assign micromatriz[11][53] = 9'b111111111;
assign micromatriz[11][54] = 9'b111111111;
assign micromatriz[11][55] = 9'b111111111;
assign micromatriz[11][56] = 9'b111111111;
assign micromatriz[11][57] = 9'b111111111;
assign micromatriz[11][58] = 9'b111111111;
assign micromatriz[11][59] = 9'b111111111;
assign micromatriz[11][60] = 9'b111111111;
assign micromatriz[11][61] = 9'b111111111;
assign micromatriz[11][62] = 9'b111111111;
assign micromatriz[11][63] = 9'b111111111;
assign micromatriz[11][64] = 9'b111111111;
assign micromatriz[11][65] = 9'b111111111;
assign micromatriz[11][66] = 9'b111111111;
assign micromatriz[11][67] = 9'b111111111;
assign micromatriz[11][68] = 9'b111111111;
assign micromatriz[11][69] = 9'b111111111;
assign micromatriz[11][70] = 9'b111111111;
assign micromatriz[11][71] = 9'b111111111;
assign micromatriz[11][72] = 9'b111111111;
assign micromatriz[11][73] = 9'b111111111;
assign micromatriz[11][74] = 9'b111111111;
assign micromatriz[11][75] = 9'b111111111;
assign micromatriz[11][76] = 9'b111111111;
assign micromatriz[11][77] = 9'b111111111;
assign micromatriz[11][78] = 9'b111111111;
assign micromatriz[11][79] = 9'b111111111;
assign micromatriz[11][80] = 9'b111111111;
assign micromatriz[11][81] = 9'b111111111;
assign micromatriz[11][82] = 9'b111111111;
assign micromatriz[11][83] = 9'b111111111;
assign micromatriz[11][84] = 9'b111111111;
assign micromatriz[11][85] = 9'b111111111;
assign micromatriz[11][86] = 9'b111111111;
assign micromatriz[11][87] = 9'b111111111;
assign micromatriz[11][88] = 9'b111111111;
assign micromatriz[11][89] = 9'b111111111;
assign micromatriz[11][90] = 9'b111111111;
assign micromatriz[11][91] = 9'b111111111;
assign micromatriz[11][92] = 9'b111111111;
assign micromatriz[11][93] = 9'b111111111;
assign micromatriz[11][94] = 9'b111111111;
assign micromatriz[11][95] = 9'b111111111;
assign micromatriz[11][96] = 9'b111111111;
assign micromatriz[11][97] = 9'b111111111;
assign micromatriz[11][98] = 9'b111111111;
assign micromatriz[11][99] = 9'b111111111;
assign micromatriz[12][0] = 9'b111111111;
assign micromatriz[12][1] = 9'b111111111;
assign micromatriz[12][2] = 9'b111111111;
assign micromatriz[12][3] = 9'b111111111;
assign micromatriz[12][4] = 9'b111111111;
assign micromatriz[12][5] = 9'b111111111;
assign micromatriz[12][6] = 9'b111111111;
assign micromatriz[12][7] = 9'b111111111;
assign micromatriz[12][8] = 9'b111111111;
assign micromatriz[12][9] = 9'b111111111;
assign micromatriz[12][10] = 9'b111111111;
assign micromatriz[12][11] = 9'b111111111;
assign micromatriz[12][12] = 9'b111111111;
assign micromatriz[12][13] = 9'b111111111;
assign micromatriz[12][14] = 9'b111111111;
assign micromatriz[12][15] = 9'b111111111;
assign micromatriz[12][16] = 9'b111111111;
assign micromatriz[12][17] = 9'b111111111;
assign micromatriz[12][18] = 9'b111111111;
assign micromatriz[12][19] = 9'b111111111;
assign micromatriz[12][20] = 9'b111111111;
assign micromatriz[12][21] = 9'b111111111;
assign micromatriz[12][22] = 9'b111111111;
assign micromatriz[12][23] = 9'b111111111;
assign micromatriz[12][24] = 9'b111111111;
assign micromatriz[12][25] = 9'b111111111;
assign micromatriz[12][26] = 9'b111111111;
assign micromatriz[12][27] = 9'b111111111;
assign micromatriz[12][28] = 9'b111111111;
assign micromatriz[12][29] = 9'b111111111;
assign micromatriz[12][30] = 9'b111111111;
assign micromatriz[12][31] = 9'b111111111;
assign micromatriz[12][32] = 9'b111111111;
assign micromatriz[12][33] = 9'b111111111;
assign micromatriz[12][34] = 9'b111111111;
assign micromatriz[12][35] = 9'b111111111;
assign micromatriz[12][36] = 9'b111111111;
assign micromatriz[12][37] = 9'b111111111;
assign micromatriz[12][38] = 9'b111111111;
assign micromatriz[12][39] = 9'b111111111;
assign micromatriz[12][40] = 9'b111111111;
assign micromatriz[12][41] = 9'b111111111;
assign micromatriz[12][42] = 9'b111111111;
assign micromatriz[12][43] = 9'b111111111;
assign micromatriz[12][44] = 9'b111111111;
assign micromatriz[12][45] = 9'b111111111;
assign micromatriz[12][46] = 9'b111111111;
assign micromatriz[12][47] = 9'b111111111;
assign micromatriz[12][48] = 9'b111111111;
assign micromatriz[12][49] = 9'b111111111;
assign micromatriz[12][50] = 9'b111111111;
assign micromatriz[12][51] = 9'b111111111;
assign micromatriz[12][52] = 9'b111111111;
assign micromatriz[12][53] = 9'b111111111;
assign micromatriz[12][54] = 9'b111111111;
assign micromatriz[12][55] = 9'b111111111;
assign micromatriz[12][56] = 9'b111111111;
assign micromatriz[12][57] = 9'b111111111;
assign micromatriz[12][58] = 9'b111111111;
assign micromatriz[12][59] = 9'b111111111;
assign micromatriz[12][60] = 9'b111111111;
assign micromatriz[12][61] = 9'b111111111;
assign micromatriz[12][62] = 9'b111111111;
assign micromatriz[12][63] = 9'b111111111;
assign micromatriz[12][64] = 9'b111111111;
assign micromatriz[12][65] = 9'b111111111;
assign micromatriz[12][66] = 9'b111111111;
assign micromatriz[12][67] = 9'b111111111;
assign micromatriz[12][68] = 9'b111111111;
assign micromatriz[12][69] = 9'b111111111;
assign micromatriz[12][70] = 9'b111111111;
assign micromatriz[12][71] = 9'b111111111;
assign micromatriz[12][72] = 9'b111111111;
assign micromatriz[12][73] = 9'b111111111;
assign micromatriz[12][74] = 9'b111111111;
assign micromatriz[12][75] = 9'b111111111;
assign micromatriz[12][76] = 9'b111111111;
assign micromatriz[12][77] = 9'b111111111;
assign micromatriz[12][78] = 9'b111111111;
assign micromatriz[12][79] = 9'b111111111;
assign micromatriz[12][80] = 9'b111111111;
assign micromatriz[12][81] = 9'b111111111;
assign micromatriz[12][82] = 9'b111111111;
assign micromatriz[12][83] = 9'b111111111;
assign micromatriz[12][84] = 9'b111111111;
assign micromatriz[12][85] = 9'b111111111;
assign micromatriz[12][86] = 9'b111111111;
assign micromatriz[12][87] = 9'b111111111;
assign micromatriz[12][88] = 9'b111111111;
assign micromatriz[12][89] = 9'b111111111;
assign micromatriz[12][90] = 9'b111111111;
assign micromatriz[12][91] = 9'b111111111;
assign micromatriz[12][92] = 9'b111111111;
assign micromatriz[12][93] = 9'b111111111;
assign micromatriz[12][94] = 9'b111111111;
assign micromatriz[12][95] = 9'b111111111;
assign micromatriz[12][96] = 9'b111111111;
assign micromatriz[12][97] = 9'b111111111;
assign micromatriz[12][98] = 9'b111111111;
assign micromatriz[12][99] = 9'b111111111;
assign micromatriz[13][0] = 9'b111111111;
assign micromatriz[13][1] = 9'b111111111;
assign micromatriz[13][2] = 9'b111111111;
assign micromatriz[13][3] = 9'b111111111;
assign micromatriz[13][4] = 9'b111111111;
assign micromatriz[13][5] = 9'b111111111;
assign micromatriz[13][6] = 9'b111111111;
assign micromatriz[13][7] = 9'b111111111;
assign micromatriz[13][8] = 9'b111111111;
assign micromatriz[13][9] = 9'b111111111;
assign micromatriz[13][10] = 9'b111111111;
assign micromatriz[13][11] = 9'b111111111;
assign micromatriz[13][12] = 9'b111111111;
assign micromatriz[13][13] = 9'b111111111;
assign micromatriz[13][14] = 9'b111111111;
assign micromatriz[13][15] = 9'b111111111;
assign micromatriz[13][16] = 9'b111111111;
assign micromatriz[13][17] = 9'b111111111;
assign micromatriz[13][18] = 9'b111111111;
assign micromatriz[13][19] = 9'b111111111;
assign micromatriz[13][20] = 9'b111111111;
assign micromatriz[13][21] = 9'b111111111;
assign micromatriz[13][22] = 9'b111111111;
assign micromatriz[13][23] = 9'b111111111;
assign micromatriz[13][24] = 9'b111111111;
assign micromatriz[13][25] = 9'b111111111;
assign micromatriz[13][26] = 9'b111111111;
assign micromatriz[13][27] = 9'b111111111;
assign micromatriz[13][28] = 9'b111111111;
assign micromatriz[13][29] = 9'b111111111;
assign micromatriz[13][30] = 9'b111111111;
assign micromatriz[13][31] = 9'b111111111;
assign micromatriz[13][32] = 9'b111111111;
assign micromatriz[13][33] = 9'b111111111;
assign micromatriz[13][34] = 9'b111111111;
assign micromatriz[13][35] = 9'b111111111;
assign micromatriz[13][36] = 9'b111111111;
assign micromatriz[13][37] = 9'b111111111;
assign micromatriz[13][38] = 9'b111111111;
assign micromatriz[13][39] = 9'b111111111;
assign micromatriz[13][40] = 9'b111111111;
assign micromatriz[13][41] = 9'b111111111;
assign micromatriz[13][42] = 9'b111111111;
assign micromatriz[13][43] = 9'b111111111;
assign micromatriz[13][44] = 9'b111111111;
assign micromatriz[13][45] = 9'b111111111;
assign micromatriz[13][46] = 9'b111111111;
assign micromatriz[13][47] = 9'b111111111;
assign micromatriz[13][48] = 9'b111111111;
assign micromatriz[13][49] = 9'b111111111;
assign micromatriz[13][50] = 9'b111111111;
assign micromatriz[13][51] = 9'b111111111;
assign micromatriz[13][52] = 9'b111111111;
assign micromatriz[13][53] = 9'b111111111;
assign micromatriz[13][54] = 9'b111111111;
assign micromatriz[13][55] = 9'b111111111;
assign micromatriz[13][56] = 9'b111111111;
assign micromatriz[13][57] = 9'b111111111;
assign micromatriz[13][58] = 9'b111111111;
assign micromatriz[13][59] = 9'b111111111;
assign micromatriz[13][60] = 9'b111111111;
assign micromatriz[13][61] = 9'b111111111;
assign micromatriz[13][62] = 9'b111111111;
assign micromatriz[13][63] = 9'b111111111;
assign micromatriz[13][64] = 9'b111111111;
assign micromatriz[13][65] = 9'b111111111;
assign micromatriz[13][66] = 9'b111111111;
assign micromatriz[13][67] = 9'b111111111;
assign micromatriz[13][68] = 9'b111111111;
assign micromatriz[13][69] = 9'b111111111;
assign micromatriz[13][70] = 9'b111111111;
assign micromatriz[13][71] = 9'b111111111;
assign micromatriz[13][72] = 9'b111111111;
assign micromatriz[13][73] = 9'b111111111;
assign micromatriz[13][74] = 9'b111111111;
assign micromatriz[13][75] = 9'b111111111;
assign micromatriz[13][76] = 9'b111111111;
assign micromatriz[13][77] = 9'b111111111;
assign micromatriz[13][78] = 9'b111111111;
assign micromatriz[13][79] = 9'b111111111;
assign micromatriz[13][80] = 9'b111111111;
assign micromatriz[13][81] = 9'b111111111;
assign micromatriz[13][82] = 9'b111111111;
assign micromatriz[13][83] = 9'b111111111;
assign micromatriz[13][84] = 9'b111111111;
assign micromatriz[13][85] = 9'b111111111;
assign micromatriz[13][86] = 9'b111111111;
assign micromatriz[13][87] = 9'b111111111;
assign micromatriz[13][88] = 9'b111111111;
assign micromatriz[13][89] = 9'b111111111;
assign micromatriz[13][90] = 9'b111111111;
assign micromatriz[13][91] = 9'b111111111;
assign micromatriz[13][92] = 9'b111111111;
assign micromatriz[13][93] = 9'b111111111;
assign micromatriz[13][94] = 9'b111111111;
assign micromatriz[13][95] = 9'b111111111;
assign micromatriz[13][96] = 9'b111111111;
assign micromatriz[13][97] = 9'b111111111;
assign micromatriz[13][98] = 9'b111111111;
assign micromatriz[13][99] = 9'b111111111;
assign micromatriz[14][0] = 9'b111111111;
assign micromatriz[14][1] = 9'b111111111;
assign micromatriz[14][2] = 9'b111111111;
assign micromatriz[14][3] = 9'b111111111;
assign micromatriz[14][4] = 9'b111111111;
assign micromatriz[14][5] = 9'b111111111;
assign micromatriz[14][6] = 9'b111111111;
assign micromatriz[14][7] = 9'b111111111;
assign micromatriz[14][8] = 9'b111111111;
assign micromatriz[14][9] = 9'b111111111;
assign micromatriz[14][10] = 9'b111111111;
assign micromatriz[14][11] = 9'b111111111;
assign micromatriz[14][12] = 9'b111111111;
assign micromatriz[14][13] = 9'b111111111;
assign micromatriz[14][14] = 9'b111111111;
assign micromatriz[14][15] = 9'b111111111;
assign micromatriz[14][16] = 9'b111111111;
assign micromatriz[14][17] = 9'b111111111;
assign micromatriz[14][18] = 9'b111111111;
assign micromatriz[14][19] = 9'b111111111;
assign micromatriz[14][20] = 9'b111111111;
assign micromatriz[14][21] = 9'b111111111;
assign micromatriz[14][22] = 9'b111111111;
assign micromatriz[14][23] = 9'b111111111;
assign micromatriz[14][24] = 9'b111111111;
assign micromatriz[14][25] = 9'b111111111;
assign micromatriz[14][26] = 9'b111111111;
assign micromatriz[14][27] = 9'b111111111;
assign micromatriz[14][28] = 9'b111111111;
assign micromatriz[14][29] = 9'b111111111;
assign micromatriz[14][30] = 9'b111111111;
assign micromatriz[14][31] = 9'b111111111;
assign micromatriz[14][32] = 9'b111111111;
assign micromatriz[14][33] = 9'b111111111;
assign micromatriz[14][34] = 9'b111111111;
assign micromatriz[14][35] = 9'b111111111;
assign micromatriz[14][36] = 9'b111111111;
assign micromatriz[14][37] = 9'b111111111;
assign micromatriz[14][38] = 9'b111111111;
assign micromatriz[14][39] = 9'b111111111;
assign micromatriz[14][40] = 9'b111111111;
assign micromatriz[14][41] = 9'b111111111;
assign micromatriz[14][42] = 9'b111111111;
assign micromatriz[14][43] = 9'b111111111;
assign micromatriz[14][44] = 9'b111111111;
assign micromatriz[14][45] = 9'b111111111;
assign micromatriz[14][46] = 9'b111111111;
assign micromatriz[14][47] = 9'b111111111;
assign micromatriz[14][48] = 9'b111111111;
assign micromatriz[14][49] = 9'b111111111;
assign micromatriz[14][50] = 9'b111111111;
assign micromatriz[14][51] = 9'b111111111;
assign micromatriz[14][52] = 9'b111111111;
assign micromatriz[14][53] = 9'b111111111;
assign micromatriz[14][54] = 9'b111111111;
assign micromatriz[14][55] = 9'b111111111;
assign micromatriz[14][56] = 9'b111111111;
assign micromatriz[14][57] = 9'b111111111;
assign micromatriz[14][58] = 9'b111111111;
assign micromatriz[14][59] = 9'b111111111;
assign micromatriz[14][60] = 9'b111111111;
assign micromatriz[14][61] = 9'b111111111;
assign micromatriz[14][62] = 9'b111111111;
assign micromatriz[14][63] = 9'b111111111;
assign micromatriz[14][64] = 9'b111111111;
assign micromatriz[14][65] = 9'b111111111;
assign micromatriz[14][66] = 9'b111111111;
assign micromatriz[14][67] = 9'b111111111;
assign micromatriz[14][68] = 9'b111111111;
assign micromatriz[14][69] = 9'b111111111;
assign micromatriz[14][70] = 9'b111111111;
assign micromatriz[14][71] = 9'b111111111;
assign micromatriz[14][72] = 9'b111111111;
assign micromatriz[14][73] = 9'b111111111;
assign micromatriz[14][74] = 9'b111111111;
assign micromatriz[14][75] = 9'b111111111;
assign micromatriz[14][76] = 9'b111111111;
assign micromatriz[14][77] = 9'b111111111;
assign micromatriz[14][78] = 9'b111111111;
assign micromatriz[14][79] = 9'b111111111;
assign micromatriz[14][80] = 9'b111111111;
assign micromatriz[14][81] = 9'b111111111;
assign micromatriz[14][82] = 9'b111111111;
assign micromatriz[14][83] = 9'b111111111;
assign micromatriz[14][84] = 9'b111111111;
assign micromatriz[14][85] = 9'b111111111;
assign micromatriz[14][86] = 9'b111111111;
assign micromatriz[14][87] = 9'b111111111;
assign micromatriz[14][88] = 9'b111111111;
assign micromatriz[14][89] = 9'b111111111;
assign micromatriz[14][90] = 9'b111111111;
assign micromatriz[14][91] = 9'b111111111;
assign micromatriz[14][92] = 9'b111111111;
assign micromatriz[14][93] = 9'b111111111;
assign micromatriz[14][94] = 9'b111111111;
assign micromatriz[14][95] = 9'b111111111;
assign micromatriz[14][96] = 9'b111111111;
assign micromatriz[14][97] = 9'b111111111;
assign micromatriz[14][98] = 9'b111111111;
assign micromatriz[14][99] = 9'b111111111;
assign micromatriz[15][0] = 9'b111111111;
assign micromatriz[15][1] = 9'b111111111;
assign micromatriz[15][2] = 9'b111111111;
assign micromatriz[15][3] = 9'b111111111;
assign micromatriz[15][4] = 9'b111111111;
assign micromatriz[15][5] = 9'b111111111;
assign micromatriz[15][6] = 9'b111111111;
assign micromatriz[15][7] = 9'b111111111;
assign micromatriz[15][8] = 9'b111111111;
assign micromatriz[15][9] = 9'b111111111;
assign micromatriz[15][10] = 9'b111111111;
assign micromatriz[15][11] = 9'b111111111;
assign micromatriz[15][12] = 9'b111111111;
assign micromatriz[15][13] = 9'b111111111;
assign micromatriz[15][14] = 9'b111111111;
assign micromatriz[15][15] = 9'b111111111;
assign micromatriz[15][16] = 9'b111111111;
assign micromatriz[15][17] = 9'b111111111;
assign micromatriz[15][18] = 9'b111111111;
assign micromatriz[15][19] = 9'b111111111;
assign micromatriz[15][20] = 9'b111111111;
assign micromatriz[15][21] = 9'b111111111;
assign micromatriz[15][22] = 9'b111111111;
assign micromatriz[15][23] = 9'b111111111;
assign micromatriz[15][24] = 9'b111111111;
assign micromatriz[15][25] = 9'b111111111;
assign micromatriz[15][26] = 9'b111111111;
assign micromatriz[15][27] = 9'b111111111;
assign micromatriz[15][28] = 9'b111111111;
assign micromatriz[15][29] = 9'b111111111;
assign micromatriz[15][30] = 9'b111111111;
assign micromatriz[15][31] = 9'b111111111;
assign micromatriz[15][32] = 9'b111111111;
assign micromatriz[15][33] = 9'b111111111;
assign micromatriz[15][34] = 9'b111111111;
assign micromatriz[15][35] = 9'b111111111;
assign micromatriz[15][36] = 9'b111111111;
assign micromatriz[15][37] = 9'b111111111;
assign micromatriz[15][38] = 9'b111111111;
assign micromatriz[15][39] = 9'b111111111;
assign micromatriz[15][40] = 9'b111111111;
assign micromatriz[15][41] = 9'b111111111;
assign micromatriz[15][42] = 9'b111111111;
assign micromatriz[15][43] = 9'b111111111;
assign micromatriz[15][44] = 9'b111111111;
assign micromatriz[15][45] = 9'b111111111;
assign micromatriz[15][46] = 9'b111111111;
assign micromatriz[15][47] = 9'b111111111;
assign micromatriz[15][48] = 9'b111111111;
assign micromatriz[15][49] = 9'b111111111;
assign micromatriz[15][50] = 9'b111111111;
assign micromatriz[15][51] = 9'b111111111;
assign micromatriz[15][52] = 9'b111111111;
assign micromatriz[15][53] = 9'b111111111;
assign micromatriz[15][54] = 9'b111111111;
assign micromatriz[15][55] = 9'b111111111;
assign micromatriz[15][56] = 9'b111111111;
assign micromatriz[15][57] = 9'b111111111;
assign micromatriz[15][58] = 9'b111111111;
assign micromatriz[15][59] = 9'b111111111;
assign micromatriz[15][60] = 9'b111111111;
assign micromatriz[15][61] = 9'b111111111;
assign micromatriz[15][62] = 9'b111111111;
assign micromatriz[15][63] = 9'b111111111;
assign micromatriz[15][64] = 9'b111111111;
assign micromatriz[15][65] = 9'b111111111;
assign micromatriz[15][66] = 9'b111111111;
assign micromatriz[15][67] = 9'b111111111;
assign micromatriz[15][68] = 9'b111111111;
assign micromatriz[15][69] = 9'b111111111;
assign micromatriz[15][70] = 9'b111111111;
assign micromatriz[15][71] = 9'b111111111;
assign micromatriz[15][72] = 9'b111111111;
assign micromatriz[15][73] = 9'b111111111;
assign micromatriz[15][74] = 9'b111111111;
assign micromatriz[15][75] = 9'b111111111;
assign micromatriz[15][76] = 9'b111111111;
assign micromatriz[15][77] = 9'b111111111;
assign micromatriz[15][78] = 9'b111111111;
assign micromatriz[15][79] = 9'b111111111;
assign micromatriz[15][80] = 9'b111111111;
assign micromatriz[15][81] = 9'b111111111;
assign micromatriz[15][82] = 9'b111111111;
assign micromatriz[15][83] = 9'b111111111;
assign micromatriz[15][84] = 9'b111111111;
assign micromatriz[15][85] = 9'b111111111;
assign micromatriz[15][86] = 9'b111111111;
assign micromatriz[15][87] = 9'b111111111;
assign micromatriz[15][88] = 9'b111111111;
assign micromatriz[15][89] = 9'b111111111;
assign micromatriz[15][90] = 9'b111111111;
assign micromatriz[15][91] = 9'b111111111;
assign micromatriz[15][92] = 9'b111111111;
assign micromatriz[15][93] = 9'b111111111;
assign micromatriz[15][94] = 9'b111111111;
assign micromatriz[15][95] = 9'b111111111;
assign micromatriz[15][96] = 9'b111111111;
assign micromatriz[15][97] = 9'b111111111;
assign micromatriz[15][98] = 9'b111111111;
assign micromatriz[15][99] = 9'b111111111;
assign micromatriz[16][0] = 9'b111111111;
assign micromatriz[16][1] = 9'b111111111;
assign micromatriz[16][2] = 9'b111111111;
assign micromatriz[16][3] = 9'b111111111;
assign micromatriz[16][4] = 9'b111111111;
assign micromatriz[16][5] = 9'b111111111;
assign micromatriz[16][6] = 9'b111111111;
assign micromatriz[16][7] = 9'b111111111;
assign micromatriz[16][8] = 9'b111111111;
assign micromatriz[16][9] = 9'b111111111;
assign micromatriz[16][10] = 9'b111111111;
assign micromatriz[16][11] = 9'b111111111;
assign micromatriz[16][12] = 9'b111111111;
assign micromatriz[16][13] = 9'b111111111;
assign micromatriz[16][14] = 9'b111111111;
assign micromatriz[16][15] = 9'b111111111;
assign micromatriz[16][16] = 9'b111111111;
assign micromatriz[16][17] = 9'b111111111;
assign micromatriz[16][18] = 9'b111111111;
assign micromatriz[16][19] = 9'b111111111;
assign micromatriz[16][20] = 9'b111111111;
assign micromatriz[16][21] = 9'b111111111;
assign micromatriz[16][22] = 9'b111111111;
assign micromatriz[16][23] = 9'b111111111;
assign micromatriz[16][24] = 9'b111111111;
assign micromatriz[16][25] = 9'b111111111;
assign micromatriz[16][26] = 9'b111111111;
assign micromatriz[16][27] = 9'b111111111;
assign micromatriz[16][28] = 9'b111111111;
assign micromatriz[16][29] = 9'b111111111;
assign micromatriz[16][30] = 9'b111111111;
assign micromatriz[16][31] = 9'b111111111;
assign micromatriz[16][32] = 9'b111111111;
assign micromatriz[16][33] = 9'b111111111;
assign micromatriz[16][34] = 9'b111111111;
assign micromatriz[16][35] = 9'b111111111;
assign micromatriz[16][36] = 9'b111111111;
assign micromatriz[16][37] = 9'b111111111;
assign micromatriz[16][38] = 9'b111111111;
assign micromatriz[16][39] = 9'b111111111;
assign micromatriz[16][40] = 9'b111111111;
assign micromatriz[16][41] = 9'b111111111;
assign micromatriz[16][42] = 9'b111111111;
assign micromatriz[16][43] = 9'b111111111;
assign micromatriz[16][44] = 9'b111111111;
assign micromatriz[16][45] = 9'b111111111;
assign micromatriz[16][46] = 9'b111111111;
assign micromatriz[16][47] = 9'b111111111;
assign micromatriz[16][48] = 9'b111111111;
assign micromatriz[16][49] = 9'b111111111;
assign micromatriz[16][50] = 9'b111111111;
assign micromatriz[16][51] = 9'b111111111;
assign micromatriz[16][52] = 9'b111111111;
assign micromatriz[16][53] = 9'b111111111;
assign micromatriz[16][54] = 9'b111111111;
assign micromatriz[16][55] = 9'b111111111;
assign micromatriz[16][56] = 9'b111111111;
assign micromatriz[16][57] = 9'b111111111;
assign micromatriz[16][58] = 9'b111111111;
assign micromatriz[16][59] = 9'b111111111;
assign micromatriz[16][60] = 9'b111111111;
assign micromatriz[16][61] = 9'b111111111;
assign micromatriz[16][62] = 9'b111111111;
assign micromatriz[16][63] = 9'b111111111;
assign micromatriz[16][64] = 9'b111111111;
assign micromatriz[16][65] = 9'b111111111;
assign micromatriz[16][66] = 9'b111111111;
assign micromatriz[16][67] = 9'b111111111;
assign micromatriz[16][68] = 9'b111111111;
assign micromatriz[16][69] = 9'b111111111;
assign micromatriz[16][70] = 9'b111111111;
assign micromatriz[16][71] = 9'b111111111;
assign micromatriz[16][72] = 9'b111111111;
assign micromatriz[16][73] = 9'b111111111;
assign micromatriz[16][74] = 9'b111111111;
assign micromatriz[16][75] = 9'b111111111;
assign micromatriz[16][76] = 9'b111111111;
assign micromatriz[16][77] = 9'b111111111;
assign micromatriz[16][78] = 9'b111111111;
assign micromatriz[16][79] = 9'b111111111;
assign micromatriz[16][80] = 9'b111111111;
assign micromatriz[16][81] = 9'b111111111;
assign micromatriz[16][82] = 9'b111111111;
assign micromatriz[16][83] = 9'b111111111;
assign micromatriz[16][84] = 9'b111111111;
assign micromatriz[16][85] = 9'b111111111;
assign micromatriz[16][86] = 9'b111111111;
assign micromatriz[16][87] = 9'b111111111;
assign micromatriz[16][88] = 9'b111111111;
assign micromatriz[16][89] = 9'b111111111;
assign micromatriz[16][90] = 9'b111111111;
assign micromatriz[16][91] = 9'b111111111;
assign micromatriz[16][92] = 9'b111111111;
assign micromatriz[16][93] = 9'b111111111;
assign micromatriz[16][94] = 9'b111111111;
assign micromatriz[16][95] = 9'b111111111;
assign micromatriz[16][96] = 9'b111111111;
assign micromatriz[16][97] = 9'b111111111;
assign micromatriz[16][98] = 9'b111111111;
assign micromatriz[16][99] = 9'b111111111;
assign micromatriz[17][0] = 9'b111111111;
assign micromatriz[17][1] = 9'b111111111;
assign micromatriz[17][2] = 9'b111111111;
assign micromatriz[17][3] = 9'b111111111;
assign micromatriz[17][4] = 9'b111111111;
assign micromatriz[17][5] = 9'b111111111;
assign micromatriz[17][6] = 9'b111111111;
assign micromatriz[17][7] = 9'b111111111;
assign micromatriz[17][8] = 9'b111111111;
assign micromatriz[17][9] = 9'b111111111;
assign micromatriz[17][10] = 9'b111111111;
assign micromatriz[17][11] = 9'b111111111;
assign micromatriz[17][12] = 9'b111111111;
assign micromatriz[17][13] = 9'b111111111;
assign micromatriz[17][14] = 9'b111111111;
assign micromatriz[17][15] = 9'b111111111;
assign micromatriz[17][16] = 9'b111111111;
assign micromatriz[17][17] = 9'b111111111;
assign micromatriz[17][18] = 9'b111111111;
assign micromatriz[17][19] = 9'b111111111;
assign micromatriz[17][20] = 9'b111111111;
assign micromatriz[17][21] = 9'b111111111;
assign micromatriz[17][22] = 9'b111111111;
assign micromatriz[17][23] = 9'b111111111;
assign micromatriz[17][24] = 9'b111111111;
assign micromatriz[17][25] = 9'b111111111;
assign micromatriz[17][26] = 9'b111111111;
assign micromatriz[17][27] = 9'b111111111;
assign micromatriz[17][28] = 9'b111111111;
assign micromatriz[17][29] = 9'b111111111;
assign micromatriz[17][30] = 9'b111111111;
assign micromatriz[17][31] = 9'b111111111;
assign micromatriz[17][32] = 9'b111111111;
assign micromatriz[17][33] = 9'b111111111;
assign micromatriz[17][34] = 9'b111111111;
assign micromatriz[17][35] = 9'b111111111;
assign micromatriz[17][36] = 9'b111111111;
assign micromatriz[17][37] = 9'b111111111;
assign micromatriz[17][38] = 9'b111111111;
assign micromatriz[17][39] = 9'b111111111;
assign micromatriz[17][40] = 9'b111111111;
assign micromatriz[17][41] = 9'b111111111;
assign micromatriz[17][42] = 9'b111111111;
assign micromatriz[17][43] = 9'b111111111;
assign micromatriz[17][44] = 9'b111111111;
assign micromatriz[17][45] = 9'b111111111;
assign micromatriz[17][46] = 9'b111111111;
assign micromatriz[17][47] = 9'b111111111;
assign micromatriz[17][48] = 9'b111111111;
assign micromatriz[17][49] = 9'b111111111;
assign micromatriz[17][50] = 9'b111111111;
assign micromatriz[17][51] = 9'b111111111;
assign micromatriz[17][52] = 9'b111111111;
assign micromatriz[17][53] = 9'b111111111;
assign micromatriz[17][54] = 9'b111111111;
assign micromatriz[17][55] = 9'b111111111;
assign micromatriz[17][56] = 9'b111111111;
assign micromatriz[17][57] = 9'b111111111;
assign micromatriz[17][58] = 9'b111111111;
assign micromatriz[17][59] = 9'b111111111;
assign micromatriz[17][60] = 9'b111111111;
assign micromatriz[17][61] = 9'b111111111;
assign micromatriz[17][62] = 9'b111111111;
assign micromatriz[17][63] = 9'b111111111;
assign micromatriz[17][64] = 9'b111111111;
assign micromatriz[17][65] = 9'b111111111;
assign micromatriz[17][66] = 9'b111111111;
assign micromatriz[17][67] = 9'b111111111;
assign micromatriz[17][68] = 9'b111111111;
assign micromatriz[17][69] = 9'b111111111;
assign micromatriz[17][70] = 9'b111111111;
assign micromatriz[17][71] = 9'b111111111;
assign micromatriz[17][72] = 9'b111111111;
assign micromatriz[17][73] = 9'b111111111;
assign micromatriz[17][74] = 9'b111111111;
assign micromatriz[17][75] = 9'b111111111;
assign micromatriz[17][76] = 9'b111111111;
assign micromatriz[17][77] = 9'b111111111;
assign micromatriz[17][78] = 9'b111111111;
assign micromatriz[17][79] = 9'b111111111;
assign micromatriz[17][80] = 9'b111111111;
assign micromatriz[17][81] = 9'b111111111;
assign micromatriz[17][82] = 9'b111111111;
assign micromatriz[17][83] = 9'b111111111;
assign micromatriz[17][84] = 9'b111111111;
assign micromatriz[17][85] = 9'b111111111;
assign micromatriz[17][86] = 9'b111111111;
assign micromatriz[17][87] = 9'b111111111;
assign micromatriz[17][88] = 9'b111111111;
assign micromatriz[17][89] = 9'b111111111;
assign micromatriz[17][90] = 9'b111111111;
assign micromatriz[17][91] = 9'b111111111;
assign micromatriz[17][92] = 9'b111111111;
assign micromatriz[17][93] = 9'b111111111;
assign micromatriz[17][94] = 9'b111111111;
assign micromatriz[17][95] = 9'b111111111;
assign micromatriz[17][96] = 9'b111111111;
assign micromatriz[17][97] = 9'b111111111;
assign micromatriz[17][98] = 9'b111111111;
assign micromatriz[17][99] = 9'b111111111;
assign micromatriz[18][0] = 9'b111111111;
assign micromatriz[18][1] = 9'b111111111;
assign micromatriz[18][2] = 9'b111111111;
assign micromatriz[18][3] = 9'b111111111;
assign micromatriz[18][4] = 9'b111111111;
assign micromatriz[18][5] = 9'b111111111;
assign micromatriz[18][6] = 9'b111111111;
assign micromatriz[18][7] = 9'b111111111;
assign micromatriz[18][8] = 9'b111111111;
assign micromatriz[18][9] = 9'b111111111;
assign micromatriz[18][10] = 9'b111111111;
assign micromatriz[18][11] = 9'b111111111;
assign micromatriz[18][12] = 9'b111111111;
assign micromatriz[18][13] = 9'b111111111;
assign micromatriz[18][14] = 9'b111111111;
assign micromatriz[18][15] = 9'b111111111;
assign micromatriz[18][16] = 9'b111111111;
assign micromatriz[18][17] = 9'b111111111;
assign micromatriz[18][18] = 9'b111111111;
assign micromatriz[18][19] = 9'b111111111;
assign micromatriz[18][20] = 9'b111111111;
assign micromatriz[18][21] = 9'b111111111;
assign micromatriz[18][22] = 9'b111111111;
assign micromatriz[18][23] = 9'b111111111;
assign micromatriz[18][24] = 9'b111111111;
assign micromatriz[18][25] = 9'b111111111;
assign micromatriz[18][26] = 9'b111111111;
assign micromatriz[18][27] = 9'b111111111;
assign micromatriz[18][28] = 9'b111111111;
assign micromatriz[18][29] = 9'b111111111;
assign micromatriz[18][30] = 9'b111111111;
assign micromatriz[18][31] = 9'b111111111;
assign micromatriz[18][32] = 9'b111111111;
assign micromatriz[18][33] = 9'b111111111;
assign micromatriz[18][34] = 9'b111111111;
assign micromatriz[18][35] = 9'b111111111;
assign micromatriz[18][36] = 9'b111111111;
assign micromatriz[18][37] = 9'b111111111;
assign micromatriz[18][38] = 9'b111111111;
assign micromatriz[18][39] = 9'b111111111;
assign micromatriz[18][40] = 9'b111111111;
assign micromatriz[18][41] = 9'b111111111;
assign micromatriz[18][42] = 9'b111111111;
assign micromatriz[18][43] = 9'b111111111;
assign micromatriz[18][44] = 9'b111111111;
assign micromatriz[18][45] = 9'b111111111;
assign micromatriz[18][46] = 9'b111111111;
assign micromatriz[18][47] = 9'b111111111;
assign micromatriz[18][48] = 9'b111111111;
assign micromatriz[18][49] = 9'b111111111;
assign micromatriz[18][50] = 9'b111111111;
assign micromatriz[18][51] = 9'b111111111;
assign micromatriz[18][52] = 9'b111111111;
assign micromatriz[18][53] = 9'b111111111;
assign micromatriz[18][54] = 9'b111111111;
assign micromatriz[18][55] = 9'b111111111;
assign micromatriz[18][56] = 9'b111111111;
assign micromatriz[18][57] = 9'b111111111;
assign micromatriz[18][58] = 9'b111111111;
assign micromatriz[18][59] = 9'b111111111;
assign micromatriz[18][60] = 9'b111111111;
assign micromatriz[18][61] = 9'b111111111;
assign micromatriz[18][62] = 9'b111111111;
assign micromatriz[18][63] = 9'b111111111;
assign micromatriz[18][64] = 9'b111111111;
assign micromatriz[18][65] = 9'b111111111;
assign micromatriz[18][66] = 9'b111111111;
assign micromatriz[18][67] = 9'b111111111;
assign micromatriz[18][68] = 9'b111111111;
assign micromatriz[18][69] = 9'b111111111;
assign micromatriz[18][70] = 9'b111111111;
assign micromatriz[18][71] = 9'b111111111;
assign micromatriz[18][72] = 9'b111111111;
assign micromatriz[18][73] = 9'b111111111;
assign micromatriz[18][74] = 9'b111111111;
assign micromatriz[18][75] = 9'b111111111;
assign micromatriz[18][76] = 9'b111111111;
assign micromatriz[18][77] = 9'b111111111;
assign micromatriz[18][78] = 9'b111111111;
assign micromatriz[18][79] = 9'b111111111;
assign micromatriz[18][80] = 9'b111111111;
assign micromatriz[18][81] = 9'b111111111;
assign micromatriz[18][82] = 9'b111111111;
assign micromatriz[18][83] = 9'b111111111;
assign micromatriz[18][84] = 9'b111111111;
assign micromatriz[18][85] = 9'b111111111;
assign micromatriz[18][86] = 9'b111111111;
assign micromatriz[18][87] = 9'b111111111;
assign micromatriz[18][88] = 9'b111111111;
assign micromatriz[18][89] = 9'b111111111;
assign micromatriz[18][90] = 9'b111111111;
assign micromatriz[18][91] = 9'b111111111;
assign micromatriz[18][92] = 9'b111111111;
assign micromatriz[18][93] = 9'b111111111;
assign micromatriz[18][94] = 9'b111111111;
assign micromatriz[18][95] = 9'b111111111;
assign micromatriz[18][96] = 9'b111111111;
assign micromatriz[18][97] = 9'b111111111;
assign micromatriz[18][98] = 9'b111111111;
assign micromatriz[18][99] = 9'b111111111;
assign micromatriz[19][0] = 9'b111111111;
assign micromatriz[19][1] = 9'b111111111;
assign micromatriz[19][2] = 9'b111111111;
assign micromatriz[19][3] = 9'b111111111;
assign micromatriz[19][4] = 9'b111111111;
assign micromatriz[19][5] = 9'b111111111;
assign micromatriz[19][6] = 9'b111111111;
assign micromatriz[19][7] = 9'b111111111;
assign micromatriz[19][8] = 9'b111111111;
assign micromatriz[19][9] = 9'b111111111;
assign micromatriz[19][10] = 9'b111111111;
assign micromatriz[19][11] = 9'b111111111;
assign micromatriz[19][12] = 9'b111111111;
assign micromatriz[19][13] = 9'b111111111;
assign micromatriz[19][14] = 9'b111111111;
assign micromatriz[19][15] = 9'b111111111;
assign micromatriz[19][16] = 9'b111111111;
assign micromatriz[19][17] = 9'b111111111;
assign micromatriz[19][18] = 9'b111111111;
assign micromatriz[19][19] = 9'b111111111;
assign micromatriz[19][20] = 9'b111111111;
assign micromatriz[19][21] = 9'b111111111;
assign micromatriz[19][22] = 9'b111111111;
assign micromatriz[19][23] = 9'b111111111;
assign micromatriz[19][24] = 9'b111111111;
assign micromatriz[19][25] = 9'b111111111;
assign micromatriz[19][26] = 9'b111111111;
assign micromatriz[19][27] = 9'b111111111;
assign micromatriz[19][28] = 9'b111111111;
assign micromatriz[19][29] = 9'b111111111;
assign micromatriz[19][30] = 9'b111111111;
assign micromatriz[19][31] = 9'b111111111;
assign micromatriz[19][32] = 9'b111111111;
assign micromatriz[19][33] = 9'b111111111;
assign micromatriz[19][34] = 9'b111111111;
assign micromatriz[19][35] = 9'b111111111;
assign micromatriz[19][36] = 9'b111111111;
assign micromatriz[19][37] = 9'b111111111;
assign micromatriz[19][38] = 9'b111111111;
assign micromatriz[19][39] = 9'b111111111;
assign micromatriz[19][40] = 9'b111111111;
assign micromatriz[19][41] = 9'b111111111;
assign micromatriz[19][42] = 9'b111111111;
assign micromatriz[19][43] = 9'b111111111;
assign micromatriz[19][44] = 9'b111111111;
assign micromatriz[19][45] = 9'b111111111;
assign micromatriz[19][46] = 9'b111111111;
assign micromatriz[19][47] = 9'b111111111;
assign micromatriz[19][48] = 9'b111111111;
assign micromatriz[19][49] = 9'b111111111;
assign micromatriz[19][50] = 9'b111111111;
assign micromatriz[19][51] = 9'b111111111;
assign micromatriz[19][52] = 9'b111111111;
assign micromatriz[19][53] = 9'b111111111;
assign micromatriz[19][54] = 9'b111111111;
assign micromatriz[19][55] = 9'b111111111;
assign micromatriz[19][56] = 9'b111111111;
assign micromatriz[19][57] = 9'b111111111;
assign micromatriz[19][58] = 9'b111111111;
assign micromatriz[19][59] = 9'b111111111;
assign micromatriz[19][60] = 9'b111111111;
assign micromatriz[19][61] = 9'b111111111;
assign micromatriz[19][62] = 9'b111111111;
assign micromatriz[19][63] = 9'b111111111;
assign micromatriz[19][64] = 9'b111111111;
assign micromatriz[19][65] = 9'b111111111;
assign micromatriz[19][66] = 9'b111111111;
assign micromatriz[19][67] = 9'b111111111;
assign micromatriz[19][68] = 9'b111111111;
assign micromatriz[19][69] = 9'b111111111;
assign micromatriz[19][70] = 9'b111111111;
assign micromatriz[19][71] = 9'b111111111;
assign micromatriz[19][72] = 9'b111111111;
assign micromatriz[19][73] = 9'b111111111;
assign micromatriz[19][74] = 9'b111111111;
assign micromatriz[19][75] = 9'b111111111;
assign micromatriz[19][76] = 9'b111111111;
assign micromatriz[19][77] = 9'b111111111;
assign micromatriz[19][78] = 9'b111111111;
assign micromatriz[19][79] = 9'b111111111;
assign micromatriz[19][80] = 9'b111111111;
assign micromatriz[19][81] = 9'b111111111;
assign micromatriz[19][82] = 9'b111111111;
assign micromatriz[19][83] = 9'b111111111;
assign micromatriz[19][84] = 9'b111111111;
assign micromatriz[19][85] = 9'b111111111;
assign micromatriz[19][86] = 9'b111111111;
assign micromatriz[19][87] = 9'b111111111;
assign micromatriz[19][88] = 9'b111111111;
assign micromatriz[19][89] = 9'b111111111;
assign micromatriz[19][90] = 9'b111111111;
assign micromatriz[19][91] = 9'b111111111;
assign micromatriz[19][92] = 9'b111111111;
assign micromatriz[19][93] = 9'b111111111;
assign micromatriz[19][94] = 9'b111111111;
assign micromatriz[19][95] = 9'b111111111;
assign micromatriz[19][96] = 9'b111111111;
assign micromatriz[19][97] = 9'b111111111;
assign micromatriz[19][98] = 9'b111111111;
assign micromatriz[19][99] = 9'b111111111;
assign micromatriz[20][0] = 9'b111111111;
assign micromatriz[20][1] = 9'b111111111;
assign micromatriz[20][2] = 9'b111111111;
assign micromatriz[20][3] = 9'b111111111;
assign micromatriz[20][4] = 9'b111111111;
assign micromatriz[20][5] = 9'b111111111;
assign micromatriz[20][6] = 9'b111111111;
assign micromatriz[20][7] = 9'b111111111;
assign micromatriz[20][8] = 9'b111111111;
assign micromatriz[20][9] = 9'b111111111;
assign micromatriz[20][10] = 9'b111111111;
assign micromatriz[20][11] = 9'b111111111;
assign micromatriz[20][12] = 9'b111111111;
assign micromatriz[20][13] = 9'b111111111;
assign micromatriz[20][14] = 9'b111111111;
assign micromatriz[20][15] = 9'b111111111;
assign micromatriz[20][16] = 9'b111111111;
assign micromatriz[20][17] = 9'b111111111;
assign micromatriz[20][18] = 9'b111111111;
assign micromatriz[20][19] = 9'b111111111;
assign micromatriz[20][20] = 9'b111111111;
assign micromatriz[20][21] = 9'b111111111;
assign micromatriz[20][22] = 9'b111111111;
assign micromatriz[20][23] = 9'b111111111;
assign micromatriz[20][24] = 9'b111111111;
assign micromatriz[20][25] = 9'b111111111;
assign micromatriz[20][26] = 9'b111111111;
assign micromatriz[20][27] = 9'b111111111;
assign micromatriz[20][28] = 9'b111111111;
assign micromatriz[20][29] = 9'b111111111;
assign micromatriz[20][30] = 9'b111111111;
assign micromatriz[20][31] = 9'b111111111;
assign micromatriz[20][32] = 9'b111111111;
assign micromatriz[20][33] = 9'b111111111;
assign micromatriz[20][34] = 9'b111111111;
assign micromatriz[20][35] = 9'b111111111;
assign micromatriz[20][36] = 9'b111111111;
assign micromatriz[20][37] = 9'b111111111;
assign micromatriz[20][38] = 9'b111111111;
assign micromatriz[20][39] = 9'b111111111;
assign micromatriz[20][40] = 9'b111111111;
assign micromatriz[20][41] = 9'b111111111;
assign micromatriz[20][42] = 9'b111111111;
assign micromatriz[20][43] = 9'b111111111;
assign micromatriz[20][44] = 9'b111111111;
assign micromatriz[20][45] = 9'b111111111;
assign micromatriz[20][46] = 9'b111111111;
assign micromatriz[20][47] = 9'b111111111;
assign micromatriz[20][48] = 9'b111111111;
assign micromatriz[20][49] = 9'b111111111;
assign micromatriz[20][50] = 9'b111111111;
assign micromatriz[20][51] = 9'b111111111;
assign micromatriz[20][52] = 9'b111111111;
assign micromatriz[20][53] = 9'b111111111;
assign micromatriz[20][54] = 9'b111111111;
assign micromatriz[20][55] = 9'b111111111;
assign micromatriz[20][56] = 9'b111111111;
assign micromatriz[20][57] = 9'b111111111;
assign micromatriz[20][58] = 9'b111111111;
assign micromatriz[20][59] = 9'b111111111;
assign micromatriz[20][60] = 9'b111111111;
assign micromatriz[20][61] = 9'b111111111;
assign micromatriz[20][62] = 9'b111111111;
assign micromatriz[20][63] = 9'b111111111;
assign micromatriz[20][64] = 9'b111111111;
assign micromatriz[20][65] = 9'b111111111;
assign micromatriz[20][66] = 9'b111111111;
assign micromatriz[20][67] = 9'b111111111;
assign micromatriz[20][68] = 9'b111111111;
assign micromatriz[20][69] = 9'b111111111;
assign micromatriz[20][70] = 9'b111111111;
assign micromatriz[20][71] = 9'b111111111;
assign micromatriz[20][72] = 9'b111111111;
assign micromatriz[20][73] = 9'b111111111;
assign micromatriz[20][74] = 9'b111111111;
assign micromatriz[20][75] = 9'b111111111;
assign micromatriz[20][76] = 9'b111111111;
assign micromatriz[20][77] = 9'b111111111;
assign micromatriz[20][78] = 9'b111111111;
assign micromatriz[20][79] = 9'b111111111;
assign micromatriz[20][80] = 9'b111111111;
assign micromatriz[20][81] = 9'b111111111;
assign micromatriz[20][82] = 9'b111111111;
assign micromatriz[20][83] = 9'b111111111;
assign micromatriz[20][84] = 9'b111111111;
assign micromatriz[20][85] = 9'b111111111;
assign micromatriz[20][86] = 9'b111111111;
assign micromatriz[20][87] = 9'b111111111;
assign micromatriz[20][88] = 9'b111111111;
assign micromatriz[20][89] = 9'b111111111;
assign micromatriz[20][90] = 9'b111111111;
assign micromatriz[20][91] = 9'b111111111;
assign micromatriz[20][92] = 9'b111111111;
assign micromatriz[20][93] = 9'b111111111;
assign micromatriz[20][94] = 9'b111111111;
assign micromatriz[20][95] = 9'b111111111;
assign micromatriz[20][96] = 9'b111111111;
assign micromatriz[20][97] = 9'b111111111;
assign micromatriz[20][98] = 9'b111111111;
assign micromatriz[20][99] = 9'b111111111;
assign micromatriz[21][0] = 9'b111111111;
assign micromatriz[21][1] = 9'b111111111;
assign micromatriz[21][2] = 9'b111111111;
assign micromatriz[21][3] = 9'b111111111;
assign micromatriz[21][4] = 9'b111111111;
assign micromatriz[21][5] = 9'b111111111;
assign micromatriz[21][6] = 9'b111111111;
assign micromatriz[21][7] = 9'b111111111;
assign micromatriz[21][8] = 9'b111111111;
assign micromatriz[21][9] = 9'b111111111;
assign micromatriz[21][10] = 9'b111111111;
assign micromatriz[21][11] = 9'b111111111;
assign micromatriz[21][12] = 9'b111111111;
assign micromatriz[21][13] = 9'b111111111;
assign micromatriz[21][14] = 9'b111111111;
assign micromatriz[21][15] = 9'b111111111;
assign micromatriz[21][16] = 9'b111111111;
assign micromatriz[21][17] = 9'b111111111;
assign micromatriz[21][18] = 9'b111111111;
assign micromatriz[21][19] = 9'b111111111;
assign micromatriz[21][20] = 9'b111111111;
assign micromatriz[21][21] = 9'b111111111;
assign micromatriz[21][22] = 9'b111111111;
assign micromatriz[21][23] = 9'b111111111;
assign micromatriz[21][24] = 9'b111111111;
assign micromatriz[21][25] = 9'b111111111;
assign micromatriz[21][26] = 9'b111111111;
assign micromatriz[21][27] = 9'b111111111;
assign micromatriz[21][28] = 9'b111111111;
assign micromatriz[21][29] = 9'b111111111;
assign micromatriz[21][30] = 9'b111111111;
assign micromatriz[21][31] = 9'b111111111;
assign micromatriz[21][32] = 9'b111111111;
assign micromatriz[21][33] = 9'b111111111;
assign micromatriz[21][34] = 9'b111111111;
assign micromatriz[21][35] = 9'b111111111;
assign micromatriz[21][36] = 9'b111111111;
assign micromatriz[21][37] = 9'b111111111;
assign micromatriz[21][38] = 9'b111111111;
assign micromatriz[21][39] = 9'b111111111;
assign micromatriz[21][40] = 9'b111111111;
assign micromatriz[21][41] = 9'b111111111;
assign micromatriz[21][42] = 9'b111111111;
assign micromatriz[21][43] = 9'b111111111;
assign micromatriz[21][44] = 9'b111111111;
assign micromatriz[21][45] = 9'b111111111;
assign micromatriz[21][46] = 9'b111111111;
assign micromatriz[21][47] = 9'b111111111;
assign micromatriz[21][48] = 9'b111111111;
assign micromatriz[21][49] = 9'b111111111;
assign micromatriz[21][50] = 9'b111111111;
assign micromatriz[21][51] = 9'b111111111;
assign micromatriz[21][52] = 9'b111111111;
assign micromatriz[21][53] = 9'b111111111;
assign micromatriz[21][54] = 9'b111111111;
assign micromatriz[21][55] = 9'b111111111;
assign micromatriz[21][56] = 9'b111111111;
assign micromatriz[21][57] = 9'b111111111;
assign micromatriz[21][58] = 9'b111111111;
assign micromatriz[21][59] = 9'b111111111;
assign micromatriz[21][60] = 9'b111111111;
assign micromatriz[21][61] = 9'b111111111;
assign micromatriz[21][62] = 9'b111111111;
assign micromatriz[21][63] = 9'b111111111;
assign micromatriz[21][64] = 9'b111111111;
assign micromatriz[21][65] = 9'b111111111;
assign micromatriz[21][66] = 9'b111111111;
assign micromatriz[21][67] = 9'b111111111;
assign micromatriz[21][68] = 9'b111111111;
assign micromatriz[21][69] = 9'b111111111;
assign micromatriz[21][70] = 9'b111111111;
assign micromatriz[21][71] = 9'b111111111;
assign micromatriz[21][72] = 9'b111111111;
assign micromatriz[21][73] = 9'b111111111;
assign micromatriz[21][74] = 9'b111111111;
assign micromatriz[21][75] = 9'b111111111;
assign micromatriz[21][76] = 9'b111111111;
assign micromatriz[21][77] = 9'b111111111;
assign micromatriz[21][78] = 9'b111111111;
assign micromatriz[21][79] = 9'b111111111;
assign micromatriz[21][80] = 9'b111111111;
assign micromatriz[21][81] = 9'b111111111;
assign micromatriz[21][82] = 9'b111111111;
assign micromatriz[21][83] = 9'b111111111;
assign micromatriz[21][84] = 9'b111111111;
assign micromatriz[21][85] = 9'b111111111;
assign micromatriz[21][86] = 9'b111111111;
assign micromatriz[21][87] = 9'b111111111;
assign micromatriz[21][88] = 9'b111111111;
assign micromatriz[21][89] = 9'b111111111;
assign micromatriz[21][90] = 9'b111111111;
assign micromatriz[21][91] = 9'b111111111;
assign micromatriz[21][92] = 9'b111111111;
assign micromatriz[21][93] = 9'b111111111;
assign micromatriz[21][94] = 9'b111111111;
assign micromatriz[21][95] = 9'b111111111;
assign micromatriz[21][96] = 9'b111111111;
assign micromatriz[21][97] = 9'b111111111;
assign micromatriz[21][98] = 9'b111111111;
assign micromatriz[21][99] = 9'b111111111;
assign micromatriz[22][0] = 9'b111111111;
assign micromatriz[22][1] = 9'b111111111;
assign micromatriz[22][2] = 9'b111111111;
assign micromatriz[22][3] = 9'b111111111;
assign micromatriz[22][4] = 9'b111111111;
assign micromatriz[22][5] = 9'b111111111;
assign micromatriz[22][6] = 9'b111111111;
assign micromatriz[22][7] = 9'b111111111;
assign micromatriz[22][8] = 9'b111111111;
assign micromatriz[22][9] = 9'b111111111;
assign micromatriz[22][10] = 9'b111111111;
assign micromatriz[22][11] = 9'b111111111;
assign micromatriz[22][12] = 9'b111111111;
assign micromatriz[22][13] = 9'b111111111;
assign micromatriz[22][14] = 9'b111111111;
assign micromatriz[22][15] = 9'b111111111;
assign micromatriz[22][16] = 9'b111111111;
assign micromatriz[22][17] = 9'b111111111;
assign micromatriz[22][18] = 9'b111111111;
assign micromatriz[22][19] = 9'b111111111;
assign micromatriz[22][20] = 9'b111111111;
assign micromatriz[22][21] = 9'b111111111;
assign micromatriz[22][22] = 9'b111111111;
assign micromatriz[22][23] = 9'b111111111;
assign micromatriz[22][24] = 9'b111111111;
assign micromatriz[22][25] = 9'b111111111;
assign micromatriz[22][26] = 9'b111111111;
assign micromatriz[22][27] = 9'b111111111;
assign micromatriz[22][28] = 9'b111111111;
assign micromatriz[22][29] = 9'b111111111;
assign micromatriz[22][30] = 9'b111111111;
assign micromatriz[22][31] = 9'b111111111;
assign micromatriz[22][32] = 9'b111111111;
assign micromatriz[22][33] = 9'b111111111;
assign micromatriz[22][34] = 9'b111111111;
assign micromatriz[22][35] = 9'b111111111;
assign micromatriz[22][36] = 9'b111111111;
assign micromatriz[22][37] = 9'b111111111;
assign micromatriz[22][38] = 9'b111111111;
assign micromatriz[22][39] = 9'b111111111;
assign micromatriz[22][40] = 9'b111111111;
assign micromatriz[22][41] = 9'b111111111;
assign micromatriz[22][42] = 9'b111111111;
assign micromatriz[22][43] = 9'b111111111;
assign micromatriz[22][44] = 9'b111111111;
assign micromatriz[22][45] = 9'b111111111;
assign micromatriz[22][46] = 9'b111111111;
assign micromatriz[22][47] = 9'b111111111;
assign micromatriz[22][48] = 9'b111111111;
assign micromatriz[22][49] = 9'b111111111;
assign micromatriz[22][50] = 9'b111111111;
assign micromatriz[22][51] = 9'b111111111;
assign micromatriz[22][52] = 9'b111111111;
assign micromatriz[22][53] = 9'b111111111;
assign micromatriz[22][54] = 9'b111111111;
assign micromatriz[22][55] = 9'b111111111;
assign micromatriz[22][56] = 9'b111111111;
assign micromatriz[22][57] = 9'b111111111;
assign micromatriz[22][58] = 9'b111111111;
assign micromatriz[22][59] = 9'b111111111;
assign micromatriz[22][60] = 9'b111111111;
assign micromatriz[22][61] = 9'b111111111;
assign micromatriz[22][62] = 9'b111111111;
assign micromatriz[22][63] = 9'b111111111;
assign micromatriz[22][64] = 9'b111111111;
assign micromatriz[22][65] = 9'b111111111;
assign micromatriz[22][66] = 9'b111111111;
assign micromatriz[22][67] = 9'b111111111;
assign micromatriz[22][68] = 9'b111111111;
assign micromatriz[22][69] = 9'b111111111;
assign micromatriz[22][70] = 9'b111111111;
assign micromatriz[22][71] = 9'b111111111;
assign micromatriz[22][72] = 9'b111111111;
assign micromatriz[22][73] = 9'b111111111;
assign micromatriz[22][74] = 9'b111111111;
assign micromatriz[22][75] = 9'b111111111;
assign micromatriz[22][76] = 9'b111111111;
assign micromatriz[22][77] = 9'b111111111;
assign micromatriz[22][78] = 9'b111111111;
assign micromatriz[22][79] = 9'b111111111;
assign micromatriz[22][80] = 9'b111111111;
assign micromatriz[22][81] = 9'b111111111;
assign micromatriz[22][82] = 9'b111111111;
assign micromatriz[22][83] = 9'b111111111;
assign micromatriz[22][84] = 9'b111111111;
assign micromatriz[22][85] = 9'b111111111;
assign micromatriz[22][86] = 9'b111111111;
assign micromatriz[22][87] = 9'b111111111;
assign micromatriz[22][88] = 9'b111111111;
assign micromatriz[22][89] = 9'b111111111;
assign micromatriz[22][90] = 9'b111111111;
assign micromatriz[22][91] = 9'b111111111;
assign micromatriz[22][92] = 9'b111111111;
assign micromatriz[22][93] = 9'b111111111;
assign micromatriz[22][94] = 9'b111111111;
assign micromatriz[22][95] = 9'b111111111;
assign micromatriz[22][96] = 9'b111111111;
assign micromatriz[22][97] = 9'b111111111;
assign micromatriz[22][98] = 9'b111111111;
assign micromatriz[22][99] = 9'b111111111;
assign micromatriz[23][0] = 9'b111111111;
assign micromatriz[23][1] = 9'b111111111;
assign micromatriz[23][2] = 9'b111111111;
assign micromatriz[23][3] = 9'b111111111;
assign micromatriz[23][4] = 9'b111111111;
assign micromatriz[23][5] = 9'b111111111;
assign micromatriz[23][6] = 9'b111111111;
assign micromatriz[23][7] = 9'b111111111;
assign micromatriz[23][8] = 9'b111111111;
assign micromatriz[23][9] = 9'b111111111;
assign micromatriz[23][10] = 9'b111111111;
assign micromatriz[23][11] = 9'b111111111;
assign micromatriz[23][12] = 9'b111111111;
assign micromatriz[23][13] = 9'b111111111;
assign micromatriz[23][14] = 9'b111111111;
assign micromatriz[23][15] = 9'b111111111;
assign micromatriz[23][16] = 9'b111111111;
assign micromatriz[23][17] = 9'b111111111;
assign micromatriz[23][18] = 9'b111111111;
assign micromatriz[23][19] = 9'b111111111;
assign micromatriz[23][20] = 9'b111111111;
assign micromatriz[23][21] = 9'b111111111;
assign micromatriz[23][22] = 9'b111111111;
assign micromatriz[23][23] = 9'b111111111;
assign micromatriz[23][24] = 9'b111111111;
assign micromatriz[23][25] = 9'b111111111;
assign micromatriz[23][26] = 9'b111111111;
assign micromatriz[23][27] = 9'b111111111;
assign micromatriz[23][28] = 9'b111111111;
assign micromatriz[23][29] = 9'b111111111;
assign micromatriz[23][30] = 9'b111111111;
assign micromatriz[23][31] = 9'b111111111;
assign micromatriz[23][32] = 9'b111111111;
assign micromatriz[23][33] = 9'b111111111;
assign micromatriz[23][34] = 9'b111111111;
assign micromatriz[23][35] = 9'b111111111;
assign micromatriz[23][36] = 9'b111111111;
assign micromatriz[23][37] = 9'b111111111;
assign micromatriz[23][38] = 9'b111111111;
assign micromatriz[23][39] = 9'b111111111;
assign micromatriz[23][40] = 9'b111111111;
assign micromatriz[23][41] = 9'b111111111;
assign micromatriz[23][42] = 9'b111111111;
assign micromatriz[23][43] = 9'b111111111;
assign micromatriz[23][44] = 9'b111111111;
assign micromatriz[23][45] = 9'b111111111;
assign micromatriz[23][46] = 9'b111111111;
assign micromatriz[23][47] = 9'b111111111;
assign micromatriz[23][48] = 9'b111111111;
assign micromatriz[23][49] = 9'b111111111;
assign micromatriz[23][50] = 9'b111111111;
assign micromatriz[23][51] = 9'b111111111;
assign micromatriz[23][52] = 9'b111111111;
assign micromatriz[23][53] = 9'b111111111;
assign micromatriz[23][54] = 9'b111111111;
assign micromatriz[23][55] = 9'b111111111;
assign micromatriz[23][56] = 9'b111111111;
assign micromatriz[23][57] = 9'b111111111;
assign micromatriz[23][58] = 9'b111111111;
assign micromatriz[23][59] = 9'b111111111;
assign micromatriz[23][60] = 9'b111111111;
assign micromatriz[23][61] = 9'b111111111;
assign micromatriz[23][62] = 9'b111111111;
assign micromatriz[23][63] = 9'b111111111;
assign micromatriz[23][64] = 9'b111111111;
assign micromatriz[23][65] = 9'b111111111;
assign micromatriz[23][66] = 9'b111111111;
assign micromatriz[23][67] = 9'b111111111;
assign micromatriz[23][68] = 9'b111111111;
assign micromatriz[23][69] = 9'b111111111;
assign micromatriz[23][70] = 9'b111111111;
assign micromatriz[23][71] = 9'b111111111;
assign micromatriz[23][72] = 9'b111111111;
assign micromatriz[23][73] = 9'b111111111;
assign micromatriz[23][74] = 9'b111111111;
assign micromatriz[23][75] = 9'b111111111;
assign micromatriz[23][76] = 9'b111111111;
assign micromatriz[23][77] = 9'b111111111;
assign micromatriz[23][78] = 9'b111111111;
assign micromatriz[23][79] = 9'b111111111;
assign micromatriz[23][80] = 9'b111111111;
assign micromatriz[23][81] = 9'b111111111;
assign micromatriz[23][82] = 9'b111111111;
assign micromatriz[23][83] = 9'b111111111;
assign micromatriz[23][84] = 9'b111111111;
assign micromatriz[23][85] = 9'b111111111;
assign micromatriz[23][86] = 9'b111111111;
assign micromatriz[23][87] = 9'b111111111;
assign micromatriz[23][88] = 9'b111111111;
assign micromatriz[23][89] = 9'b111111111;
assign micromatriz[23][90] = 9'b111111111;
assign micromatriz[23][91] = 9'b111111111;
assign micromatriz[23][92] = 9'b111111111;
assign micromatriz[23][93] = 9'b111111111;
assign micromatriz[23][94] = 9'b111111111;
assign micromatriz[23][95] = 9'b111111111;
assign micromatriz[23][96] = 9'b111111111;
assign micromatriz[23][97] = 9'b111111111;
assign micromatriz[23][98] = 9'b111111111;
assign micromatriz[23][99] = 9'b111111111;
assign micromatriz[24][0] = 9'b111111111;
assign micromatriz[24][1] = 9'b111111111;
assign micromatriz[24][2] = 9'b111111111;
assign micromatriz[24][3] = 9'b111111111;
assign micromatriz[24][4] = 9'b111111111;
assign micromatriz[24][5] = 9'b111111111;
assign micromatriz[24][6] = 9'b111111111;
assign micromatriz[24][7] = 9'b111111111;
assign micromatriz[24][8] = 9'b111111111;
assign micromatriz[24][9] = 9'b111111111;
assign micromatriz[24][10] = 9'b111111111;
assign micromatriz[24][11] = 9'b111111111;
assign micromatriz[24][12] = 9'b111111111;
assign micromatriz[24][13] = 9'b111111111;
assign micromatriz[24][14] = 9'b111111111;
assign micromatriz[24][15] = 9'b111111111;
assign micromatriz[24][16] = 9'b111111111;
assign micromatriz[24][17] = 9'b111111111;
assign micromatriz[24][18] = 9'b111111111;
assign micromatriz[24][19] = 9'b111111111;
assign micromatriz[24][20] = 9'b111111111;
assign micromatriz[24][21] = 9'b111111111;
assign micromatriz[24][22] = 9'b111111111;
assign micromatriz[24][23] = 9'b111111111;
assign micromatriz[24][24] = 9'b111111111;
assign micromatriz[24][25] = 9'b111111111;
assign micromatriz[24][26] = 9'b111111111;
assign micromatriz[24][27] = 9'b111111111;
assign micromatriz[24][28] = 9'b111111111;
assign micromatriz[24][29] = 9'b111111111;
assign micromatriz[24][30] = 9'b111111111;
assign micromatriz[24][31] = 9'b111111111;
assign micromatriz[24][32] = 9'b111111111;
assign micromatriz[24][33] = 9'b111111111;
assign micromatriz[24][34] = 9'b111111111;
assign micromatriz[24][35] = 9'b111111111;
assign micromatriz[24][36] = 9'b111111111;
assign micromatriz[24][37] = 9'b111111111;
assign micromatriz[24][38] = 9'b111111111;
assign micromatriz[24][39] = 9'b111111111;
assign micromatriz[24][40] = 9'b111111111;
assign micromatriz[24][41] = 9'b111111111;
assign micromatriz[24][42] = 9'b111111111;
assign micromatriz[24][43] = 9'b111111111;
assign micromatriz[24][44] = 9'b111111111;
assign micromatriz[24][45] = 9'b111111111;
assign micromatriz[24][46] = 9'b111111111;
assign micromatriz[24][47] = 9'b111111111;
assign micromatriz[24][48] = 9'b111111111;
assign micromatriz[24][49] = 9'b111111111;
assign micromatriz[24][50] = 9'b111111111;
assign micromatriz[24][51] = 9'b111111111;
assign micromatriz[24][52] = 9'b111111111;
assign micromatriz[24][53] = 9'b111111111;
assign micromatriz[24][54] = 9'b111111111;
assign micromatriz[24][55] = 9'b111111111;
assign micromatriz[24][56] = 9'b111111111;
assign micromatriz[24][57] = 9'b111111111;
assign micromatriz[24][58] = 9'b111111111;
assign micromatriz[24][59] = 9'b111111111;
assign micromatriz[24][60] = 9'b111111111;
assign micromatriz[24][61] = 9'b111111111;
assign micromatriz[24][62] = 9'b111111111;
assign micromatriz[24][63] = 9'b111111111;
assign micromatriz[24][64] = 9'b111111111;
assign micromatriz[24][65] = 9'b111111111;
assign micromatriz[24][66] = 9'b111111111;
assign micromatriz[24][67] = 9'b111111111;
assign micromatriz[24][68] = 9'b111111111;
assign micromatriz[24][69] = 9'b111111111;
assign micromatriz[24][70] = 9'b111111111;
assign micromatriz[24][71] = 9'b111111111;
assign micromatriz[24][72] = 9'b111111111;
assign micromatriz[24][73] = 9'b111111111;
assign micromatriz[24][74] = 9'b111111111;
assign micromatriz[24][75] = 9'b111111111;
assign micromatriz[24][76] = 9'b111111111;
assign micromatriz[24][77] = 9'b111111111;
assign micromatriz[24][78] = 9'b111111111;
assign micromatriz[24][79] = 9'b111111111;
assign micromatriz[24][80] = 9'b111111111;
assign micromatriz[24][81] = 9'b111111111;
assign micromatriz[24][82] = 9'b111111111;
assign micromatriz[24][83] = 9'b111111111;
assign micromatriz[24][84] = 9'b111111111;
assign micromatriz[24][85] = 9'b111111111;
assign micromatriz[24][86] = 9'b111111111;
assign micromatriz[24][87] = 9'b111111111;
assign micromatriz[24][88] = 9'b111111111;
assign micromatriz[24][89] = 9'b111111111;
assign micromatriz[24][90] = 9'b111111111;
assign micromatriz[24][91] = 9'b111111111;
assign micromatriz[24][92] = 9'b111111111;
assign micromatriz[24][93] = 9'b111111111;
assign micromatriz[24][94] = 9'b111111111;
assign micromatriz[24][95] = 9'b111111111;
assign micromatriz[24][96] = 9'b111111111;
assign micromatriz[24][97] = 9'b111111111;
assign micromatriz[24][98] = 9'b111111111;
assign micromatriz[24][99] = 9'b111111111;
assign micromatriz[25][0] = 9'b111111111;
assign micromatriz[25][1] = 9'b111111111;
assign micromatriz[25][2] = 9'b111111111;
assign micromatriz[25][3] = 9'b111111111;
assign micromatriz[25][4] = 9'b111111111;
assign micromatriz[25][5] = 9'b111111111;
assign micromatriz[25][6] = 9'b111111111;
assign micromatriz[25][7] = 9'b111111111;
assign micromatriz[25][8] = 9'b111111111;
assign micromatriz[25][9] = 9'b111111111;
assign micromatriz[25][10] = 9'b111111111;
assign micromatriz[25][11] = 9'b111111111;
assign micromatriz[25][12] = 9'b111111111;
assign micromatriz[25][13] = 9'b111111111;
assign micromatriz[25][14] = 9'b111111111;
assign micromatriz[25][15] = 9'b111111111;
assign micromatriz[25][16] = 9'b111111111;
assign micromatriz[25][17] = 9'b111111111;
assign micromatriz[25][18] = 9'b111111111;
assign micromatriz[25][19] = 9'b111111111;
assign micromatriz[25][20] = 9'b111111111;
assign micromatriz[25][21] = 9'b111111111;
assign micromatriz[25][22] = 9'b111111111;
assign micromatriz[25][23] = 9'b111111111;
assign micromatriz[25][24] = 9'b111111111;
assign micromatriz[25][25] = 9'b111111111;
assign micromatriz[25][26] = 9'b111111111;
assign micromatriz[25][27] = 9'b111111111;
assign micromatriz[25][28] = 9'b111111111;
assign micromatriz[25][29] = 9'b111111111;
assign micromatriz[25][30] = 9'b111111111;
assign micromatriz[25][31] = 9'b111111111;
assign micromatriz[25][32] = 9'b111111111;
assign micromatriz[25][33] = 9'b111111111;
assign micromatriz[25][34] = 9'b111111111;
assign micromatriz[25][35] = 9'b111111111;
assign micromatriz[25][36] = 9'b111111111;
assign micromatriz[25][37] = 9'b111111111;
assign micromatriz[25][38] = 9'b111111111;
assign micromatriz[25][39] = 9'b111111111;
assign micromatriz[25][40] = 9'b111111111;
assign micromatriz[25][41] = 9'b111111111;
assign micromatriz[25][42] = 9'b111111111;
assign micromatriz[25][43] = 9'b111111111;
assign micromatriz[25][44] = 9'b111111111;
assign micromatriz[25][45] = 9'b111111111;
assign micromatriz[25][46] = 9'b111111111;
assign micromatriz[25][47] = 9'b111111111;
assign micromatriz[25][48] = 9'b111111111;
assign micromatriz[25][49] = 9'b111111111;
assign micromatriz[25][50] = 9'b111111111;
assign micromatriz[25][51] = 9'b111111111;
assign micromatriz[25][52] = 9'b111111111;
assign micromatriz[25][53] = 9'b111111111;
assign micromatriz[25][54] = 9'b111111111;
assign micromatriz[25][55] = 9'b111111111;
assign micromatriz[25][56] = 9'b111111111;
assign micromatriz[25][57] = 9'b111111111;
assign micromatriz[25][58] = 9'b111111111;
assign micromatriz[25][59] = 9'b111111111;
assign micromatriz[25][60] = 9'b111111111;
assign micromatriz[25][61] = 9'b111111111;
assign micromatriz[25][62] = 9'b111111111;
assign micromatriz[25][63] = 9'b111111111;
assign micromatriz[25][64] = 9'b111111111;
assign micromatriz[25][65] = 9'b111111111;
assign micromatriz[25][66] = 9'b111111111;
assign micromatriz[25][67] = 9'b111111111;
assign micromatriz[25][68] = 9'b111111111;
assign micromatriz[25][69] = 9'b111111111;
assign micromatriz[25][70] = 9'b111111111;
assign micromatriz[25][71] = 9'b111111111;
assign micromatriz[25][72] = 9'b111111111;
assign micromatriz[25][73] = 9'b111111111;
assign micromatriz[25][74] = 9'b111111111;
assign micromatriz[25][75] = 9'b111111111;
assign micromatriz[25][76] = 9'b111111111;
assign micromatriz[25][77] = 9'b111111111;
assign micromatriz[25][78] = 9'b111111111;
assign micromatriz[25][79] = 9'b111111111;
assign micromatriz[25][80] = 9'b111111111;
assign micromatriz[25][81] = 9'b111111111;
assign micromatriz[25][82] = 9'b111111111;
assign micromatriz[25][83] = 9'b111111111;
assign micromatriz[25][84] = 9'b111111111;
assign micromatriz[25][85] = 9'b111111111;
assign micromatriz[25][86] = 9'b111111111;
assign micromatriz[25][87] = 9'b111111111;
assign micromatriz[25][88] = 9'b111111111;
assign micromatriz[25][89] = 9'b111111111;
assign micromatriz[25][90] = 9'b111111111;
assign micromatriz[25][91] = 9'b111111111;
assign micromatriz[25][92] = 9'b111111111;
assign micromatriz[25][93] = 9'b111111111;
assign micromatriz[25][94] = 9'b111111111;
assign micromatriz[25][95] = 9'b111111111;
assign micromatriz[25][96] = 9'b111111111;
assign micromatriz[25][97] = 9'b111111111;
assign micromatriz[25][98] = 9'b111111111;
assign micromatriz[25][99] = 9'b111111111;
assign micromatriz[26][0] = 9'b111111111;
assign micromatriz[26][1] = 9'b111111111;
assign micromatriz[26][2] = 9'b111111111;
assign micromatriz[26][3] = 9'b111111111;
assign micromatriz[26][4] = 9'b111111111;
assign micromatriz[26][5] = 9'b111111111;
assign micromatriz[26][6] = 9'b111111111;
assign micromatriz[26][7] = 9'b111111111;
assign micromatriz[26][8] = 9'b111111111;
assign micromatriz[26][9] = 9'b111111111;
assign micromatriz[26][10] = 9'b111111111;
assign micromatriz[26][11] = 9'b111111111;
assign micromatriz[26][12] = 9'b111111111;
assign micromatriz[26][13] = 9'b111111111;
assign micromatriz[26][14] = 9'b111111111;
assign micromatriz[26][15] = 9'b111111111;
assign micromatriz[26][16] = 9'b111111111;
assign micromatriz[26][17] = 9'b111111111;
assign micromatriz[26][18] = 9'b111111111;
assign micromatriz[26][19] = 9'b111111111;
assign micromatriz[26][20] = 9'b111111111;
assign micromatriz[26][21] = 9'b111111111;
assign micromatriz[26][22] = 9'b111111111;
assign micromatriz[26][23] = 9'b111111111;
assign micromatriz[26][24] = 9'b111111111;
assign micromatriz[26][25] = 9'b111111111;
assign micromatriz[26][26] = 9'b111111111;
assign micromatriz[26][27] = 9'b111111111;
assign micromatriz[26][28] = 9'b111111111;
assign micromatriz[26][29] = 9'b111111111;
assign micromatriz[26][30] = 9'b111111111;
assign micromatriz[26][31] = 9'b111111111;
assign micromatriz[26][32] = 9'b111111111;
assign micromatriz[26][33] = 9'b111111111;
assign micromatriz[26][34] = 9'b111111111;
assign micromatriz[26][35] = 9'b111111111;
assign micromatriz[26][36] = 9'b111111111;
assign micromatriz[26][37] = 9'b111111111;
assign micromatriz[26][38] = 9'b111111111;
assign micromatriz[26][39] = 9'b111111111;
assign micromatriz[26][40] = 9'b111111111;
assign micromatriz[26][41] = 9'b111111111;
assign micromatriz[26][42] = 9'b111111111;
assign micromatriz[26][43] = 9'b111111111;
assign micromatriz[26][44] = 9'b111111111;
assign micromatriz[26][45] = 9'b111111111;
assign micromatriz[26][46] = 9'b111111111;
assign micromatriz[26][47] = 9'b111111111;
assign micromatriz[26][48] = 9'b111111111;
assign micromatriz[26][49] = 9'b111111111;
assign micromatriz[26][50] = 9'b111111111;
assign micromatriz[26][51] = 9'b111111111;
assign micromatriz[26][52] = 9'b111111111;
assign micromatriz[26][53] = 9'b111111111;
assign micromatriz[26][54] = 9'b111111111;
assign micromatriz[26][55] = 9'b111111111;
assign micromatriz[26][56] = 9'b111111111;
assign micromatriz[26][57] = 9'b111111111;
assign micromatriz[26][58] = 9'b111111111;
assign micromatriz[26][59] = 9'b111111111;
assign micromatriz[26][60] = 9'b111111111;
assign micromatriz[26][61] = 9'b111111111;
assign micromatriz[26][62] = 9'b111111111;
assign micromatriz[26][63] = 9'b111111111;
assign micromatriz[26][64] = 9'b111111111;
assign micromatriz[26][65] = 9'b111111111;
assign micromatriz[26][66] = 9'b111111111;
assign micromatriz[26][67] = 9'b111111111;
assign micromatriz[26][68] = 9'b111111111;
assign micromatriz[26][69] = 9'b111111111;
assign micromatriz[26][70] = 9'b111111111;
assign micromatriz[26][71] = 9'b111111111;
assign micromatriz[26][72] = 9'b111111111;
assign micromatriz[26][73] = 9'b111111111;
assign micromatriz[26][74] = 9'b111111111;
assign micromatriz[26][75] = 9'b111111111;
assign micromatriz[26][76] = 9'b111111111;
assign micromatriz[26][77] = 9'b111111111;
assign micromatriz[26][78] = 9'b111111111;
assign micromatriz[26][79] = 9'b111111111;
assign micromatriz[26][80] = 9'b111111111;
assign micromatriz[26][81] = 9'b111111111;
assign micromatriz[26][82] = 9'b111111111;
assign micromatriz[26][83] = 9'b111111111;
assign micromatriz[26][84] = 9'b111111111;
assign micromatriz[26][85] = 9'b111111111;
assign micromatriz[26][86] = 9'b111111111;
assign micromatriz[26][87] = 9'b111111111;
assign micromatriz[26][88] = 9'b111111111;
assign micromatriz[26][89] = 9'b111111111;
assign micromatriz[26][90] = 9'b111111111;
assign micromatriz[26][91] = 9'b111111111;
assign micromatriz[26][92] = 9'b111111111;
assign micromatriz[26][93] = 9'b111111111;
assign micromatriz[26][94] = 9'b111111111;
assign micromatriz[26][95] = 9'b111111111;
assign micromatriz[26][96] = 9'b111111111;
assign micromatriz[26][97] = 9'b111111111;
assign micromatriz[26][98] = 9'b111111111;
assign micromatriz[26][99] = 9'b111111111;
assign micromatriz[27][0] = 9'b111111111;
assign micromatriz[27][1] = 9'b111111111;
assign micromatriz[27][2] = 9'b111111111;
assign micromatriz[27][3] = 9'b111111111;
assign micromatriz[27][4] = 9'b111111111;
assign micromatriz[27][5] = 9'b111111111;
assign micromatriz[27][6] = 9'b111111111;
assign micromatriz[27][7] = 9'b111111111;
assign micromatriz[27][8] = 9'b111111111;
assign micromatriz[27][9] = 9'b111111111;
assign micromatriz[27][10] = 9'b111111111;
assign micromatriz[27][11] = 9'b111111111;
assign micromatriz[27][12] = 9'b111111111;
assign micromatriz[27][13] = 9'b111111111;
assign micromatriz[27][14] = 9'b111111111;
assign micromatriz[27][15] = 9'b111111111;
assign micromatriz[27][16] = 9'b111111111;
assign micromatriz[27][17] = 9'b111111111;
assign micromatriz[27][18] = 9'b111111111;
assign micromatriz[27][19] = 9'b111111111;
assign micromatriz[27][20] = 9'b111111111;
assign micromatriz[27][21] = 9'b111111111;
assign micromatriz[27][22] = 9'b111111111;
assign micromatriz[27][23] = 9'b111111111;
assign micromatriz[27][24] = 9'b111111111;
assign micromatriz[27][25] = 9'b111111111;
assign micromatriz[27][26] = 9'b111111111;
assign micromatriz[27][27] = 9'b111111111;
assign micromatriz[27][28] = 9'b111111111;
assign micromatriz[27][29] = 9'b111111111;
assign micromatriz[27][30] = 9'b111111111;
assign micromatriz[27][31] = 9'b111111111;
assign micromatriz[27][32] = 9'b111111111;
assign micromatriz[27][33] = 9'b111111111;
assign micromatriz[27][34] = 9'b111111111;
assign micromatriz[27][35] = 9'b111111111;
assign micromatriz[27][36] = 9'b111111111;
assign micromatriz[27][37] = 9'b111111111;
assign micromatriz[27][38] = 9'b111111111;
assign micromatriz[27][39] = 9'b111111111;
assign micromatriz[27][40] = 9'b111111111;
assign micromatriz[27][41] = 9'b111111111;
assign micromatriz[27][42] = 9'b111111111;
assign micromatriz[27][43] = 9'b111111111;
assign micromatriz[27][44] = 9'b111111111;
assign micromatriz[27][45] = 9'b111111111;
assign micromatriz[27][46] = 9'b111111111;
assign micromatriz[27][47] = 9'b111111111;
assign micromatriz[27][48] = 9'b111111111;
assign micromatriz[27][49] = 9'b111111111;
assign micromatriz[27][50] = 9'b111111111;
assign micromatriz[27][51] = 9'b111111111;
assign micromatriz[27][52] = 9'b111111111;
assign micromatriz[27][53] = 9'b111111111;
assign micromatriz[27][54] = 9'b111111111;
assign micromatriz[27][55] = 9'b111111111;
assign micromatriz[27][56] = 9'b111111111;
assign micromatriz[27][57] = 9'b111111111;
assign micromatriz[27][58] = 9'b111111111;
assign micromatriz[27][59] = 9'b111111111;
assign micromatriz[27][60] = 9'b111111111;
assign micromatriz[27][61] = 9'b111111111;
assign micromatriz[27][62] = 9'b111111111;
assign micromatriz[27][63] = 9'b111111111;
assign micromatriz[27][64] = 9'b111111111;
assign micromatriz[27][65] = 9'b111111111;
assign micromatriz[27][66] = 9'b111111111;
assign micromatriz[27][67] = 9'b111111111;
assign micromatriz[27][68] = 9'b111111111;
assign micromatriz[27][69] = 9'b111111111;
assign micromatriz[27][70] = 9'b111111111;
assign micromatriz[27][71] = 9'b111111111;
assign micromatriz[27][72] = 9'b111111111;
assign micromatriz[27][73] = 9'b111111111;
assign micromatriz[27][74] = 9'b111111111;
assign micromatriz[27][75] = 9'b111111111;
assign micromatriz[27][76] = 9'b111111111;
assign micromatriz[27][77] = 9'b111111111;
assign micromatriz[27][78] = 9'b111111111;
assign micromatriz[27][79] = 9'b111111111;
assign micromatriz[27][80] = 9'b111111111;
assign micromatriz[27][81] = 9'b111111111;
assign micromatriz[27][82] = 9'b111111111;
assign micromatriz[27][83] = 9'b111111111;
assign micromatriz[27][84] = 9'b111111111;
assign micromatriz[27][85] = 9'b111111111;
assign micromatriz[27][86] = 9'b111111111;
assign micromatriz[27][87] = 9'b111111111;
assign micromatriz[27][88] = 9'b111111111;
assign micromatriz[27][89] = 9'b111111111;
assign micromatriz[27][90] = 9'b111111111;
assign micromatriz[27][91] = 9'b111111111;
assign micromatriz[27][92] = 9'b111111111;
assign micromatriz[27][93] = 9'b111111111;
assign micromatriz[27][94] = 9'b111111111;
assign micromatriz[27][95] = 9'b111111111;
assign micromatriz[27][96] = 9'b111111111;
assign micromatriz[27][97] = 9'b111111111;
assign micromatriz[27][98] = 9'b111111111;
assign micromatriz[27][99] = 9'b111111111;
assign micromatriz[28][0] = 9'b111111111;
assign micromatriz[28][1] = 9'b111111111;
assign micromatriz[28][2] = 9'b111111111;
assign micromatriz[28][3] = 9'b111111111;
assign micromatriz[28][4] = 9'b111111111;
assign micromatriz[28][5] = 9'b111111111;
assign micromatriz[28][6] = 9'b111111111;
assign micromatriz[28][7] = 9'b111111111;
assign micromatriz[28][8] = 9'b111111111;
assign micromatriz[28][9] = 9'b111111111;
assign micromatriz[28][10] = 9'b111111111;
assign micromatriz[28][11] = 9'b111111111;
assign micromatriz[28][12] = 9'b111111111;
assign micromatriz[28][13] = 9'b111111111;
assign micromatriz[28][14] = 9'b111111111;
assign micromatriz[28][15] = 9'b111111111;
assign micromatriz[28][16] = 9'b110110110;
assign micromatriz[28][17] = 9'b101101101;
assign micromatriz[28][18] = 9'b101101101;
assign micromatriz[28][19] = 9'b101101101;
assign micromatriz[28][20] = 9'b101101101;
assign micromatriz[28][21] = 9'b101101101;
assign micromatriz[28][22] = 9'b101101101;
assign micromatriz[28][23] = 9'b101101101;
assign micromatriz[28][24] = 9'b101101101;
assign micromatriz[28][25] = 9'b101101101;
assign micromatriz[28][26] = 9'b101101101;
assign micromatriz[28][27] = 9'b101101101;
assign micromatriz[28][28] = 9'b101101101;
assign micromatriz[28][29] = 9'b101101101;
assign micromatriz[28][30] = 9'b101101101;
assign micromatriz[28][31] = 9'b101101101;
assign micromatriz[28][32] = 9'b101101101;
assign micromatriz[28][33] = 9'b101101101;
assign micromatriz[28][34] = 9'b101101101;
assign micromatriz[28][35] = 9'b101101101;
assign micromatriz[28][36] = 9'b101101101;
assign micromatriz[28][37] = 9'b101101101;
assign micromatriz[28][38] = 9'b101101101;
assign micromatriz[28][39] = 9'b101101101;
assign micromatriz[28][40] = 9'b101101101;
assign micromatriz[28][41] = 9'b101101101;
assign micromatriz[28][42] = 9'b101101101;
assign micromatriz[28][43] = 9'b101101101;
assign micromatriz[28][44] = 9'b101101101;
assign micromatriz[28][45] = 9'b101101101;
assign micromatriz[28][46] = 9'b101101101;
assign micromatriz[28][47] = 9'b101101101;
assign micromatriz[28][48] = 9'b101101101;
assign micromatriz[28][49] = 9'b101101101;
assign micromatriz[28][50] = 9'b101101101;
assign micromatriz[28][51] = 9'b101101101;
assign micromatriz[28][52] = 9'b101101101;
assign micromatriz[28][53] = 9'b101101101;
assign micromatriz[28][54] = 9'b101101101;
assign micromatriz[28][55] = 9'b101101101;
assign micromatriz[28][56] = 9'b101101101;
assign micromatriz[28][57] = 9'b101101101;
assign micromatriz[28][58] = 9'b101101101;
assign micromatriz[28][59] = 9'b101101101;
assign micromatriz[28][60] = 9'b101101101;
assign micromatriz[28][61] = 9'b101101101;
assign micromatriz[28][62] = 9'b101101101;
assign micromatriz[28][63] = 9'b101101101;
assign micromatriz[28][64] = 9'b101101101;
assign micromatriz[28][65] = 9'b101101101;
assign micromatriz[28][66] = 9'b101101101;
assign micromatriz[28][67] = 9'b101101101;
assign micromatriz[28][68] = 9'b101101101;
assign micromatriz[28][69] = 9'b101101101;
assign micromatriz[28][70] = 9'b101101101;
assign micromatriz[28][71] = 9'b101101101;
assign micromatriz[28][72] = 9'b101101101;
assign micromatriz[28][73] = 9'b101101101;
assign micromatriz[28][74] = 9'b101101101;
assign micromatriz[28][75] = 9'b101101101;
assign micromatriz[28][76] = 9'b101101101;
assign micromatriz[28][77] = 9'b101101101;
assign micromatriz[28][78] = 9'b101101101;
assign micromatriz[28][79] = 9'b101101101;
assign micromatriz[28][80] = 9'b101101101;
assign micromatriz[28][81] = 9'b101101101;
assign micromatriz[28][82] = 9'b101101101;
assign micromatriz[28][83] = 9'b110110110;
assign micromatriz[28][84] = 9'b111111111;
assign micromatriz[28][85] = 9'b111111111;
assign micromatriz[28][86] = 9'b111111111;
assign micromatriz[28][87] = 9'b111111111;
assign micromatriz[28][88] = 9'b111111111;
assign micromatriz[28][89] = 9'b111111111;
assign micromatriz[28][90] = 9'b111111111;
assign micromatriz[28][91] = 9'b111111111;
assign micromatriz[28][92] = 9'b111111111;
assign micromatriz[28][93] = 9'b111111111;
assign micromatriz[28][94] = 9'b111111111;
assign micromatriz[28][95] = 9'b111111111;
assign micromatriz[28][96] = 9'b111111111;
assign micromatriz[28][97] = 9'b111111111;
assign micromatriz[28][98] = 9'b111111111;
assign micromatriz[28][99] = 9'b111111111;
assign micromatriz[29][0] = 9'b111111111;
assign micromatriz[29][1] = 9'b111111111;
assign micromatriz[29][2] = 9'b111111111;
assign micromatriz[29][3] = 9'b111111111;
assign micromatriz[29][4] = 9'b111111111;
assign micromatriz[29][5] = 9'b111111111;
assign micromatriz[29][6] = 9'b111111111;
assign micromatriz[29][7] = 9'b111111111;
assign micromatriz[29][8] = 9'b111111111;
assign micromatriz[29][9] = 9'b111111111;
assign micromatriz[29][10] = 9'b111111111;
assign micromatriz[29][11] = 9'b111111111;
assign micromatriz[29][12] = 9'b111111111;
assign micromatriz[29][13] = 9'b111111111;
assign micromatriz[29][14] = 9'b111111111;
assign micromatriz[29][15] = 9'b111111111;
assign micromatriz[29][16] = 9'b101101101;
assign micromatriz[29][17] = 9'b100000000;
assign micromatriz[29][18] = 9'b100000000;
assign micromatriz[29][19] = 9'b100000000;
assign micromatriz[29][20] = 9'b100000000;
assign micromatriz[29][21] = 9'b100000000;
assign micromatriz[29][22] = 9'b100000000;
assign micromatriz[29][23] = 9'b100000000;
assign micromatriz[29][24] = 9'b100000000;
assign micromatriz[29][25] = 9'b100000000;
assign micromatriz[29][26] = 9'b100000000;
assign micromatriz[29][27] = 9'b100000000;
assign micromatriz[29][28] = 9'b100000000;
assign micromatriz[29][29] = 9'b100000000;
assign micromatriz[29][30] = 9'b100000000;
assign micromatriz[29][31] = 9'b100000000;
assign micromatriz[29][32] = 9'b100000000;
assign micromatriz[29][33] = 9'b100000000;
assign micromatriz[29][34] = 9'b100000000;
assign micromatriz[29][35] = 9'b100000000;
assign micromatriz[29][36] = 9'b100000000;
assign micromatriz[29][37] = 9'b100000000;
assign micromatriz[29][38] = 9'b100000000;
assign micromatriz[29][39] = 9'b100000000;
assign micromatriz[29][40] = 9'b100000000;
assign micromatriz[29][41] = 9'b100000000;
assign micromatriz[29][42] = 9'b100000000;
assign micromatriz[29][43] = 9'b100000000;
assign micromatriz[29][44] = 9'b100000000;
assign micromatriz[29][45] = 9'b100000000;
assign micromatriz[29][46] = 9'b100000000;
assign micromatriz[29][47] = 9'b100000000;
assign micromatriz[29][48] = 9'b100000000;
assign micromatriz[29][49] = 9'b100000000;
assign micromatriz[29][50] = 9'b100000000;
assign micromatriz[29][51] = 9'b100000000;
assign micromatriz[29][52] = 9'b100000000;
assign micromatriz[29][53] = 9'b100000000;
assign micromatriz[29][54] = 9'b100000000;
assign micromatriz[29][55] = 9'b100000000;
assign micromatriz[29][56] = 9'b100000000;
assign micromatriz[29][57] = 9'b100000000;
assign micromatriz[29][58] = 9'b100000000;
assign micromatriz[29][59] = 9'b100000000;
assign micromatriz[29][60] = 9'b100000000;
assign micromatriz[29][61] = 9'b100000000;
assign micromatriz[29][62] = 9'b100000000;
assign micromatriz[29][63] = 9'b100000000;
assign micromatriz[29][64] = 9'b100000000;
assign micromatriz[29][65] = 9'b100000000;
assign micromatriz[29][66] = 9'b100000000;
assign micromatriz[29][67] = 9'b100000000;
assign micromatriz[29][68] = 9'b100000000;
assign micromatriz[29][69] = 9'b100000000;
assign micromatriz[29][70] = 9'b100000000;
assign micromatriz[29][71] = 9'b100000000;
assign micromatriz[29][72] = 9'b100000000;
assign micromatriz[29][73] = 9'b100000000;
assign micromatriz[29][74] = 9'b100000000;
assign micromatriz[29][75] = 9'b100000000;
assign micromatriz[29][76] = 9'b100000000;
assign micromatriz[29][77] = 9'b100000000;
assign micromatriz[29][78] = 9'b100000000;
assign micromatriz[29][79] = 9'b100000000;
assign micromatriz[29][80] = 9'b100000000;
assign micromatriz[29][81] = 9'b100000000;
assign micromatriz[29][82] = 9'b100000000;
assign micromatriz[29][83] = 9'b101101101;
assign micromatriz[29][84] = 9'b111111111;
assign micromatriz[29][85] = 9'b111111111;
assign micromatriz[29][86] = 9'b111111111;
assign micromatriz[29][87] = 9'b111111111;
assign micromatriz[29][88] = 9'b111111111;
assign micromatriz[29][89] = 9'b111111111;
assign micromatriz[29][90] = 9'b111111111;
assign micromatriz[29][91] = 9'b111111111;
assign micromatriz[29][92] = 9'b111111111;
assign micromatriz[29][93] = 9'b111111111;
assign micromatriz[29][94] = 9'b111111111;
assign micromatriz[29][95] = 9'b111111111;
assign micromatriz[29][96] = 9'b111111111;
assign micromatriz[29][97] = 9'b111111111;
assign micromatriz[29][98] = 9'b111111111;
assign micromatriz[29][99] = 9'b111111111;
assign micromatriz[30][0] = 9'b111111111;
assign micromatriz[30][1] = 9'b111111111;
assign micromatriz[30][2] = 9'b111111111;
assign micromatriz[30][3] = 9'b111111111;
assign micromatriz[30][4] = 9'b111111111;
assign micromatriz[30][5] = 9'b111111111;
assign micromatriz[30][6] = 9'b111111111;
assign micromatriz[30][7] = 9'b111111111;
assign micromatriz[30][8] = 9'b111111111;
assign micromatriz[30][9] = 9'b111111111;
assign micromatriz[30][10] = 9'b111111111;
assign micromatriz[30][11] = 9'b111111111;
assign micromatriz[30][12] = 9'b111111111;
assign micromatriz[30][13] = 9'b111111111;
assign micromatriz[30][14] = 9'b111111111;
assign micromatriz[30][15] = 9'b111111111;
assign micromatriz[30][16] = 9'b101101101;
assign micromatriz[30][17] = 9'b100100100;
assign micromatriz[30][18] = 9'b100100100;
assign micromatriz[30][19] = 9'b100100100;
assign micromatriz[30][20] = 9'b100100100;
assign micromatriz[30][21] = 9'b100100100;
assign micromatriz[30][22] = 9'b100100100;
assign micromatriz[30][23] = 9'b100100100;
assign micromatriz[30][24] = 9'b100100100;
assign micromatriz[30][25] = 9'b100100100;
assign micromatriz[30][26] = 9'b100100100;
assign micromatriz[30][27] = 9'b100100100;
assign micromatriz[30][28] = 9'b100100100;
assign micromatriz[30][29] = 9'b100100100;
assign micromatriz[30][30] = 9'b100100100;
assign micromatriz[30][31] = 9'b100100100;
assign micromatriz[30][32] = 9'b100100100;
assign micromatriz[30][33] = 9'b100100100;
assign micromatriz[30][34] = 9'b100100100;
assign micromatriz[30][35] = 9'b100100100;
assign micromatriz[30][36] = 9'b100100100;
assign micromatriz[30][37] = 9'b100100100;
assign micromatriz[30][38] = 9'b100100100;
assign micromatriz[30][39] = 9'b100100100;
assign micromatriz[30][40] = 9'b100100100;
assign micromatriz[30][41] = 9'b100100100;
assign micromatriz[30][42] = 9'b100100100;
assign micromatriz[30][43] = 9'b100100100;
assign micromatriz[30][44] = 9'b100100100;
assign micromatriz[30][45] = 9'b100100100;
assign micromatriz[30][46] = 9'b100100100;
assign micromatriz[30][47] = 9'b100100100;
assign micromatriz[30][48] = 9'b100100100;
assign micromatriz[30][49] = 9'b100100100;
assign micromatriz[30][50] = 9'b100100100;
assign micromatriz[30][51] = 9'b100100100;
assign micromatriz[30][52] = 9'b100100100;
assign micromatriz[30][53] = 9'b100100100;
assign micromatriz[30][54] = 9'b100100100;
assign micromatriz[30][55] = 9'b100100100;
assign micromatriz[30][56] = 9'b100100100;
assign micromatriz[30][57] = 9'b100100100;
assign micromatriz[30][58] = 9'b100100100;
assign micromatriz[30][59] = 9'b100100100;
assign micromatriz[30][60] = 9'b100100100;
assign micromatriz[30][61] = 9'b100100100;
assign micromatriz[30][62] = 9'b100100100;
assign micromatriz[30][63] = 9'b100100100;
assign micromatriz[30][64] = 9'b100100100;
assign micromatriz[30][65] = 9'b100100100;
assign micromatriz[30][66] = 9'b100000000;
assign micromatriz[30][67] = 9'b100000000;
assign micromatriz[30][68] = 9'b100000000;
assign micromatriz[30][69] = 9'b100100100;
assign micromatriz[30][70] = 9'b100100100;
assign micromatriz[30][71] = 9'b100100100;
assign micromatriz[30][72] = 9'b100100100;
assign micromatriz[30][73] = 9'b100100100;
assign micromatriz[30][74] = 9'b100100100;
assign micromatriz[30][75] = 9'b100100100;
assign micromatriz[30][76] = 9'b100100100;
assign micromatriz[30][77] = 9'b100100100;
assign micromatriz[30][78] = 9'b100100100;
assign micromatriz[30][79] = 9'b100100100;
assign micromatriz[30][80] = 9'b100100100;
assign micromatriz[30][81] = 9'b100100100;
assign micromatriz[30][82] = 9'b100100100;
assign micromatriz[30][83] = 9'b101101101;
assign micromatriz[30][84] = 9'b111111111;
assign micromatriz[30][85] = 9'b111111111;
assign micromatriz[30][86] = 9'b111111111;
assign micromatriz[30][87] = 9'b111111111;
assign micromatriz[30][88] = 9'b111111111;
assign micromatriz[30][89] = 9'b111111111;
assign micromatriz[30][90] = 9'b111111111;
assign micromatriz[30][91] = 9'b111111111;
assign micromatriz[30][92] = 9'b111111111;
assign micromatriz[30][93] = 9'b111111111;
assign micromatriz[30][94] = 9'b111111111;
assign micromatriz[30][95] = 9'b111111111;
assign micromatriz[30][96] = 9'b111111111;
assign micromatriz[30][97] = 9'b111111111;
assign micromatriz[30][98] = 9'b111111111;
assign micromatriz[30][99] = 9'b111111111;
assign micromatriz[31][0] = 9'b111111111;
assign micromatriz[31][1] = 9'b111111111;
assign micromatriz[31][2] = 9'b111111111;
assign micromatriz[31][3] = 9'b111111111;
assign micromatriz[31][4] = 9'b111111111;
assign micromatriz[31][5] = 9'b111111111;
assign micromatriz[31][6] = 9'b111111111;
assign micromatriz[31][7] = 9'b111111111;
assign micromatriz[31][8] = 9'b111111111;
assign micromatriz[31][9] = 9'b111111111;
assign micromatriz[31][10] = 9'b111111111;
assign micromatriz[31][11] = 9'b111111111;
assign micromatriz[31][12] = 9'b111111111;
assign micromatriz[31][13] = 9'b111111111;
assign micromatriz[31][14] = 9'b100100100;
assign micromatriz[31][15] = 9'b100000000;
assign micromatriz[31][16] = 9'b101101101;
assign micromatriz[31][17] = 9'b111111111;
assign micromatriz[31][18] = 9'b111111111;
assign micromatriz[31][19] = 9'b111111111;
assign micromatriz[31][20] = 9'b111111111;
assign micromatriz[31][21] = 9'b111111111;
assign micromatriz[31][22] = 9'b111111111;
assign micromatriz[31][23] = 9'b111111111;
assign micromatriz[31][24] = 9'b111111111;
assign micromatriz[31][25] = 9'b111111111;
assign micromatriz[31][26] = 9'b111111111;
assign micromatriz[31][27] = 9'b111111111;
assign micromatriz[31][28] = 9'b111111111;
assign micromatriz[31][29] = 9'b111111111;
assign micromatriz[31][30] = 9'b111111111;
assign micromatriz[31][31] = 9'b111111111;
assign micromatriz[31][32] = 9'b111111111;
assign micromatriz[31][33] = 9'b111111111;
assign micromatriz[31][34] = 9'b111111111;
assign micromatriz[31][35] = 9'b111111111;
assign micromatriz[31][36] = 9'b111111111;
assign micromatriz[31][37] = 9'b111111111;
assign micromatriz[31][38] = 9'b111111111;
assign micromatriz[31][39] = 9'b111111111;
assign micromatriz[31][40] = 9'b111111111;
assign micromatriz[31][41] = 9'b111111111;
assign micromatriz[31][42] = 9'b111111111;
assign micromatriz[31][43] = 9'b111111111;
assign micromatriz[31][44] = 9'b111111111;
assign micromatriz[31][45] = 9'b111111111;
assign micromatriz[31][46] = 9'b111111111;
assign micromatriz[31][47] = 9'b111111111;
assign micromatriz[31][48] = 9'b111111111;
assign micromatriz[31][49] = 9'b111111111;
assign micromatriz[31][50] = 9'b111111111;
assign micromatriz[31][51] = 9'b111111111;
assign micromatriz[31][52] = 9'b111111111;
assign micromatriz[31][53] = 9'b111111111;
assign micromatriz[31][54] = 9'b111111111;
assign micromatriz[31][55] = 9'b111111111;
assign micromatriz[31][56] = 9'b111111111;
assign micromatriz[31][57] = 9'b111111111;
assign micromatriz[31][58] = 9'b111111111;
assign micromatriz[31][59] = 9'b111111111;
assign micromatriz[31][60] = 9'b111111111;
assign micromatriz[31][61] = 9'b111111111;
assign micromatriz[31][62] = 9'b111111111;
assign micromatriz[31][63] = 9'b111111111;
assign micromatriz[31][64] = 9'b111111111;
assign micromatriz[31][65] = 9'b111111111;
assign micromatriz[31][66] = 9'b110010010;
assign micromatriz[31][67] = 9'b100000000;
assign micromatriz[31][68] = 9'b100000000;
assign micromatriz[31][69] = 9'b111111111;
assign micromatriz[31][70] = 9'b111111111;
assign micromatriz[31][71] = 9'b111111111;
assign micromatriz[31][72] = 9'b111111111;
assign micromatriz[31][73] = 9'b111111111;
assign micromatriz[31][74] = 9'b111111111;
assign micromatriz[31][75] = 9'b111111111;
assign micromatriz[31][76] = 9'b111111111;
assign micromatriz[31][77] = 9'b111111111;
assign micromatriz[31][78] = 9'b111111111;
assign micromatriz[31][79] = 9'b111111111;
assign micromatriz[31][80] = 9'b111111111;
assign micromatriz[31][81] = 9'b111111111;
assign micromatriz[31][82] = 9'b111111111;
assign micromatriz[31][83] = 9'b101101101;
assign micromatriz[31][84] = 9'b100000000;
assign micromatriz[31][85] = 9'b100100100;
assign micromatriz[31][86] = 9'b111111111;
assign micromatriz[31][87] = 9'b111111111;
assign micromatriz[31][88] = 9'b111111111;
assign micromatriz[31][89] = 9'b111111111;
assign micromatriz[31][90] = 9'b111111111;
assign micromatriz[31][91] = 9'b111111111;
assign micromatriz[31][92] = 9'b111111111;
assign micromatriz[31][93] = 9'b111111111;
assign micromatriz[31][94] = 9'b111111111;
assign micromatriz[31][95] = 9'b111111111;
assign micromatriz[31][96] = 9'b111111111;
assign micromatriz[31][97] = 9'b111111111;
assign micromatriz[31][98] = 9'b111111111;
assign micromatriz[31][99] = 9'b111111111;
assign micromatriz[32][0] = 9'b111111111;
assign micromatriz[32][1] = 9'b111111111;
assign micromatriz[32][2] = 9'b111111111;
assign micromatriz[32][3] = 9'b111111111;
assign micromatriz[32][4] = 9'b111111111;
assign micromatriz[32][5] = 9'b111111111;
assign micromatriz[32][6] = 9'b111111111;
assign micromatriz[32][7] = 9'b111111111;
assign micromatriz[32][8] = 9'b111111111;
assign micromatriz[32][9] = 9'b111111111;
assign micromatriz[32][10] = 9'b111111111;
assign micromatriz[32][11] = 9'b111111111;
assign micromatriz[32][12] = 9'b111111111;
assign micromatriz[32][13] = 9'b111111111;
assign micromatriz[32][14] = 9'b100100100;
assign micromatriz[32][15] = 9'b100000000;
assign micromatriz[32][16] = 9'b101101101;
assign micromatriz[32][17] = 9'b111111111;
assign micromatriz[32][18] = 9'b111111111;
assign micromatriz[32][19] = 9'b111111111;
assign micromatriz[32][20] = 9'b111111111;
assign micromatriz[32][21] = 9'b111111111;
assign micromatriz[32][22] = 9'b111111111;
assign micromatriz[32][23] = 9'b111111111;
assign micromatriz[32][24] = 9'b111111111;
assign micromatriz[32][25] = 9'b111111111;
assign micromatriz[32][26] = 9'b111111111;
assign micromatriz[32][27] = 9'b111111111;
assign micromatriz[32][28] = 9'b111111111;
assign micromatriz[32][29] = 9'b111111111;
assign micromatriz[32][30] = 9'b111111111;
assign micromatriz[32][31] = 9'b111111111;
assign micromatriz[32][32] = 9'b111111111;
assign micromatriz[32][33] = 9'b111111111;
assign micromatriz[32][34] = 9'b111111111;
assign micromatriz[32][35] = 9'b111111111;
assign micromatriz[32][36] = 9'b111111111;
assign micromatriz[32][37] = 9'b111111111;
assign micromatriz[32][38] = 9'b111111111;
assign micromatriz[32][39] = 9'b111111111;
assign micromatriz[32][40] = 9'b111111111;
assign micromatriz[32][41] = 9'b111111111;
assign micromatriz[32][42] = 9'b111111111;
assign micromatriz[32][43] = 9'b111111111;
assign micromatriz[32][44] = 9'b111111111;
assign micromatriz[32][45] = 9'b111111111;
assign micromatriz[32][46] = 9'b111111111;
assign micromatriz[32][47] = 9'b111111111;
assign micromatriz[32][48] = 9'b111111111;
assign micromatriz[32][49] = 9'b111111111;
assign micromatriz[32][50] = 9'b111111111;
assign micromatriz[32][51] = 9'b111111111;
assign micromatriz[32][52] = 9'b111111111;
assign micromatriz[32][53] = 9'b111111111;
assign micromatriz[32][54] = 9'b111111111;
assign micromatriz[32][55] = 9'b111111111;
assign micromatriz[32][56] = 9'b111111111;
assign micromatriz[32][57] = 9'b111111111;
assign micromatriz[32][58] = 9'b111111111;
assign micromatriz[32][59] = 9'b111111111;
assign micromatriz[32][60] = 9'b111111111;
assign micromatriz[32][61] = 9'b111111111;
assign micromatriz[32][62] = 9'b111111111;
assign micromatriz[32][63] = 9'b111111111;
assign micromatriz[32][64] = 9'b111111111;
assign micromatriz[32][65] = 9'b111111111;
assign micromatriz[32][66] = 9'b110010010;
assign micromatriz[32][67] = 9'b100000000;
assign micromatriz[32][68] = 9'b100000000;
assign micromatriz[32][69] = 9'b111111111;
assign micromatriz[32][70] = 9'b111111111;
assign micromatriz[32][71] = 9'b111111111;
assign micromatriz[32][72] = 9'b111111111;
assign micromatriz[32][73] = 9'b111111111;
assign micromatriz[32][74] = 9'b111111111;
assign micromatriz[32][75] = 9'b111111111;
assign micromatriz[32][76] = 9'b111111111;
assign micromatriz[32][77] = 9'b111111111;
assign micromatriz[32][78] = 9'b111111111;
assign micromatriz[32][79] = 9'b111111111;
assign micromatriz[32][80] = 9'b111111111;
assign micromatriz[32][81] = 9'b111111111;
assign micromatriz[32][82] = 9'b111111111;
assign micromatriz[32][83] = 9'b101001101;
assign micromatriz[32][84] = 9'b100000000;
assign micromatriz[32][85] = 9'b100100100;
assign micromatriz[32][86] = 9'b111111111;
assign micromatriz[32][87] = 9'b111111111;
assign micromatriz[32][88] = 9'b111111111;
assign micromatriz[32][89] = 9'b111111111;
assign micromatriz[32][90] = 9'b111111111;
assign micromatriz[32][91] = 9'b111111111;
assign micromatriz[32][92] = 9'b111111111;
assign micromatriz[32][93] = 9'b111111111;
assign micromatriz[32][94] = 9'b111111111;
assign micromatriz[32][95] = 9'b111111111;
assign micromatriz[32][96] = 9'b111111111;
assign micromatriz[32][97] = 9'b111111111;
assign micromatriz[32][98] = 9'b111111111;
assign micromatriz[32][99] = 9'b111111111;
assign micromatriz[33][0] = 9'b111111111;
assign micromatriz[33][1] = 9'b111111111;
assign micromatriz[33][2] = 9'b111111111;
assign micromatriz[33][3] = 9'b111111111;
assign micromatriz[33][4] = 9'b111111111;
assign micromatriz[33][5] = 9'b111111111;
assign micromatriz[33][6] = 9'b111111111;
assign micromatriz[33][7] = 9'b111111111;
assign micromatriz[33][8] = 9'b111111111;
assign micromatriz[33][9] = 9'b111111111;
assign micromatriz[33][10] = 9'b111111111;
assign micromatriz[33][11] = 9'b111111111;
assign micromatriz[33][12] = 9'b111111111;
assign micromatriz[33][13] = 9'b111111111;
assign micromatriz[33][14] = 9'b100100100;
assign micromatriz[33][15] = 9'b100000000;
assign micromatriz[33][16] = 9'b101101101;
assign micromatriz[33][17] = 9'b111111111;
assign micromatriz[33][18] = 9'b111111111;
assign micromatriz[33][19] = 9'b111111111;
assign micromatriz[33][20] = 9'b111111111;
assign micromatriz[33][21] = 9'b111111111;
assign micromatriz[33][22] = 9'b111111111;
assign micromatriz[33][23] = 9'b111111111;
assign micromatriz[33][24] = 9'b111111111;
assign micromatriz[33][25] = 9'b111111111;
assign micromatriz[33][26] = 9'b111111111;
assign micromatriz[33][27] = 9'b111111111;
assign micromatriz[33][28] = 9'b111111111;
assign micromatriz[33][29] = 9'b111111111;
assign micromatriz[33][30] = 9'b111111111;
assign micromatriz[33][31] = 9'b111111111;
assign micromatriz[33][32] = 9'b111111111;
assign micromatriz[33][33] = 9'b111111111;
assign micromatriz[33][34] = 9'b111111111;
assign micromatriz[33][35] = 9'b111111111;
assign micromatriz[33][36] = 9'b111111111;
assign micromatriz[33][37] = 9'b111111111;
assign micromatriz[33][38] = 9'b111111111;
assign micromatriz[33][39] = 9'b111111111;
assign micromatriz[33][40] = 9'b111111111;
assign micromatriz[33][41] = 9'b111111111;
assign micromatriz[33][42] = 9'b111111111;
assign micromatriz[33][43] = 9'b111111111;
assign micromatriz[33][44] = 9'b111111111;
assign micromatriz[33][45] = 9'b111111111;
assign micromatriz[33][46] = 9'b111111111;
assign micromatriz[33][47] = 9'b111111111;
assign micromatriz[33][48] = 9'b111111111;
assign micromatriz[33][49] = 9'b111111111;
assign micromatriz[33][50] = 9'b111111111;
assign micromatriz[33][51] = 9'b111111111;
assign micromatriz[33][52] = 9'b111111111;
assign micromatriz[33][53] = 9'b111111111;
assign micromatriz[33][54] = 9'b111111111;
assign micromatriz[33][55] = 9'b111111111;
assign micromatriz[33][56] = 9'b111111111;
assign micromatriz[33][57] = 9'b111111111;
assign micromatriz[33][58] = 9'b111111111;
assign micromatriz[33][59] = 9'b111111111;
assign micromatriz[33][60] = 9'b111111111;
assign micromatriz[33][61] = 9'b111111111;
assign micromatriz[33][62] = 9'b111111111;
assign micromatriz[33][63] = 9'b111111111;
assign micromatriz[33][64] = 9'b110111111;
assign micromatriz[33][65] = 9'b110111111;
assign micromatriz[33][66] = 9'b101110001;
assign micromatriz[33][67] = 9'b100000000;
assign micromatriz[33][68] = 9'b100000000;
assign micromatriz[33][69] = 9'b111111111;
assign micromatriz[33][70] = 9'b111111111;
assign micromatriz[33][71] = 9'b111111111;
assign micromatriz[33][72] = 9'b111111111;
assign micromatriz[33][73] = 9'b110111111;
assign micromatriz[33][74] = 9'b101001001;
assign micromatriz[33][75] = 9'b101001000;
assign micromatriz[33][76] = 9'b101001000;
assign micromatriz[33][77] = 9'b100101000;
assign micromatriz[33][78] = 9'b101101101;
assign micromatriz[33][79] = 9'b111111111;
assign micromatriz[33][80] = 9'b111111111;
assign micromatriz[33][81] = 9'b110110111;
assign micromatriz[33][82] = 9'b111111111;
assign micromatriz[33][83] = 9'b101001001;
assign micromatriz[33][84] = 9'b100000000;
assign micromatriz[33][85] = 9'b100100100;
assign micromatriz[33][86] = 9'b111111111;
assign micromatriz[33][87] = 9'b111111111;
assign micromatriz[33][88] = 9'b111111111;
assign micromatriz[33][89] = 9'b111111111;
assign micromatriz[33][90] = 9'b111111111;
assign micromatriz[33][91] = 9'b111111111;
assign micromatriz[33][92] = 9'b111111111;
assign micromatriz[33][93] = 9'b111111111;
assign micromatriz[33][94] = 9'b111111111;
assign micromatriz[33][95] = 9'b111111111;
assign micromatriz[33][96] = 9'b111111111;
assign micromatriz[33][97] = 9'b111111111;
assign micromatriz[33][98] = 9'b111111111;
assign micromatriz[33][99] = 9'b111111111;
assign micromatriz[34][0] = 9'b111111111;
assign micromatriz[34][1] = 9'b111111111;
assign micromatriz[34][2] = 9'b111111111;
assign micromatriz[34][3] = 9'b111111111;
assign micromatriz[34][4] = 9'b111111111;
assign micromatriz[34][5] = 9'b111111111;
assign micromatriz[34][6] = 9'b111111111;
assign micromatriz[34][7] = 9'b111111111;
assign micromatriz[34][8] = 9'b111111111;
assign micromatriz[34][9] = 9'b111111111;
assign micromatriz[34][10] = 9'b111111111;
assign micromatriz[34][11] = 9'b111111111;
assign micromatriz[34][12] = 9'b111111111;
assign micromatriz[34][13] = 9'b111111111;
assign micromatriz[34][14] = 9'b100100100;
assign micromatriz[34][15] = 9'b100000000;
assign micromatriz[34][16] = 9'b101101101;
assign micromatriz[34][17] = 9'b111111111;
assign micromatriz[34][18] = 9'b111111111;
assign micromatriz[34][19] = 9'b111111111;
assign micromatriz[34][20] = 9'b111111111;
assign micromatriz[34][21] = 9'b111111111;
assign micromatriz[34][22] = 9'b111111111;
assign micromatriz[34][23] = 9'b111111111;
assign micromatriz[34][24] = 9'b111111111;
assign micromatriz[34][25] = 9'b111111111;
assign micromatriz[34][26] = 9'b111111111;
assign micromatriz[34][27] = 9'b111111111;
assign micromatriz[34][28] = 9'b111111111;
assign micromatriz[34][29] = 9'b111111111;
assign micromatriz[34][30] = 9'b111111111;
assign micromatriz[34][31] = 9'b111111111;
assign micromatriz[34][32] = 9'b111111111;
assign micromatriz[34][33] = 9'b111111111;
assign micromatriz[34][34] = 9'b111111111;
assign micromatriz[34][35] = 9'b111111111;
assign micromatriz[34][36] = 9'b111111111;
assign micromatriz[34][37] = 9'b111111111;
assign micromatriz[34][38] = 9'b111111111;
assign micromatriz[34][39] = 9'b111111111;
assign micromatriz[34][40] = 9'b111111111;
assign micromatriz[34][41] = 9'b111111111;
assign micromatriz[34][42] = 9'b111111111;
assign micromatriz[34][43] = 9'b111111111;
assign micromatriz[34][44] = 9'b111111111;
assign micromatriz[34][45] = 9'b111111111;
assign micromatriz[34][46] = 9'b111111111;
assign micromatriz[34][47] = 9'b111111111;
assign micromatriz[34][48] = 9'b111111111;
assign micromatriz[34][49] = 9'b111111111;
assign micromatriz[34][50] = 9'b111111111;
assign micromatriz[34][51] = 9'b111111111;
assign micromatriz[34][52] = 9'b111111111;
assign micromatriz[34][53] = 9'b111111111;
assign micromatriz[34][54] = 9'b111111111;
assign micromatriz[34][55] = 9'b111111111;
assign micromatriz[34][56] = 9'b111111111;
assign micromatriz[34][57] = 9'b111111111;
assign micromatriz[34][58] = 9'b111111111;
assign micromatriz[34][59] = 9'b111111111;
assign micromatriz[34][60] = 9'b111111111;
assign micromatriz[34][61] = 9'b111111111;
assign micromatriz[34][62] = 9'b111111111;
assign micromatriz[34][63] = 9'b111111111;
assign micromatriz[34][64] = 9'b110110111;
assign micromatriz[34][65] = 9'b110110111;
assign micromatriz[34][66] = 9'b101101101;
assign micromatriz[34][67] = 9'b100000000;
assign micromatriz[34][68] = 9'b100000000;
assign micromatriz[34][69] = 9'b111111111;
assign micromatriz[34][70] = 9'b111111111;
assign micromatriz[34][71] = 9'b111111111;
assign micromatriz[34][72] = 9'b111111111;
assign micromatriz[34][73] = 9'b110111111;
assign micromatriz[34][74] = 9'b100000000;
assign micromatriz[34][75] = 9'b100000000;
assign micromatriz[34][76] = 9'b100000000;
assign micromatriz[34][77] = 9'b100000000;
assign micromatriz[34][78] = 9'b100100100;
assign micromatriz[34][79] = 9'b111111111;
assign micromatriz[34][80] = 9'b111111111;
assign micromatriz[34][81] = 9'b110110111;
assign micromatriz[34][82] = 9'b110111111;
assign micromatriz[34][83] = 9'b101001001;
assign micromatriz[34][84] = 9'b100000000;
assign micromatriz[34][85] = 9'b100100100;
assign micromatriz[34][86] = 9'b111111111;
assign micromatriz[34][87] = 9'b111111111;
assign micromatriz[34][88] = 9'b111111111;
assign micromatriz[34][89] = 9'b111111111;
assign micromatriz[34][90] = 9'b111111111;
assign micromatriz[34][91] = 9'b111111111;
assign micromatriz[34][92] = 9'b111111111;
assign micromatriz[34][93] = 9'b111111111;
assign micromatriz[34][94] = 9'b111111111;
assign micromatriz[34][95] = 9'b111111111;
assign micromatriz[34][96] = 9'b111111111;
assign micromatriz[34][97] = 9'b111111111;
assign micromatriz[34][98] = 9'b111111111;
assign micromatriz[34][99] = 9'b111111111;
assign micromatriz[35][0] = 9'b111111111;
assign micromatriz[35][1] = 9'b111111111;
assign micromatriz[35][2] = 9'b111111111;
assign micromatriz[35][3] = 9'b111111111;
assign micromatriz[35][4] = 9'b111111111;
assign micromatriz[35][5] = 9'b111111111;
assign micromatriz[35][6] = 9'b111111111;
assign micromatriz[35][7] = 9'b111111111;
assign micromatriz[35][8] = 9'b111111111;
assign micromatriz[35][9] = 9'b111111111;
assign micromatriz[35][10] = 9'b111111111;
assign micromatriz[35][11] = 9'b111111111;
assign micromatriz[35][12] = 9'b111111111;
assign micromatriz[35][13] = 9'b111111111;
assign micromatriz[35][14] = 9'b100100100;
assign micromatriz[35][15] = 9'b100000000;
assign micromatriz[35][16] = 9'b101101101;
assign micromatriz[35][17] = 9'b111111111;
assign micromatriz[35][18] = 9'b111111111;
assign micromatriz[35][19] = 9'b111111111;
assign micromatriz[35][20] = 9'b111111111;
assign micromatriz[35][21] = 9'b110010010;
assign micromatriz[35][22] = 9'b101101101;
assign micromatriz[35][23] = 9'b101110001;
assign micromatriz[35][24] = 9'b101110001;
assign micromatriz[35][25] = 9'b101110001;
assign micromatriz[35][26] = 9'b101110001;
assign micromatriz[35][27] = 9'b101110001;
assign micromatriz[35][28] = 9'b101110001;
assign micromatriz[35][29] = 9'b101110001;
assign micromatriz[35][30] = 9'b101110001;
assign micromatriz[35][31] = 9'b101110001;
assign micromatriz[35][32] = 9'b101110001;
assign micromatriz[35][33] = 9'b101110001;
assign micromatriz[35][34] = 9'b101110001;
assign micromatriz[35][35] = 9'b101110001;
assign micromatriz[35][36] = 9'b101110001;
assign micromatriz[35][37] = 9'b101110001;
assign micromatriz[35][38] = 9'b101110001;
assign micromatriz[35][39] = 9'b101110001;
assign micromatriz[35][40] = 9'b101110001;
assign micromatriz[35][41] = 9'b101110001;
assign micromatriz[35][42] = 9'b101110001;
assign micromatriz[35][43] = 9'b101110001;
assign micromatriz[35][44] = 9'b101110001;
assign micromatriz[35][45] = 9'b101110001;
assign micromatriz[35][46] = 9'b101110001;
assign micromatriz[35][47] = 9'b101110001;
assign micromatriz[35][48] = 9'b101110001;
assign micromatriz[35][49] = 9'b101110001;
assign micromatriz[35][50] = 9'b101110001;
assign micromatriz[35][51] = 9'b101110001;
assign micromatriz[35][52] = 9'b101110001;
assign micromatriz[35][53] = 9'b101110001;
assign micromatriz[35][54] = 9'b101110001;
assign micromatriz[35][55] = 9'b101110001;
assign micromatriz[35][56] = 9'b101110001;
assign micromatriz[35][57] = 9'b101110001;
assign micromatriz[35][58] = 9'b101110001;
assign micromatriz[35][59] = 9'b101110001;
assign micromatriz[35][60] = 9'b101110001;
assign micromatriz[35][61] = 9'b110010001;
assign micromatriz[35][62] = 9'b111111111;
assign micromatriz[35][63] = 9'b111111111;
assign micromatriz[35][64] = 9'b110110111;
assign micromatriz[35][65] = 9'b110110111;
assign micromatriz[35][66] = 9'b101101101;
assign micromatriz[35][67] = 9'b100000000;
assign micromatriz[35][68] = 9'b100000000;
assign micromatriz[35][69] = 9'b111111111;
assign micromatriz[35][70] = 9'b111111111;
assign micromatriz[35][71] = 9'b110110111;
assign micromatriz[35][72] = 9'b101101101;
assign micromatriz[35][73] = 9'b101101101;
assign micromatriz[35][74] = 9'b101001001;
assign micromatriz[35][75] = 9'b101001001;
assign micromatriz[35][76] = 9'b101001001;
assign micromatriz[35][77] = 9'b101001001;
assign micromatriz[35][78] = 9'b101001001;
assign micromatriz[35][79] = 9'b101110001;
assign micromatriz[35][80] = 9'b101110001;
assign micromatriz[35][81] = 9'b110010110;
assign micromatriz[35][82] = 9'b110111111;
assign micromatriz[35][83] = 9'b101001001;
assign micromatriz[35][84] = 9'b100000000;
assign micromatriz[35][85] = 9'b100100100;
assign micromatriz[35][86] = 9'b111111111;
assign micromatriz[35][87] = 9'b111111111;
assign micromatriz[35][88] = 9'b111111111;
assign micromatriz[35][89] = 9'b111111111;
assign micromatriz[35][90] = 9'b111111111;
assign micromatriz[35][91] = 9'b111111111;
assign micromatriz[35][92] = 9'b111111111;
assign micromatriz[35][93] = 9'b111111111;
assign micromatriz[35][94] = 9'b111111111;
assign micromatriz[35][95] = 9'b111111111;
assign micromatriz[35][96] = 9'b111111111;
assign micromatriz[35][97] = 9'b111111111;
assign micromatriz[35][98] = 9'b111111111;
assign micromatriz[35][99] = 9'b111111111;
assign micromatriz[36][0] = 9'b111111111;
assign micromatriz[36][1] = 9'b111111111;
assign micromatriz[36][2] = 9'b111111111;
assign micromatriz[36][3] = 9'b111111111;
assign micromatriz[36][4] = 9'b111111111;
assign micromatriz[36][5] = 9'b111111111;
assign micromatriz[36][6] = 9'b111111111;
assign micromatriz[36][7] = 9'b111111111;
assign micromatriz[36][8] = 9'b111111111;
assign micromatriz[36][9] = 9'b111111111;
assign micromatriz[36][10] = 9'b111111111;
assign micromatriz[36][11] = 9'b111111111;
assign micromatriz[36][12] = 9'b111111111;
assign micromatriz[36][13] = 9'b111111111;
assign micromatriz[36][14] = 9'b100100100;
assign micromatriz[36][15] = 9'b100000000;
assign micromatriz[36][16] = 9'b101101101;
assign micromatriz[36][17] = 9'b111111111;
assign micromatriz[36][18] = 9'b111111111;
assign micromatriz[36][19] = 9'b111111111;
assign micromatriz[36][20] = 9'b111111111;
assign micromatriz[36][21] = 9'b100100100;
assign micromatriz[36][22] = 9'b100000000;
assign micromatriz[36][23] = 9'b100000000;
assign micromatriz[36][24] = 9'b100000000;
assign micromatriz[36][25] = 9'b100000000;
assign micromatriz[36][26] = 9'b100000000;
assign micromatriz[36][27] = 9'b100000000;
assign micromatriz[36][28] = 9'b100000000;
assign micromatriz[36][29] = 9'b100000000;
assign micromatriz[36][30] = 9'b100000000;
assign micromatriz[36][31] = 9'b100000000;
assign micromatriz[36][32] = 9'b100000000;
assign micromatriz[36][33] = 9'b100000000;
assign micromatriz[36][34] = 9'b100000000;
assign micromatriz[36][35] = 9'b100000000;
assign micromatriz[36][36] = 9'b100000000;
assign micromatriz[36][37] = 9'b100000000;
assign micromatriz[36][38] = 9'b100000000;
assign micromatriz[36][39] = 9'b100000000;
assign micromatriz[36][40] = 9'b100000000;
assign micromatriz[36][41] = 9'b100000000;
assign micromatriz[36][42] = 9'b100000000;
assign micromatriz[36][43] = 9'b100000000;
assign micromatriz[36][44] = 9'b100000000;
assign micromatriz[36][45] = 9'b100000000;
assign micromatriz[36][46] = 9'b100000000;
assign micromatriz[36][47] = 9'b100000000;
assign micromatriz[36][48] = 9'b100000000;
assign micromatriz[36][49] = 9'b100000000;
assign micromatriz[36][50] = 9'b100000000;
assign micromatriz[36][51] = 9'b100000000;
assign micromatriz[36][52] = 9'b100000000;
assign micromatriz[36][53] = 9'b100000000;
assign micromatriz[36][54] = 9'b100000000;
assign micromatriz[36][55] = 9'b100000000;
assign micromatriz[36][56] = 9'b100000000;
assign micromatriz[36][57] = 9'b100000000;
assign micromatriz[36][58] = 9'b100000000;
assign micromatriz[36][59] = 9'b100000000;
assign micromatriz[36][60] = 9'b100000000;
assign micromatriz[36][61] = 9'b100000000;
assign micromatriz[36][62] = 9'b110111111;
assign micromatriz[36][63] = 9'b111111111;
assign micromatriz[36][64] = 9'b110110111;
assign micromatriz[36][65] = 9'b110110111;
assign micromatriz[36][66] = 9'b101101101;
assign micromatriz[36][67] = 9'b100000000;
assign micromatriz[36][68] = 9'b100000000;
assign micromatriz[36][69] = 9'b111111111;
assign micromatriz[36][70] = 9'b111111111;
assign micromatriz[36][71] = 9'b101101101;
assign micromatriz[36][72] = 9'b100000000;
assign micromatriz[36][73] = 9'b100000000;
assign micromatriz[36][74] = 9'b111111111;
assign micromatriz[36][75] = 9'b111111111;
assign micromatriz[36][76] = 9'b111111111;
assign micromatriz[36][77] = 9'b111111111;
assign micromatriz[36][78] = 9'b110010010;
assign micromatriz[36][79] = 9'b100000000;
assign micromatriz[36][80] = 9'b100000000;
assign micromatriz[36][81] = 9'b110010010;
assign micromatriz[36][82] = 9'b111111111;
assign micromatriz[36][83] = 9'b101001001;
assign micromatriz[36][84] = 9'b100000000;
assign micromatriz[36][85] = 9'b100100100;
assign micromatriz[36][86] = 9'b111111111;
assign micromatriz[36][87] = 9'b111111111;
assign micromatriz[36][88] = 9'b111111111;
assign micromatriz[36][89] = 9'b111111111;
assign micromatriz[36][90] = 9'b111111111;
assign micromatriz[36][91] = 9'b111111111;
assign micromatriz[36][92] = 9'b111111111;
assign micromatriz[36][93] = 9'b111111111;
assign micromatriz[36][94] = 9'b111111111;
assign micromatriz[36][95] = 9'b111111111;
assign micromatriz[36][96] = 9'b111111111;
assign micromatriz[36][97] = 9'b111111111;
assign micromatriz[36][98] = 9'b111111111;
assign micromatriz[36][99] = 9'b111111111;
assign micromatriz[37][0] = 9'b111111111;
assign micromatriz[37][1] = 9'b111111111;
assign micromatriz[37][2] = 9'b111111111;
assign micromatriz[37][3] = 9'b111111111;
assign micromatriz[37][4] = 9'b111111111;
assign micromatriz[37][5] = 9'b111111111;
assign micromatriz[37][6] = 9'b111111111;
assign micromatriz[37][7] = 9'b111111111;
assign micromatriz[37][8] = 9'b111111111;
assign micromatriz[37][9] = 9'b111111111;
assign micromatriz[37][10] = 9'b111111111;
assign micromatriz[37][11] = 9'b111111111;
assign micromatriz[37][12] = 9'b111111111;
assign micromatriz[37][13] = 9'b111111111;
assign micromatriz[37][14] = 9'b100100100;
assign micromatriz[37][15] = 9'b100000000;
assign micromatriz[37][16] = 9'b101101101;
assign micromatriz[37][17] = 9'b111111111;
assign micromatriz[37][18] = 9'b111111111;
assign micromatriz[37][19] = 9'b111111111;
assign micromatriz[37][20] = 9'b111111111;
assign micromatriz[37][21] = 9'b100101000;
assign micromatriz[37][22] = 9'b100000000;
assign micromatriz[37][23] = 9'b100000000;
assign micromatriz[37][24] = 9'b100000000;
assign micromatriz[37][25] = 9'b100000000;
assign micromatriz[37][26] = 9'b100000000;
assign micromatriz[37][27] = 9'b100000000;
assign micromatriz[37][28] = 9'b100000000;
assign micromatriz[37][29] = 9'b100000000;
assign micromatriz[37][30] = 9'b100000000;
assign micromatriz[37][31] = 9'b100000000;
assign micromatriz[37][32] = 9'b100000000;
assign micromatriz[37][33] = 9'b100000000;
assign micromatriz[37][34] = 9'b100000000;
assign micromatriz[37][35] = 9'b100000000;
assign micromatriz[37][36] = 9'b100000000;
assign micromatriz[37][37] = 9'b100000000;
assign micromatriz[37][38] = 9'b100000000;
assign micromatriz[37][39] = 9'b100000000;
assign micromatriz[37][40] = 9'b100000000;
assign micromatriz[37][41] = 9'b100000000;
assign micromatriz[37][42] = 9'b100000000;
assign micromatriz[37][43] = 9'b100000000;
assign micromatriz[37][44] = 9'b100000000;
assign micromatriz[37][45] = 9'b100000000;
assign micromatriz[37][46] = 9'b100000000;
assign micromatriz[37][47] = 9'b100000000;
assign micromatriz[37][48] = 9'b100000000;
assign micromatriz[37][49] = 9'b100000000;
assign micromatriz[37][50] = 9'b100000000;
assign micromatriz[37][51] = 9'b100000000;
assign micromatriz[37][52] = 9'b100000000;
assign micromatriz[37][53] = 9'b100000000;
assign micromatriz[37][54] = 9'b100000000;
assign micromatriz[37][55] = 9'b100000000;
assign micromatriz[37][56] = 9'b100000000;
assign micromatriz[37][57] = 9'b100000000;
assign micromatriz[37][58] = 9'b100000000;
assign micromatriz[37][59] = 9'b100000000;
assign micromatriz[37][60] = 9'b100000000;
assign micromatriz[37][61] = 9'b100000000;
assign micromatriz[37][62] = 9'b110111111;
assign micromatriz[37][63] = 9'b111111111;
assign micromatriz[37][64] = 9'b110110111;
assign micromatriz[37][65] = 9'b110110111;
assign micromatriz[37][66] = 9'b101101101;
assign micromatriz[37][67] = 9'b100000000;
assign micromatriz[37][68] = 9'b100000000;
assign micromatriz[37][69] = 9'b111111111;
assign micromatriz[37][70] = 9'b111111111;
assign micromatriz[37][71] = 9'b101101101;
assign micromatriz[37][72] = 9'b100000000;
assign micromatriz[37][73] = 9'b100100100;
assign micromatriz[37][74] = 9'b111111111;
assign micromatriz[37][75] = 9'b111111111;
assign micromatriz[37][76] = 9'b111111111;
assign micromatriz[37][77] = 9'b111111111;
assign micromatriz[37][78] = 9'b110010001;
assign micromatriz[37][79] = 9'b100000000;
assign micromatriz[37][80] = 9'b100000000;
assign micromatriz[37][81] = 9'b110010010;
assign micromatriz[37][82] = 9'b111111111;
assign micromatriz[37][83] = 9'b101001001;
assign micromatriz[37][84] = 9'b100000000;
assign micromatriz[37][85] = 9'b100100100;
assign micromatriz[37][86] = 9'b111111111;
assign micromatriz[37][87] = 9'b111111111;
assign micromatriz[37][88] = 9'b111111111;
assign micromatriz[37][89] = 9'b111111111;
assign micromatriz[37][90] = 9'b111111111;
assign micromatriz[37][91] = 9'b111111111;
assign micromatriz[37][92] = 9'b111111111;
assign micromatriz[37][93] = 9'b111111111;
assign micromatriz[37][94] = 9'b111111111;
assign micromatriz[37][95] = 9'b111111111;
assign micromatriz[37][96] = 9'b111111111;
assign micromatriz[37][97] = 9'b111111111;
assign micromatriz[37][98] = 9'b111111111;
assign micromatriz[37][99] = 9'b111111111;
assign micromatriz[38][0] = 9'b111111111;
assign micromatriz[38][1] = 9'b111111111;
assign micromatriz[38][2] = 9'b111111111;
assign micromatriz[38][3] = 9'b111111111;
assign micromatriz[38][4] = 9'b111111111;
assign micromatriz[38][5] = 9'b111111111;
assign micromatriz[38][6] = 9'b111111111;
assign micromatriz[38][7] = 9'b111111111;
assign micromatriz[38][8] = 9'b111111111;
assign micromatriz[38][9] = 9'b111111111;
assign micromatriz[38][10] = 9'b111111111;
assign micromatriz[38][11] = 9'b111111111;
assign micromatriz[38][12] = 9'b111111111;
assign micromatriz[38][13] = 9'b111111111;
assign micromatriz[38][14] = 9'b100100100;
assign micromatriz[38][15] = 9'b100000000;
assign micromatriz[38][16] = 9'b101101101;
assign micromatriz[38][17] = 9'b111111111;
assign micromatriz[38][18] = 9'b111111111;
assign micromatriz[38][19] = 9'b111111111;
assign micromatriz[38][20] = 9'b111111111;
assign micromatriz[38][21] = 9'b100101000;
assign micromatriz[38][22] = 9'b100000000;
assign micromatriz[38][23] = 9'b100100100;
assign micromatriz[38][24] = 9'b101101101;
assign micromatriz[38][25] = 9'b101001001;
assign micromatriz[38][26] = 9'b101001001;
assign micromatriz[38][27] = 9'b101001001;
assign micromatriz[38][28] = 9'b101001001;
assign micromatriz[38][29] = 9'b101001001;
assign micromatriz[38][30] = 9'b101001001;
assign micromatriz[38][31] = 9'b101001001;
assign micromatriz[38][32] = 9'b101001001;
assign micromatriz[38][33] = 9'b101001001;
assign micromatriz[38][34] = 9'b101001001;
assign micromatriz[38][35] = 9'b101001001;
assign micromatriz[38][36] = 9'b101001001;
assign micromatriz[38][37] = 9'b101001001;
assign micromatriz[38][38] = 9'b101001001;
assign micromatriz[38][39] = 9'b101001001;
assign micromatriz[38][40] = 9'b101001001;
assign micromatriz[38][41] = 9'b101001001;
assign micromatriz[38][42] = 9'b101001001;
assign micromatriz[38][43] = 9'b101001001;
assign micromatriz[38][44] = 9'b101001001;
assign micromatriz[38][45] = 9'b101001001;
assign micromatriz[38][46] = 9'b101001001;
assign micromatriz[38][47] = 9'b101001001;
assign micromatriz[38][48] = 9'b101001001;
assign micromatriz[38][49] = 9'b101001001;
assign micromatriz[38][50] = 9'b101001001;
assign micromatriz[38][51] = 9'b101001001;
assign micromatriz[38][52] = 9'b101001001;
assign micromatriz[38][53] = 9'b101001001;
assign micromatriz[38][54] = 9'b101001001;
assign micromatriz[38][55] = 9'b101001001;
assign micromatriz[38][56] = 9'b101001001;
assign micromatriz[38][57] = 9'b101101101;
assign micromatriz[38][58] = 9'b101101101;
assign micromatriz[38][59] = 9'b100100100;
assign micromatriz[38][60] = 9'b100000000;
assign micromatriz[38][61] = 9'b100000000;
assign micromatriz[38][62] = 9'b110111111;
assign micromatriz[38][63] = 9'b111111111;
assign micromatriz[38][64] = 9'b110110111;
assign micromatriz[38][65] = 9'b110110111;
assign micromatriz[38][66] = 9'b101101101;
assign micromatriz[38][67] = 9'b100000000;
assign micromatriz[38][68] = 9'b100000000;
assign micromatriz[38][69] = 9'b111111111;
assign micromatriz[38][70] = 9'b111111111;
assign micromatriz[38][71] = 9'b101101101;
assign micromatriz[38][72] = 9'b100000000;
assign micromatriz[38][73] = 9'b100000000;
assign micromatriz[38][74] = 9'b111111111;
assign micromatriz[38][75] = 9'b111111111;
assign micromatriz[38][76] = 9'b110110111;
assign micromatriz[38][77] = 9'b110111111;
assign micromatriz[38][78] = 9'b101101101;
assign micromatriz[38][79] = 9'b100000000;
assign micromatriz[38][80] = 9'b100000000;
assign micromatriz[38][81] = 9'b110010010;
assign micromatriz[38][82] = 9'b111111111;
assign micromatriz[38][83] = 9'b101001001;
assign micromatriz[38][84] = 9'b100000000;
assign micromatriz[38][85] = 9'b100100100;
assign micromatriz[38][86] = 9'b111111111;
assign micromatriz[38][87] = 9'b111111111;
assign micromatriz[38][88] = 9'b111111111;
assign micromatriz[38][89] = 9'b111111111;
assign micromatriz[38][90] = 9'b111111111;
assign micromatriz[38][91] = 9'b111111111;
assign micromatriz[38][92] = 9'b111111111;
assign micromatriz[38][93] = 9'b111111111;
assign micromatriz[38][94] = 9'b111111111;
assign micromatriz[38][95] = 9'b111111111;
assign micromatriz[38][96] = 9'b111111111;
assign micromatriz[38][97] = 9'b111111111;
assign micromatriz[38][98] = 9'b111111111;
assign micromatriz[38][99] = 9'b111111111;
assign micromatriz[39][0] = 9'b111111111;
assign micromatriz[39][1] = 9'b111111111;
assign micromatriz[39][2] = 9'b111111111;
assign micromatriz[39][3] = 9'b111111111;
assign micromatriz[39][4] = 9'b111111111;
assign micromatriz[39][5] = 9'b111111111;
assign micromatriz[39][6] = 9'b111111111;
assign micromatriz[39][7] = 9'b111111111;
assign micromatriz[39][8] = 9'b111111111;
assign micromatriz[39][9] = 9'b111111111;
assign micromatriz[39][10] = 9'b111111111;
assign micromatriz[39][11] = 9'b111111111;
assign micromatriz[39][12] = 9'b111111111;
assign micromatriz[39][13] = 9'b111111111;
assign micromatriz[39][14] = 9'b100100100;
assign micromatriz[39][15] = 9'b100000000;
assign micromatriz[39][16] = 9'b101101101;
assign micromatriz[39][17] = 9'b111111111;
assign micromatriz[39][18] = 9'b111111111;
assign micromatriz[39][19] = 9'b111111111;
assign micromatriz[39][20] = 9'b111111111;
assign micromatriz[39][21] = 9'b100101000;
assign micromatriz[39][22] = 9'b100000000;
assign micromatriz[39][23] = 9'b100100100;
assign micromatriz[39][24] = 9'b101101101;
assign micromatriz[39][25] = 9'b101101101;
assign micromatriz[39][26] = 9'b101101101;
assign micromatriz[39][27] = 9'b101101101;
assign micromatriz[39][28] = 9'b101101101;
assign micromatriz[39][29] = 9'b101101101;
assign micromatriz[39][30] = 9'b101101101;
assign micromatriz[39][31] = 9'b101101101;
assign micromatriz[39][32] = 9'b101101101;
assign micromatriz[39][33] = 9'b101101101;
assign micromatriz[39][34] = 9'b101101101;
assign micromatriz[39][35] = 9'b101101101;
assign micromatriz[39][36] = 9'b101101101;
assign micromatriz[39][37] = 9'b101101101;
assign micromatriz[39][38] = 9'b101101101;
assign micromatriz[39][39] = 9'b101101101;
assign micromatriz[39][40] = 9'b101101101;
assign micromatriz[39][41] = 9'b101101101;
assign micromatriz[39][42] = 9'b101101101;
assign micromatriz[39][43] = 9'b101101101;
assign micromatriz[39][44] = 9'b101101101;
assign micromatriz[39][45] = 9'b101101101;
assign micromatriz[39][46] = 9'b101101101;
assign micromatriz[39][47] = 9'b101101101;
assign micromatriz[39][48] = 9'b101101101;
assign micromatriz[39][49] = 9'b101101101;
assign micromatriz[39][50] = 9'b101101101;
assign micromatriz[39][51] = 9'b101101101;
assign micromatriz[39][52] = 9'b101101101;
assign micromatriz[39][53] = 9'b101101101;
assign micromatriz[39][54] = 9'b101101101;
assign micromatriz[39][55] = 9'b101101101;
assign micromatriz[39][56] = 9'b101101101;
assign micromatriz[39][57] = 9'b101101101;
assign micromatriz[39][58] = 9'b101101101;
assign micromatriz[39][59] = 9'b101001000;
assign micromatriz[39][60] = 9'b100000000;
assign micromatriz[39][61] = 9'b100000000;
assign micromatriz[39][62] = 9'b110111111;
assign micromatriz[39][63] = 9'b111111111;
assign micromatriz[39][64] = 9'b110110111;
assign micromatriz[39][65] = 9'b110110111;
assign micromatriz[39][66] = 9'b101101101;
assign micromatriz[39][67] = 9'b100000000;
assign micromatriz[39][68] = 9'b100000000;
assign micromatriz[39][69] = 9'b111111111;
assign micromatriz[39][70] = 9'b111111111;
assign micromatriz[39][71] = 9'b101101101;
assign micromatriz[39][72] = 9'b100000000;
assign micromatriz[39][73] = 9'b100000000;
assign micromatriz[39][74] = 9'b111111111;
assign micromatriz[39][75] = 9'b111111111;
assign micromatriz[39][76] = 9'b111111111;
assign micromatriz[39][77] = 9'b111111111;
assign micromatriz[39][78] = 9'b101101101;
assign micromatriz[39][79] = 9'b100000000;
assign micromatriz[39][80] = 9'b100000000;
assign micromatriz[39][81] = 9'b110010010;
assign micromatriz[39][82] = 9'b111111111;
assign micromatriz[39][83] = 9'b101001001;
assign micromatriz[39][84] = 9'b100000000;
assign micromatriz[39][85] = 9'b100100100;
assign micromatriz[39][86] = 9'b111111111;
assign micromatriz[39][87] = 9'b111111111;
assign micromatriz[39][88] = 9'b111111111;
assign micromatriz[39][89] = 9'b111111111;
assign micromatriz[39][90] = 9'b111111111;
assign micromatriz[39][91] = 9'b111111111;
assign micromatriz[39][92] = 9'b111111111;
assign micromatriz[39][93] = 9'b111111111;
assign micromatriz[39][94] = 9'b111111111;
assign micromatriz[39][95] = 9'b111111111;
assign micromatriz[39][96] = 9'b111111111;
assign micromatriz[39][97] = 9'b111111111;
assign micromatriz[39][98] = 9'b111111111;
assign micromatriz[39][99] = 9'b111111111;
assign micromatriz[40][0] = 9'b111111111;
assign micromatriz[40][1] = 9'b111111111;
assign micromatriz[40][2] = 9'b111111111;
assign micromatriz[40][3] = 9'b111111111;
assign micromatriz[40][4] = 9'b111111111;
assign micromatriz[40][5] = 9'b111111111;
assign micromatriz[40][6] = 9'b111111111;
assign micromatriz[40][7] = 9'b111111111;
assign micromatriz[40][8] = 9'b111111111;
assign micromatriz[40][9] = 9'b111111111;
assign micromatriz[40][10] = 9'b111111111;
assign micromatriz[40][11] = 9'b111111111;
assign micromatriz[40][12] = 9'b111111111;
assign micromatriz[40][13] = 9'b111111111;
assign micromatriz[40][14] = 9'b100100100;
assign micromatriz[40][15] = 9'b100000000;
assign micromatriz[40][16] = 9'b101101101;
assign micromatriz[40][17] = 9'b111111111;
assign micromatriz[40][18] = 9'b111111111;
assign micromatriz[40][19] = 9'b111111111;
assign micromatriz[40][20] = 9'b111111111;
assign micromatriz[40][21] = 9'b100101000;
assign micromatriz[40][22] = 9'b100000000;
assign micromatriz[40][23] = 9'b100100100;
assign micromatriz[40][24] = 9'b101101101;
assign micromatriz[40][25] = 9'b101101101;
assign micromatriz[40][26] = 9'b101101101;
assign micromatriz[40][27] = 9'b101101101;
assign micromatriz[40][28] = 9'b101101101;
assign micromatriz[40][29] = 9'b101101101;
assign micromatriz[40][30] = 9'b101101101;
assign micromatriz[40][31] = 9'b101101101;
assign micromatriz[40][32] = 9'b101101101;
assign micromatriz[40][33] = 9'b101101101;
assign micromatriz[40][34] = 9'b101101101;
assign micromatriz[40][35] = 9'b101101101;
assign micromatriz[40][36] = 9'b101101101;
assign micromatriz[40][37] = 9'b101101101;
assign micromatriz[40][38] = 9'b101101101;
assign micromatriz[40][39] = 9'b101101101;
assign micromatriz[40][40] = 9'b101101101;
assign micromatriz[40][41] = 9'b101101101;
assign micromatriz[40][42] = 9'b101101101;
assign micromatriz[40][43] = 9'b101101101;
assign micromatriz[40][44] = 9'b101101101;
assign micromatriz[40][45] = 9'b101101101;
assign micromatriz[40][46] = 9'b101101101;
assign micromatriz[40][47] = 9'b101101101;
assign micromatriz[40][48] = 9'b101101101;
assign micromatriz[40][49] = 9'b101101101;
assign micromatriz[40][50] = 9'b101101101;
assign micromatriz[40][51] = 9'b101101101;
assign micromatriz[40][52] = 9'b101101101;
assign micromatriz[40][53] = 9'b101101101;
assign micromatriz[40][54] = 9'b101101101;
assign micromatriz[40][55] = 9'b101101101;
assign micromatriz[40][56] = 9'b101101101;
assign micromatriz[40][57] = 9'b110010001;
assign micromatriz[40][58] = 9'b110010001;
assign micromatriz[40][59] = 9'b101001001;
assign micromatriz[40][60] = 9'b100000000;
assign micromatriz[40][61] = 9'b100000000;
assign micromatriz[40][62] = 9'b110111111;
assign micromatriz[40][63] = 9'b111111111;
assign micromatriz[40][64] = 9'b110110111;
assign micromatriz[40][65] = 9'b110110111;
assign micromatriz[40][66] = 9'b101101101;
assign micromatriz[40][67] = 9'b100000000;
assign micromatriz[40][68] = 9'b100000000;
assign micromatriz[40][69] = 9'b111111111;
assign micromatriz[40][70] = 9'b111111111;
assign micromatriz[40][71] = 9'b110110110;
assign micromatriz[40][72] = 9'b101101101;
assign micromatriz[40][73] = 9'b101101101;
assign micromatriz[40][74] = 9'b101001001;
assign micromatriz[40][75] = 9'b101001001;
assign micromatriz[40][76] = 9'b101001001;
assign micromatriz[40][77] = 9'b101001001;
assign micromatriz[40][78] = 9'b101001001;
assign micromatriz[40][79] = 9'b101101101;
assign micromatriz[40][80] = 9'b101101101;
assign micromatriz[40][81] = 9'b110010010;
assign micromatriz[40][82] = 9'b110111111;
assign micromatriz[40][83] = 9'b101001001;
assign micromatriz[40][84] = 9'b100000000;
assign micromatriz[40][85] = 9'b100100100;
assign micromatriz[40][86] = 9'b111111111;
assign micromatriz[40][87] = 9'b111111111;
assign micromatriz[40][88] = 9'b111111111;
assign micromatriz[40][89] = 9'b111111111;
assign micromatriz[40][90] = 9'b111111111;
assign micromatriz[40][91] = 9'b111111111;
assign micromatriz[40][92] = 9'b111111111;
assign micromatriz[40][93] = 9'b111111111;
assign micromatriz[40][94] = 9'b111111111;
assign micromatriz[40][95] = 9'b111111111;
assign micromatriz[40][96] = 9'b111111111;
assign micromatriz[40][97] = 9'b111111111;
assign micromatriz[40][98] = 9'b111111111;
assign micromatriz[40][99] = 9'b111111111;
assign micromatriz[41][0] = 9'b111111111;
assign micromatriz[41][1] = 9'b111111111;
assign micromatriz[41][2] = 9'b111111111;
assign micromatriz[41][3] = 9'b111111111;
assign micromatriz[41][4] = 9'b111111111;
assign micromatriz[41][5] = 9'b111111111;
assign micromatriz[41][6] = 9'b111111111;
assign micromatriz[41][7] = 9'b111111111;
assign micromatriz[41][8] = 9'b111111111;
assign micromatriz[41][9] = 9'b111111111;
assign micromatriz[41][10] = 9'b111111111;
assign micromatriz[41][11] = 9'b111111111;
assign micromatriz[41][12] = 9'b111111111;
assign micromatriz[41][13] = 9'b111111111;
assign micromatriz[41][14] = 9'b100100100;
assign micromatriz[41][15] = 9'b100000000;
assign micromatriz[41][16] = 9'b101101101;
assign micromatriz[41][17] = 9'b111111111;
assign micromatriz[41][18] = 9'b111111111;
assign micromatriz[41][19] = 9'b111111111;
assign micromatriz[41][20] = 9'b111111111;
assign micromatriz[41][21] = 9'b100101000;
assign micromatriz[41][22] = 9'b100000000;
assign micromatriz[41][23] = 9'b100100100;
assign micromatriz[41][24] = 9'b101101101;
assign micromatriz[41][25] = 9'b101001101;
assign micromatriz[41][26] = 9'b110010001;
assign micromatriz[41][27] = 9'b111111100;
assign micromatriz[41][28] = 9'b111111100;
assign micromatriz[41][29] = 9'b111111100;
assign micromatriz[41][30] = 9'b111111100;
assign micromatriz[41][31] = 9'b111111100;
assign micromatriz[41][32] = 9'b111111100;
assign micromatriz[41][33] = 9'b111111100;
assign micromatriz[41][34] = 9'b111111100;
assign micromatriz[41][35] = 9'b111111100;
assign micromatriz[41][36] = 9'b111111100;
assign micromatriz[41][37] = 9'b111111100;
assign micromatriz[41][38] = 9'b111111100;
assign micromatriz[41][39] = 9'b111111100;
assign micromatriz[41][40] = 9'b111111100;
assign micromatriz[41][41] = 9'b111111100;
assign micromatriz[41][42] = 9'b111111100;
assign micromatriz[41][43] = 9'b111111100;
assign micromatriz[41][44] = 9'b111111100;
assign micromatriz[41][45] = 9'b111111100;
assign micromatriz[41][46] = 9'b111111100;
assign micromatriz[41][47] = 9'b111111100;
assign micromatriz[41][48] = 9'b111111100;
assign micromatriz[41][49] = 9'b111111100;
assign micromatriz[41][50] = 9'b111111100;
assign micromatriz[41][51] = 9'b111111100;
assign micromatriz[41][52] = 9'b111111100;
assign micromatriz[41][53] = 9'b111111100;
assign micromatriz[41][54] = 9'b111111100;
assign micromatriz[41][55] = 9'b111111100;
assign micromatriz[41][56] = 9'b110010001;
assign micromatriz[41][57] = 9'b110010010;
assign micromatriz[41][58] = 9'b110110110;
assign micromatriz[41][59] = 9'b101001001;
assign micromatriz[41][60] = 9'b100000000;
assign micromatriz[41][61] = 9'b100000000;
assign micromatriz[41][62] = 9'b110111111;
assign micromatriz[41][63] = 9'b111111111;
assign micromatriz[41][64] = 9'b110110111;
assign micromatriz[41][65] = 9'b110110111;
assign micromatriz[41][66] = 9'b101101101;
assign micromatriz[41][67] = 9'b100000000;
assign micromatriz[41][68] = 9'b100000000;
assign micromatriz[41][69] = 9'b111111111;
assign micromatriz[41][70] = 9'b111111111;
assign micromatriz[41][71] = 9'b111111111;
assign micromatriz[41][72] = 9'b111111111;
assign micromatriz[41][73] = 9'b110111111;
assign micromatriz[41][74] = 9'b100000000;
assign micromatriz[41][75] = 9'b100000000;
assign micromatriz[41][76] = 9'b100000000;
assign micromatriz[41][77] = 9'b100000000;
assign micromatriz[41][78] = 9'b100100100;
assign micromatriz[41][79] = 9'b111111111;
assign micromatriz[41][80] = 9'b111111111;
assign micromatriz[41][81] = 9'b110110111;
assign micromatriz[41][82] = 9'b110111111;
assign micromatriz[41][83] = 9'b101001001;
assign micromatriz[41][84] = 9'b100000000;
assign micromatriz[41][85] = 9'b100100100;
assign micromatriz[41][86] = 9'b111111111;
assign micromatriz[41][87] = 9'b111111111;
assign micromatriz[41][88] = 9'b111111111;
assign micromatriz[41][89] = 9'b111111111;
assign micromatriz[41][90] = 9'b111111111;
assign micromatriz[41][91] = 9'b111111111;
assign micromatriz[41][92] = 9'b111111111;
assign micromatriz[41][93] = 9'b111111111;
assign micromatriz[41][94] = 9'b111111111;
assign micromatriz[41][95] = 9'b111111111;
assign micromatriz[41][96] = 9'b111111111;
assign micromatriz[41][97] = 9'b111111111;
assign micromatriz[41][98] = 9'b111111111;
assign micromatriz[41][99] = 9'b111111111;
assign micromatriz[42][0] = 9'b111111111;
assign micromatriz[42][1] = 9'b111111111;
assign micromatriz[42][2] = 9'b111111111;
assign micromatriz[42][3] = 9'b111111111;
assign micromatriz[42][4] = 9'b111111111;
assign micromatriz[42][5] = 9'b111111111;
assign micromatriz[42][6] = 9'b111111111;
assign micromatriz[42][7] = 9'b111111111;
assign micromatriz[42][8] = 9'b111111111;
assign micromatriz[42][9] = 9'b111111111;
assign micromatriz[42][10] = 9'b111111111;
assign micromatriz[42][11] = 9'b111111111;
assign micromatriz[42][12] = 9'b111111111;
assign micromatriz[42][13] = 9'b111111111;
assign micromatriz[42][14] = 9'b100100100;
assign micromatriz[42][15] = 9'b100000000;
assign micromatriz[42][16] = 9'b101101101;
assign micromatriz[42][17] = 9'b111111111;
assign micromatriz[42][18] = 9'b111111111;
assign micromatriz[42][19] = 9'b111111111;
assign micromatriz[42][20] = 9'b111111111;
assign micromatriz[42][21] = 9'b100101000;
assign micromatriz[42][22] = 9'b100000000;
assign micromatriz[42][23] = 9'b100100100;
assign micromatriz[42][24] = 9'b101101101;
assign micromatriz[42][25] = 9'b101001101;
assign micromatriz[42][26] = 9'b110001101;
assign micromatriz[42][27] = 9'b111111100;
assign micromatriz[42][28] = 9'b111111100;
assign micromatriz[42][29] = 9'b111111100;
assign micromatriz[42][30] = 9'b111111100;
assign micromatriz[42][31] = 9'b111111100;
assign micromatriz[42][32] = 9'b111111100;
assign micromatriz[42][33] = 9'b111111100;
assign micromatriz[42][34] = 9'b111111100;
assign micromatriz[42][35] = 9'b111111100;
assign micromatriz[42][36] = 9'b111111100;
assign micromatriz[42][37] = 9'b111111100;
assign micromatriz[42][38] = 9'b111111100;
assign micromatriz[42][39] = 9'b111111100;
assign micromatriz[42][40] = 9'b111111100;
assign micromatriz[42][41] = 9'b111111100;
assign micromatriz[42][42] = 9'b111111100;
assign micromatriz[42][43] = 9'b111111100;
assign micromatriz[42][44] = 9'b111111100;
assign micromatriz[42][45] = 9'b111111100;
assign micromatriz[42][46] = 9'b111111100;
assign micromatriz[42][47] = 9'b111111100;
assign micromatriz[42][48] = 9'b111111100;
assign micromatriz[42][49] = 9'b111111100;
assign micromatriz[42][50] = 9'b111111100;
assign micromatriz[42][51] = 9'b111111100;
assign micromatriz[42][52] = 9'b111111100;
assign micromatriz[42][53] = 9'b111111100;
assign micromatriz[42][54] = 9'b111111100;
assign micromatriz[42][55] = 9'b111111100;
assign micromatriz[42][56] = 9'b110010001;
assign micromatriz[42][57] = 9'b110010010;
assign micromatriz[42][58] = 9'b110110110;
assign micromatriz[42][59] = 9'b101001001;
assign micromatriz[42][60] = 9'b100000000;
assign micromatriz[42][61] = 9'b100000000;
assign micromatriz[42][62] = 9'b110111111;
assign micromatriz[42][63] = 9'b111111111;
assign micromatriz[42][64] = 9'b110110111;
assign micromatriz[42][65] = 9'b110110111;
assign micromatriz[42][66] = 9'b101101101;
assign micromatriz[42][67] = 9'b100000000;
assign micromatriz[42][68] = 9'b100000000;
assign micromatriz[42][69] = 9'b111111111;
assign micromatriz[42][70] = 9'b111111111;
assign micromatriz[42][71] = 9'b111111111;
assign micromatriz[42][72] = 9'b111111111;
assign micromatriz[42][73] = 9'b110110111;
assign micromatriz[42][74] = 9'b100100100;
assign micromatriz[42][75] = 9'b100100100;
assign micromatriz[42][76] = 9'b100100100;
assign micromatriz[42][77] = 9'b100100100;
assign micromatriz[42][78] = 9'b101001001;
assign micromatriz[42][79] = 9'b111111111;
assign micromatriz[42][80] = 9'b111111111;
assign micromatriz[42][81] = 9'b110110111;
assign micromatriz[42][82] = 9'b110111111;
assign micromatriz[42][83] = 9'b101001001;
assign micromatriz[42][84] = 9'b100000000;
assign micromatriz[42][85] = 9'b100100100;
assign micromatriz[42][86] = 9'b111111111;
assign micromatriz[42][87] = 9'b111111111;
assign micromatriz[42][88] = 9'b111111111;
assign micromatriz[42][89] = 9'b111111111;
assign micromatriz[42][90] = 9'b111111111;
assign micromatriz[42][91] = 9'b111111111;
assign micromatriz[42][92] = 9'b111111111;
assign micromatriz[42][93] = 9'b111111111;
assign micromatriz[42][94] = 9'b111111111;
assign micromatriz[42][95] = 9'b111111111;
assign micromatriz[42][96] = 9'b111111111;
assign micromatriz[42][97] = 9'b111111111;
assign micromatriz[42][98] = 9'b111111111;
assign micromatriz[42][99] = 9'b111111111;
assign micromatriz[43][0] = 9'b111111111;
assign micromatriz[43][1] = 9'b111111111;
assign micromatriz[43][2] = 9'b111111111;
assign micromatriz[43][3] = 9'b111111111;
assign micromatriz[43][4] = 9'b111111111;
assign micromatriz[43][5] = 9'b111111111;
assign micromatriz[43][6] = 9'b111111111;
assign micromatriz[43][7] = 9'b111111111;
assign micromatriz[43][8] = 9'b111111111;
assign micromatriz[43][9] = 9'b111111111;
assign micromatriz[43][10] = 9'b111111111;
assign micromatriz[43][11] = 9'b111111111;
assign micromatriz[43][12] = 9'b111111111;
assign micromatriz[43][13] = 9'b111111111;
assign micromatriz[43][14] = 9'b100100100;
assign micromatriz[43][15] = 9'b100000000;
assign micromatriz[43][16] = 9'b101101101;
assign micromatriz[43][17] = 9'b111111111;
assign micromatriz[43][18] = 9'b111111111;
assign micromatriz[43][19] = 9'b111111111;
assign micromatriz[43][20] = 9'b111111111;
assign micromatriz[43][21] = 9'b100101000;
assign micromatriz[43][22] = 9'b100000000;
assign micromatriz[43][23] = 9'b100100100;
assign micromatriz[43][24] = 9'b101101101;
assign micromatriz[43][25] = 9'b101001101;
assign micromatriz[43][26] = 9'b110001101;
assign micromatriz[43][27] = 9'b111111100;
assign micromatriz[43][28] = 9'b111111100;
assign micromatriz[43][29] = 9'b111111100;
assign micromatriz[43][30] = 9'b111111100;
assign micromatriz[43][31] = 9'b111111100;
assign micromatriz[43][32] = 9'b111111100;
assign micromatriz[43][33] = 9'b111111100;
assign micromatriz[43][34] = 9'b111111100;
assign micromatriz[43][35] = 9'b111111100;
assign micromatriz[43][36] = 9'b111111100;
assign micromatriz[43][37] = 9'b111111100;
assign micromatriz[43][38] = 9'b111111100;
assign micromatriz[43][39] = 9'b111111100;
assign micromatriz[43][40] = 9'b111111100;
assign micromatriz[43][41] = 9'b111111100;
assign micromatriz[43][42] = 9'b111111100;
assign micromatriz[43][43] = 9'b111111100;
assign micromatriz[43][44] = 9'b111111100;
assign micromatriz[43][45] = 9'b111111100;
assign micromatriz[43][46] = 9'b111111100;
assign micromatriz[43][47] = 9'b111111100;
assign micromatriz[43][48] = 9'b111111100;
assign micromatriz[43][49] = 9'b111111100;
assign micromatriz[43][50] = 9'b111111100;
assign micromatriz[43][51] = 9'b111111100;
assign micromatriz[43][52] = 9'b111111100;
assign micromatriz[43][53] = 9'b111111100;
assign micromatriz[43][54] = 9'b111111100;
assign micromatriz[43][55] = 9'b111111100;
assign micromatriz[43][56] = 9'b110010001;
assign micromatriz[43][57] = 9'b110010010;
assign micromatriz[43][58] = 9'b110110110;
assign micromatriz[43][59] = 9'b101001001;
assign micromatriz[43][60] = 9'b100000000;
assign micromatriz[43][61] = 9'b100000000;
assign micromatriz[43][62] = 9'b110111111;
assign micromatriz[43][63] = 9'b111111111;
assign micromatriz[43][64] = 9'b110110111;
assign micromatriz[43][65] = 9'b110110111;
assign micromatriz[43][66] = 9'b101101101;
assign micromatriz[43][67] = 9'b100000000;
assign micromatriz[43][68] = 9'b100000000;
assign micromatriz[43][69] = 9'b111111111;
assign micromatriz[43][70] = 9'b111111111;
assign micromatriz[43][71] = 9'b111111111;
assign micromatriz[43][72] = 9'b111111111;
assign micromatriz[43][73] = 9'b111111111;
assign micromatriz[43][74] = 9'b111111111;
assign micromatriz[43][75] = 9'b111111111;
assign micromatriz[43][76] = 9'b111111111;
assign micromatriz[43][77] = 9'b111111111;
assign micromatriz[43][78] = 9'b111111111;
assign micromatriz[43][79] = 9'b111111111;
assign micromatriz[43][80] = 9'b111111111;
assign micromatriz[43][81] = 9'b110110111;
assign micromatriz[43][82] = 9'b110111111;
assign micromatriz[43][83] = 9'b101001001;
assign micromatriz[43][84] = 9'b100000000;
assign micromatriz[43][85] = 9'b100100100;
assign micromatriz[43][86] = 9'b111111111;
assign micromatriz[43][87] = 9'b111111111;
assign micromatriz[43][88] = 9'b111111111;
assign micromatriz[43][89] = 9'b111111111;
assign micromatriz[43][90] = 9'b111111111;
assign micromatriz[43][91] = 9'b111111111;
assign micromatriz[43][92] = 9'b111111111;
assign micromatriz[43][93] = 9'b111111111;
assign micromatriz[43][94] = 9'b111111111;
assign micromatriz[43][95] = 9'b111111111;
assign micromatriz[43][96] = 9'b111111111;
assign micromatriz[43][97] = 9'b111111111;
assign micromatriz[43][98] = 9'b111111111;
assign micromatriz[43][99] = 9'b111111111;
assign micromatriz[44][0] = 9'b111111111;
assign micromatriz[44][1] = 9'b111111111;
assign micromatriz[44][2] = 9'b111111111;
assign micromatriz[44][3] = 9'b111111111;
assign micromatriz[44][4] = 9'b111111111;
assign micromatriz[44][5] = 9'b111111111;
assign micromatriz[44][6] = 9'b111111111;
assign micromatriz[44][7] = 9'b111111111;
assign micromatriz[44][8] = 9'b111111111;
assign micromatriz[44][9] = 9'b111111111;
assign micromatriz[44][10] = 9'b111111111;
assign micromatriz[44][11] = 9'b111111111;
assign micromatriz[44][12] = 9'b111111111;
assign micromatriz[44][13] = 9'b111111111;
assign micromatriz[44][14] = 9'b100100100;
assign micromatriz[44][15] = 9'b100000000;
assign micromatriz[44][16] = 9'b101101101;
assign micromatriz[44][17] = 9'b111111111;
assign micromatriz[44][18] = 9'b111111111;
assign micromatriz[44][19] = 9'b111111111;
assign micromatriz[44][20] = 9'b111111111;
assign micromatriz[44][21] = 9'b100101000;
assign micromatriz[44][22] = 9'b100000000;
assign micromatriz[44][23] = 9'b100100100;
assign micromatriz[44][24] = 9'b101101101;
assign micromatriz[44][25] = 9'b101001101;
assign micromatriz[44][26] = 9'b110001101;
assign micromatriz[44][27] = 9'b111111100;
assign micromatriz[44][28] = 9'b111111100;
assign micromatriz[44][29] = 9'b111111100;
assign micromatriz[44][30] = 9'b111111100;
assign micromatriz[44][31] = 9'b111111100;
assign micromatriz[44][32] = 9'b111111100;
assign micromatriz[44][33] = 9'b111111100;
assign micromatriz[44][34] = 9'b111111100;
assign micromatriz[44][35] = 9'b111111100;
assign micromatriz[44][36] = 9'b111111100;
assign micromatriz[44][37] = 9'b111111100;
assign micromatriz[44][38] = 9'b111111100;
assign micromatriz[44][39] = 9'b111111100;
assign micromatriz[44][40] = 9'b111111100;
assign micromatriz[44][41] = 9'b111111100;
assign micromatriz[44][42] = 9'b111111100;
assign micromatriz[44][43] = 9'b111111100;
assign micromatriz[44][44] = 9'b111111100;
assign micromatriz[44][45] = 9'b111111100;
assign micromatriz[44][46] = 9'b111111100;
assign micromatriz[44][47] = 9'b111111100;
assign micromatriz[44][48] = 9'b111111100;
assign micromatriz[44][49] = 9'b111111100;
assign micromatriz[44][50] = 9'b111111100;
assign micromatriz[44][51] = 9'b111111100;
assign micromatriz[44][52] = 9'b111111100;
assign micromatriz[44][53] = 9'b111111100;
assign micromatriz[44][54] = 9'b111111100;
assign micromatriz[44][55] = 9'b111111100;
assign micromatriz[44][56] = 9'b110010001;
assign micromatriz[44][57] = 9'b110010010;
assign micromatriz[44][58] = 9'b110110110;
assign micromatriz[44][59] = 9'b101001001;
assign micromatriz[44][60] = 9'b100000000;
assign micromatriz[44][61] = 9'b100000000;
assign micromatriz[44][62] = 9'b110111111;
assign micromatriz[44][63] = 9'b111111111;
assign micromatriz[44][64] = 9'b110110111;
assign micromatriz[44][65] = 9'b110110111;
assign micromatriz[44][66] = 9'b101101101;
assign micromatriz[44][67] = 9'b100000000;
assign micromatriz[44][68] = 9'b100000000;
assign micromatriz[44][69] = 9'b111111111;
assign micromatriz[44][70] = 9'b111111111;
assign micromatriz[44][71] = 9'b111111111;
assign micromatriz[44][72] = 9'b111111111;
assign micromatriz[44][73] = 9'b111111111;
assign micromatriz[44][74] = 9'b111111111;
assign micromatriz[44][75] = 9'b111111111;
assign micromatriz[44][76] = 9'b111111111;
assign micromatriz[44][77] = 9'b111111111;
assign micromatriz[44][78] = 9'b111111111;
assign micromatriz[44][79] = 9'b111111111;
assign micromatriz[44][80] = 9'b111111111;
assign micromatriz[44][81] = 9'b110110111;
assign micromatriz[44][82] = 9'b110111111;
assign micromatriz[44][83] = 9'b101001001;
assign micromatriz[44][84] = 9'b100000000;
assign micromatriz[44][85] = 9'b100100100;
assign micromatriz[44][86] = 9'b111111111;
assign micromatriz[44][87] = 9'b111111111;
assign micromatriz[44][88] = 9'b111111111;
assign micromatriz[44][89] = 9'b111111111;
assign micromatriz[44][90] = 9'b111111111;
assign micromatriz[44][91] = 9'b111111111;
assign micromatriz[44][92] = 9'b111111111;
assign micromatriz[44][93] = 9'b111111111;
assign micromatriz[44][94] = 9'b111111111;
assign micromatriz[44][95] = 9'b111111111;
assign micromatriz[44][96] = 9'b111111111;
assign micromatriz[44][97] = 9'b111111111;
assign micromatriz[44][98] = 9'b111111111;
assign micromatriz[44][99] = 9'b111111111;
assign micromatriz[45][0] = 9'b111111111;
assign micromatriz[45][1] = 9'b111111111;
assign micromatriz[45][2] = 9'b111111111;
assign micromatriz[45][3] = 9'b111111111;
assign micromatriz[45][4] = 9'b111111111;
assign micromatriz[45][5] = 9'b111111111;
assign micromatriz[45][6] = 9'b111111111;
assign micromatriz[45][7] = 9'b111111111;
assign micromatriz[45][8] = 9'b111111111;
assign micromatriz[45][9] = 9'b111111111;
assign micromatriz[45][10] = 9'b111111111;
assign micromatriz[45][11] = 9'b111111111;
assign micromatriz[45][12] = 9'b111111111;
assign micromatriz[45][13] = 9'b111111111;
assign micromatriz[45][14] = 9'b100100100;
assign micromatriz[45][15] = 9'b100000000;
assign micromatriz[45][16] = 9'b101101101;
assign micromatriz[45][17] = 9'b111111111;
assign micromatriz[45][18] = 9'b111111111;
assign micromatriz[45][19] = 9'b111111111;
assign micromatriz[45][20] = 9'b111111111;
assign micromatriz[45][21] = 9'b100101000;
assign micromatriz[45][22] = 9'b100000000;
assign micromatriz[45][23] = 9'b100100100;
assign micromatriz[45][24] = 9'b101101101;
assign micromatriz[45][25] = 9'b101001101;
assign micromatriz[45][26] = 9'b110001101;
assign micromatriz[45][27] = 9'b111111100;
assign micromatriz[45][28] = 9'b111111100;
assign micromatriz[45][29] = 9'b111111100;
assign micromatriz[45][30] = 9'b111111100;
assign micromatriz[45][31] = 9'b111111100;
assign micromatriz[45][32] = 9'b111111100;
assign micromatriz[45][33] = 9'b111111100;
assign micromatriz[45][34] = 9'b111111100;
assign micromatriz[45][35] = 9'b111111100;
assign micromatriz[45][36] = 9'b111111100;
assign micromatriz[45][37] = 9'b111111100;
assign micromatriz[45][38] = 9'b111111100;
assign micromatriz[45][39] = 9'b111111100;
assign micromatriz[45][40] = 9'b111111100;
assign micromatriz[45][41] = 9'b111111100;
assign micromatriz[45][42] = 9'b111111100;
assign micromatriz[45][43] = 9'b111111100;
assign micromatriz[45][44] = 9'b111111100;
assign micromatriz[45][45] = 9'b111111100;
assign micromatriz[45][46] = 9'b111111100;
assign micromatriz[45][47] = 9'b111111100;
assign micromatriz[45][48] = 9'b111111100;
assign micromatriz[45][49] = 9'b111111100;
assign micromatriz[45][50] = 9'b111111100;
assign micromatriz[45][51] = 9'b111111100;
assign micromatriz[45][52] = 9'b111111100;
assign micromatriz[45][53] = 9'b111111100;
assign micromatriz[45][54] = 9'b111111100;
assign micromatriz[45][55] = 9'b111111100;
assign micromatriz[45][56] = 9'b110010001;
assign micromatriz[45][57] = 9'b110010010;
assign micromatriz[45][58] = 9'b110110110;
assign micromatriz[45][59] = 9'b101001001;
assign micromatriz[45][60] = 9'b100000000;
assign micromatriz[45][61] = 9'b100000000;
assign micromatriz[45][62] = 9'b110111111;
assign micromatriz[45][63] = 9'b111111111;
assign micromatriz[45][64] = 9'b110110111;
assign micromatriz[45][65] = 9'b110110111;
assign micromatriz[45][66] = 9'b101101101;
assign micromatriz[45][67] = 9'b100000000;
assign micromatriz[45][68] = 9'b100000000;
assign micromatriz[45][69] = 9'b111111111;
assign micromatriz[45][70] = 9'b111111111;
assign micromatriz[45][71] = 9'b111111111;
assign micromatriz[45][72] = 9'b111111111;
assign micromatriz[45][73] = 9'b110110111;
assign micromatriz[45][74] = 9'b100100100;
assign micromatriz[45][75] = 9'b100100100;
assign micromatriz[45][76] = 9'b100100100;
assign micromatriz[45][77] = 9'b100100100;
assign micromatriz[45][78] = 9'b101001101;
assign micromatriz[45][79] = 9'b111111111;
assign micromatriz[45][80] = 9'b111111111;
assign micromatriz[45][81] = 9'b110110111;
assign micromatriz[45][82] = 9'b110111111;
assign micromatriz[45][83] = 9'b101001001;
assign micromatriz[45][84] = 9'b100000000;
assign micromatriz[45][85] = 9'b100100100;
assign micromatriz[45][86] = 9'b111111111;
assign micromatriz[45][87] = 9'b111111111;
assign micromatriz[45][88] = 9'b111111111;
assign micromatriz[45][89] = 9'b111111111;
assign micromatriz[45][90] = 9'b111111111;
assign micromatriz[45][91] = 9'b111111111;
assign micromatriz[45][92] = 9'b111111111;
assign micromatriz[45][93] = 9'b111111111;
assign micromatriz[45][94] = 9'b111111111;
assign micromatriz[45][95] = 9'b111111111;
assign micromatriz[45][96] = 9'b111111111;
assign micromatriz[45][97] = 9'b111111111;
assign micromatriz[45][98] = 9'b111111111;
assign micromatriz[45][99] = 9'b111111111;
assign micromatriz[46][0] = 9'b111111111;
assign micromatriz[46][1] = 9'b111111111;
assign micromatriz[46][2] = 9'b111111111;
assign micromatriz[46][3] = 9'b111111111;
assign micromatriz[46][4] = 9'b111111111;
assign micromatriz[46][5] = 9'b111111111;
assign micromatriz[46][6] = 9'b111111111;
assign micromatriz[46][7] = 9'b111111111;
assign micromatriz[46][8] = 9'b111111111;
assign micromatriz[46][9] = 9'b111111111;
assign micromatriz[46][10] = 9'b111111111;
assign micromatriz[46][11] = 9'b111111111;
assign micromatriz[46][12] = 9'b111111111;
assign micromatriz[46][13] = 9'b111111111;
assign micromatriz[46][14] = 9'b100100100;
assign micromatriz[46][15] = 9'b100000000;
assign micromatriz[46][16] = 9'b101101101;
assign micromatriz[46][17] = 9'b111111111;
assign micromatriz[46][18] = 9'b111111111;
assign micromatriz[46][19] = 9'b111111111;
assign micromatriz[46][20] = 9'b111111111;
assign micromatriz[46][21] = 9'b100101000;
assign micromatriz[46][22] = 9'b100000000;
assign micromatriz[46][23] = 9'b100100100;
assign micromatriz[46][24] = 9'b101101101;
assign micromatriz[46][25] = 9'b101001101;
assign micromatriz[46][26] = 9'b110001101;
assign micromatriz[46][27] = 9'b111111100;
assign micromatriz[46][28] = 9'b111111100;
assign micromatriz[46][29] = 9'b111111100;
assign micromatriz[46][30] = 9'b111111100;
assign micromatriz[46][31] = 9'b111111100;
assign micromatriz[46][32] = 9'b111111100;
assign micromatriz[46][33] = 9'b111111100;
assign micromatriz[46][34] = 9'b111111100;
assign micromatriz[46][35] = 9'b111111100;
assign micromatriz[46][36] = 9'b111111100;
assign micromatriz[46][37] = 9'b111111100;
assign micromatriz[46][38] = 9'b111111100;
assign micromatriz[46][39] = 9'b111111100;
assign micromatriz[46][40] = 9'b111111100;
assign micromatriz[46][41] = 9'b111111100;
assign micromatriz[46][42] = 9'b111111100;
assign micromatriz[46][43] = 9'b111111100;
assign micromatriz[46][44] = 9'b111111100;
assign micromatriz[46][45] = 9'b111111100;
assign micromatriz[46][46] = 9'b111111100;
assign micromatriz[46][47] = 9'b111111100;
assign micromatriz[46][48] = 9'b111111100;
assign micromatriz[46][49] = 9'b111111100;
assign micromatriz[46][50] = 9'b111111100;
assign micromatriz[46][51] = 9'b111111100;
assign micromatriz[46][52] = 9'b111111100;
assign micromatriz[46][53] = 9'b111111100;
assign micromatriz[46][54] = 9'b111111100;
assign micromatriz[46][55] = 9'b111111100;
assign micromatriz[46][56] = 9'b110010001;
assign micromatriz[46][57] = 9'b110010010;
assign micromatriz[46][58] = 9'b110110110;
assign micromatriz[46][59] = 9'b101001001;
assign micromatriz[46][60] = 9'b100000000;
assign micromatriz[46][61] = 9'b100000000;
assign micromatriz[46][62] = 9'b110111111;
assign micromatriz[46][63] = 9'b111111111;
assign micromatriz[46][64] = 9'b110110111;
assign micromatriz[46][65] = 9'b110110111;
assign micromatriz[46][66] = 9'b101101101;
assign micromatriz[46][67] = 9'b100000000;
assign micromatriz[46][68] = 9'b100000000;
assign micromatriz[46][69] = 9'b111111111;
assign micromatriz[46][70] = 9'b111111111;
assign micromatriz[46][71] = 9'b111111111;
assign micromatriz[46][72] = 9'b111111111;
assign micromatriz[46][73] = 9'b110111111;
assign micromatriz[46][74] = 9'b100000000;
assign micromatriz[46][75] = 9'b100000000;
assign micromatriz[46][76] = 9'b100000000;
assign micromatriz[46][77] = 9'b100000000;
assign micromatriz[46][78] = 9'b100100100;
assign micromatriz[46][79] = 9'b111111111;
assign micromatriz[46][80] = 9'b111111111;
assign micromatriz[46][81] = 9'b110110111;
assign micromatriz[46][82] = 9'b110111111;
assign micromatriz[46][83] = 9'b101001001;
assign micromatriz[46][84] = 9'b100000000;
assign micromatriz[46][85] = 9'b100100100;
assign micromatriz[46][86] = 9'b111111111;
assign micromatriz[46][87] = 9'b111111111;
assign micromatriz[46][88] = 9'b111111111;
assign micromatriz[46][89] = 9'b111111111;
assign micromatriz[46][90] = 9'b111111111;
assign micromatriz[46][91] = 9'b111111111;
assign micromatriz[46][92] = 9'b111111111;
assign micromatriz[46][93] = 9'b111111111;
assign micromatriz[46][94] = 9'b111111111;
assign micromatriz[46][95] = 9'b111111111;
assign micromatriz[46][96] = 9'b111111111;
assign micromatriz[46][97] = 9'b111111111;
assign micromatriz[46][98] = 9'b111111111;
assign micromatriz[46][99] = 9'b111111111;
assign micromatriz[47][0] = 9'b111111111;
assign micromatriz[47][1] = 9'b111111111;
assign micromatriz[47][2] = 9'b111111111;
assign micromatriz[47][3] = 9'b111111111;
assign micromatriz[47][4] = 9'b111111111;
assign micromatriz[47][5] = 9'b111111111;
assign micromatriz[47][6] = 9'b111111111;
assign micromatriz[47][7] = 9'b111111111;
assign micromatriz[47][8] = 9'b111111111;
assign micromatriz[47][9] = 9'b111111111;
assign micromatriz[47][10] = 9'b111111111;
assign micromatriz[47][11] = 9'b111111111;
assign micromatriz[47][12] = 9'b111111111;
assign micromatriz[47][13] = 9'b111111111;
assign micromatriz[47][14] = 9'b100100100;
assign micromatriz[47][15] = 9'b100000000;
assign micromatriz[47][16] = 9'b101101101;
assign micromatriz[47][17] = 9'b111111111;
assign micromatriz[47][18] = 9'b111111111;
assign micromatriz[47][19] = 9'b111111111;
assign micromatriz[47][20] = 9'b111111111;
assign micromatriz[47][21] = 9'b100101000;
assign micromatriz[47][22] = 9'b100000000;
assign micromatriz[47][23] = 9'b100100100;
assign micromatriz[47][24] = 9'b101101101;
assign micromatriz[47][25] = 9'b101001101;
assign micromatriz[47][26] = 9'b110001101;
assign micromatriz[47][27] = 9'b111111100;
assign micromatriz[47][28] = 9'b111111100;
assign micromatriz[47][29] = 9'b111111100;
assign micromatriz[47][30] = 9'b111111100;
assign micromatriz[47][31] = 9'b111111100;
assign micromatriz[47][32] = 9'b111111100;
assign micromatriz[47][33] = 9'b111111100;
assign micromatriz[47][34] = 9'b111111100;
assign micromatriz[47][35] = 9'b111111100;
assign micromatriz[47][36] = 9'b111111100;
assign micromatriz[47][37] = 9'b111111100;
assign micromatriz[47][38] = 9'b111111100;
assign micromatriz[47][39] = 9'b111111100;
assign micromatriz[47][40] = 9'b111111100;
assign micromatriz[47][41] = 9'b111111100;
assign micromatriz[47][42] = 9'b111111100;
assign micromatriz[47][43] = 9'b111111100;
assign micromatriz[47][44] = 9'b111111100;
assign micromatriz[47][45] = 9'b111111100;
assign micromatriz[47][46] = 9'b111111100;
assign micromatriz[47][47] = 9'b111111100;
assign micromatriz[47][48] = 9'b111111100;
assign micromatriz[47][49] = 9'b111111100;
assign micromatriz[47][50] = 9'b111111100;
assign micromatriz[47][51] = 9'b111111100;
assign micromatriz[47][52] = 9'b111111100;
assign micromatriz[47][53] = 9'b111111100;
assign micromatriz[47][54] = 9'b111111100;
assign micromatriz[47][55] = 9'b111111100;
assign micromatriz[47][56] = 9'b110010001;
assign micromatriz[47][57] = 9'b110010010;
assign micromatriz[47][58] = 9'b110110110;
assign micromatriz[47][59] = 9'b101001001;
assign micromatriz[47][60] = 9'b100000000;
assign micromatriz[47][61] = 9'b100000000;
assign micromatriz[47][62] = 9'b110111111;
assign micromatriz[47][63] = 9'b111111111;
assign micromatriz[47][64] = 9'b110110111;
assign micromatriz[47][65] = 9'b110110111;
assign micromatriz[47][66] = 9'b101101101;
assign micromatriz[47][67] = 9'b100000000;
assign micromatriz[47][68] = 9'b100000000;
assign micromatriz[47][69] = 9'b111111111;
assign micromatriz[47][70] = 9'b111111111;
assign micromatriz[47][71] = 9'b110110111;
assign micromatriz[47][72] = 9'b101101101;
assign micromatriz[47][73] = 9'b101101101;
assign micromatriz[47][74] = 9'b101001001;
assign micromatriz[47][75] = 9'b101001001;
assign micromatriz[47][76] = 9'b101001001;
assign micromatriz[47][77] = 9'b101001001;
assign micromatriz[47][78] = 9'b101001001;
assign micromatriz[47][79] = 9'b101101101;
assign micromatriz[47][80] = 9'b101101101;
assign micromatriz[47][81] = 9'b110010110;
assign micromatriz[47][82] = 9'b110111111;
assign micromatriz[47][83] = 9'b101001001;
assign micromatriz[47][84] = 9'b100000000;
assign micromatriz[47][85] = 9'b100100100;
assign micromatriz[47][86] = 9'b111111111;
assign micromatriz[47][87] = 9'b111111111;
assign micromatriz[47][88] = 9'b111111111;
assign micromatriz[47][89] = 9'b111111111;
assign micromatriz[47][90] = 9'b111111111;
assign micromatriz[47][91] = 9'b111111111;
assign micromatriz[47][92] = 9'b111111111;
assign micromatriz[47][93] = 9'b111111111;
assign micromatriz[47][94] = 9'b111111111;
assign micromatriz[47][95] = 9'b111111111;
assign micromatriz[47][96] = 9'b111111111;
assign micromatriz[47][97] = 9'b111111111;
assign micromatriz[47][98] = 9'b111111111;
assign micromatriz[47][99] = 9'b111111111;
assign micromatriz[48][0] = 9'b111111111;
assign micromatriz[48][1] = 9'b111111111;
assign micromatriz[48][2] = 9'b111111111;
assign micromatriz[48][3] = 9'b111111111;
assign micromatriz[48][4] = 9'b111111111;
assign micromatriz[48][5] = 9'b111111111;
assign micromatriz[48][6] = 9'b111111111;
assign micromatriz[48][7] = 9'b111111111;
assign micromatriz[48][8] = 9'b111111111;
assign micromatriz[48][9] = 9'b111111111;
assign micromatriz[48][10] = 9'b111111111;
assign micromatriz[48][11] = 9'b111111111;
assign micromatriz[48][12] = 9'b111111111;
assign micromatriz[48][13] = 9'b111111111;
assign micromatriz[48][14] = 9'b100100100;
assign micromatriz[48][15] = 9'b100000000;
assign micromatriz[48][16] = 9'b101101101;
assign micromatriz[48][17] = 9'b111111111;
assign micromatriz[48][18] = 9'b111111111;
assign micromatriz[48][19] = 9'b111111111;
assign micromatriz[48][20] = 9'b111111111;
assign micromatriz[48][21] = 9'b100101000;
assign micromatriz[48][22] = 9'b100000000;
assign micromatriz[48][23] = 9'b100100100;
assign micromatriz[48][24] = 9'b101101101;
assign micromatriz[48][25] = 9'b101001101;
assign micromatriz[48][26] = 9'b110001101;
assign micromatriz[48][27] = 9'b111111100;
assign micromatriz[48][28] = 9'b111111100;
assign micromatriz[48][29] = 9'b111111100;
assign micromatriz[48][30] = 9'b111111100;
assign micromatriz[48][31] = 9'b111111100;
assign micromatriz[48][32] = 9'b111111100;
assign micromatriz[48][33] = 9'b111111100;
assign micromatriz[48][34] = 9'b111111100;
assign micromatriz[48][35] = 9'b111111100;
assign micromatriz[48][36] = 9'b111111100;
assign micromatriz[48][37] = 9'b111111100;
assign micromatriz[48][38] = 9'b111111100;
assign micromatriz[48][39] = 9'b111111100;
assign micromatriz[48][40] = 9'b111111100;
assign micromatriz[48][41] = 9'b111111100;
assign micromatriz[48][42] = 9'b111111100;
assign micromatriz[48][43] = 9'b111111100;
assign micromatriz[48][44] = 9'b111111100;
assign micromatriz[48][45] = 9'b111111100;
assign micromatriz[48][46] = 9'b111111100;
assign micromatriz[48][47] = 9'b111111100;
assign micromatriz[48][48] = 9'b111111100;
assign micromatriz[48][49] = 9'b111111100;
assign micromatriz[48][50] = 9'b111111100;
assign micromatriz[48][51] = 9'b111111100;
assign micromatriz[48][52] = 9'b111111100;
assign micromatriz[48][53] = 9'b111111100;
assign micromatriz[48][54] = 9'b111111100;
assign micromatriz[48][55] = 9'b111111100;
assign micromatriz[48][56] = 9'b110010001;
assign micromatriz[48][57] = 9'b110010010;
assign micromatriz[48][58] = 9'b110110110;
assign micromatriz[48][59] = 9'b101001001;
assign micromatriz[48][60] = 9'b100000000;
assign micromatriz[48][61] = 9'b100000000;
assign micromatriz[48][62] = 9'b110111111;
assign micromatriz[48][63] = 9'b111111111;
assign micromatriz[48][64] = 9'b110110111;
assign micromatriz[48][65] = 9'b110110111;
assign micromatriz[48][66] = 9'b101101101;
assign micromatriz[48][67] = 9'b100000000;
assign micromatriz[48][68] = 9'b100000000;
assign micromatriz[48][69] = 9'b111111111;
assign micromatriz[48][70] = 9'b111111111;
assign micromatriz[48][71] = 9'b101101101;
assign micromatriz[48][72] = 9'b100000000;
assign micromatriz[48][73] = 9'b100000000;
assign micromatriz[48][74] = 9'b111111111;
assign micromatriz[48][75] = 9'b111111111;
assign micromatriz[48][76] = 9'b111111111;
assign micromatriz[48][77] = 9'b111111111;
assign micromatriz[48][78] = 9'b110010010;
assign micromatriz[48][79] = 9'b100000000;
assign micromatriz[48][80] = 9'b100000000;
assign micromatriz[48][81] = 9'b110010010;
assign micromatriz[48][82] = 9'b111111111;
assign micromatriz[48][83] = 9'b101001001;
assign micromatriz[48][84] = 9'b100000000;
assign micromatriz[48][85] = 9'b100100100;
assign micromatriz[48][86] = 9'b111111111;
assign micromatriz[48][87] = 9'b111111111;
assign micromatriz[48][88] = 9'b111111111;
assign micromatriz[48][89] = 9'b111111111;
assign micromatriz[48][90] = 9'b111111111;
assign micromatriz[48][91] = 9'b111111111;
assign micromatriz[48][92] = 9'b111111111;
assign micromatriz[48][93] = 9'b111111111;
assign micromatriz[48][94] = 9'b111111111;
assign micromatriz[48][95] = 9'b111111111;
assign micromatriz[48][96] = 9'b111111111;
assign micromatriz[48][97] = 9'b111111111;
assign micromatriz[48][98] = 9'b111111111;
assign micromatriz[48][99] = 9'b111111111;
assign micromatriz[49][0] = 9'b111111111;
assign micromatriz[49][1] = 9'b111111111;
assign micromatriz[49][2] = 9'b111111111;
assign micromatriz[49][3] = 9'b111111111;
assign micromatriz[49][4] = 9'b111111111;
assign micromatriz[49][5] = 9'b111111111;
assign micromatriz[49][6] = 9'b111111111;
assign micromatriz[49][7] = 9'b111111111;
assign micromatriz[49][8] = 9'b111111111;
assign micromatriz[49][9] = 9'b111111111;
assign micromatriz[49][10] = 9'b111111111;
assign micromatriz[49][11] = 9'b111111111;
assign micromatriz[49][12] = 9'b111111111;
assign micromatriz[49][13] = 9'b111111111;
assign micromatriz[49][14] = 9'b100100100;
assign micromatriz[49][15] = 9'b100000000;
assign micromatriz[49][16] = 9'b101101101;
assign micromatriz[49][17] = 9'b111111111;
assign micromatriz[49][18] = 9'b111111111;
assign micromatriz[49][19] = 9'b111111111;
assign micromatriz[49][20] = 9'b111111111;
assign micromatriz[49][21] = 9'b100101000;
assign micromatriz[49][22] = 9'b100000000;
assign micromatriz[49][23] = 9'b100100100;
assign micromatriz[49][24] = 9'b101101101;
assign micromatriz[49][25] = 9'b101001101;
assign micromatriz[49][26] = 9'b110001101;
assign micromatriz[49][27] = 9'b111111100;
assign micromatriz[49][28] = 9'b111111100;
assign micromatriz[49][29] = 9'b111111100;
assign micromatriz[49][30] = 9'b111111100;
assign micromatriz[49][31] = 9'b111111100;
assign micromatriz[49][32] = 9'b111111100;
assign micromatriz[49][33] = 9'b111111100;
assign micromatriz[49][34] = 9'b111111100;
assign micromatriz[49][35] = 9'b111111100;
assign micromatriz[49][36] = 9'b111111100;
assign micromatriz[49][37] = 9'b111111100;
assign micromatriz[49][38] = 9'b111111100;
assign micromatriz[49][39] = 9'b111111100;
assign micromatriz[49][40] = 9'b111111100;
assign micromatriz[49][41] = 9'b111111100;
assign micromatriz[49][42] = 9'b111111100;
assign micromatriz[49][43] = 9'b111111100;
assign micromatriz[49][44] = 9'b111111100;
assign micromatriz[49][45] = 9'b111111100;
assign micromatriz[49][46] = 9'b111111100;
assign micromatriz[49][47] = 9'b111111100;
assign micromatriz[49][48] = 9'b111111100;
assign micromatriz[49][49] = 9'b111111100;
assign micromatriz[49][50] = 9'b111111100;
assign micromatriz[49][51] = 9'b111111100;
assign micromatriz[49][52] = 9'b111111100;
assign micromatriz[49][53] = 9'b111111100;
assign micromatriz[49][54] = 9'b111111100;
assign micromatriz[49][55] = 9'b111111100;
assign micromatriz[49][56] = 9'b110010001;
assign micromatriz[49][57] = 9'b110010010;
assign micromatriz[49][58] = 9'b110110110;
assign micromatriz[49][59] = 9'b101001001;
assign micromatriz[49][60] = 9'b100000000;
assign micromatriz[49][61] = 9'b100000000;
assign micromatriz[49][62] = 9'b110111111;
assign micromatriz[49][63] = 9'b111111111;
assign micromatriz[49][64] = 9'b110110111;
assign micromatriz[49][65] = 9'b110110111;
assign micromatriz[49][66] = 9'b101101101;
assign micromatriz[49][67] = 9'b100000000;
assign micromatriz[49][68] = 9'b100000000;
assign micromatriz[49][69] = 9'b111111111;
assign micromatriz[49][70] = 9'b111111111;
assign micromatriz[49][71] = 9'b101101101;
assign micromatriz[49][72] = 9'b100000000;
assign micromatriz[49][73] = 9'b100000100;
assign micromatriz[49][74] = 9'b111111111;
assign micromatriz[49][75] = 9'b111111111;
assign micromatriz[49][76] = 9'b111111111;
assign micromatriz[49][77] = 9'b111111111;
assign micromatriz[49][78] = 9'b110010001;
assign micromatriz[49][79] = 9'b100000000;
assign micromatriz[49][80] = 9'b100000000;
assign micromatriz[49][81] = 9'b110010010;
assign micromatriz[49][82] = 9'b111111111;
assign micromatriz[49][83] = 9'b101001001;
assign micromatriz[49][84] = 9'b100000000;
assign micromatriz[49][85] = 9'b100100100;
assign micromatriz[49][86] = 9'b111111111;
assign micromatriz[49][87] = 9'b111111111;
assign micromatriz[49][88] = 9'b111111111;
assign micromatriz[49][89] = 9'b111111111;
assign micromatriz[49][90] = 9'b111111111;
assign micromatriz[49][91] = 9'b111111111;
assign micromatriz[49][92] = 9'b111111111;
assign micromatriz[49][93] = 9'b111111111;
assign micromatriz[49][94] = 9'b111111111;
assign micromatriz[49][95] = 9'b111111111;
assign micromatriz[49][96] = 9'b111111111;
assign micromatriz[49][97] = 9'b111111111;
assign micromatriz[49][98] = 9'b111111111;
assign micromatriz[49][99] = 9'b111111111;
assign micromatriz[50][0] = 9'b111111111;
assign micromatriz[50][1] = 9'b111111111;
assign micromatriz[50][2] = 9'b111111111;
assign micromatriz[50][3] = 9'b111111111;
assign micromatriz[50][4] = 9'b111111111;
assign micromatriz[50][5] = 9'b111111111;
assign micromatriz[50][6] = 9'b111111111;
assign micromatriz[50][7] = 9'b111111111;
assign micromatriz[50][8] = 9'b111111111;
assign micromatriz[50][9] = 9'b111111111;
assign micromatriz[50][10] = 9'b111111111;
assign micromatriz[50][11] = 9'b111111111;
assign micromatriz[50][12] = 9'b111111111;
assign micromatriz[50][13] = 9'b111111111;
assign micromatriz[50][14] = 9'b100100100;
assign micromatriz[50][15] = 9'b100000000;
assign micromatriz[50][16] = 9'b101101101;
assign micromatriz[50][17] = 9'b111111111;
assign micromatriz[50][18] = 9'b111111111;
assign micromatriz[50][19] = 9'b111111111;
assign micromatriz[50][20] = 9'b111111111;
assign micromatriz[50][21] = 9'b100101000;
assign micromatriz[50][22] = 9'b100000000;
assign micromatriz[50][23] = 9'b100100100;
assign micromatriz[50][24] = 9'b101101101;
assign micromatriz[50][25] = 9'b101001101;
assign micromatriz[50][26] = 9'b110001101;
assign micromatriz[50][27] = 9'b111111100;
assign micromatriz[50][28] = 9'b111111100;
assign micromatriz[50][29] = 9'b111111100;
assign micromatriz[50][30] = 9'b111111100;
assign micromatriz[50][31] = 9'b111111100;
assign micromatriz[50][32] = 9'b111111100;
assign micromatriz[50][33] = 9'b111111100;
assign micromatriz[50][34] = 9'b111111100;
assign micromatriz[50][35] = 9'b111111100;
assign micromatriz[50][36] = 9'b111111100;
assign micromatriz[50][37] = 9'b111111100;
assign micromatriz[50][38] = 9'b111111100;
assign micromatriz[50][39] = 9'b111111100;
assign micromatriz[50][40] = 9'b111111100;
assign micromatriz[50][41] = 9'b111111100;
assign micromatriz[50][42] = 9'b111111100;
assign micromatriz[50][43] = 9'b111111100;
assign micromatriz[50][44] = 9'b111111100;
assign micromatriz[50][45] = 9'b111111100;
assign micromatriz[50][46] = 9'b111111100;
assign micromatriz[50][47] = 9'b111111100;
assign micromatriz[50][48] = 9'b111111100;
assign micromatriz[50][49] = 9'b111111100;
assign micromatriz[50][50] = 9'b111111100;
assign micromatriz[50][51] = 9'b111111100;
assign micromatriz[50][52] = 9'b111111100;
assign micromatriz[50][53] = 9'b111111100;
assign micromatriz[50][54] = 9'b111111100;
assign micromatriz[50][55] = 9'b111111100;
assign micromatriz[50][56] = 9'b110010001;
assign micromatriz[50][57] = 9'b110010010;
assign micromatriz[50][58] = 9'b110110110;
assign micromatriz[50][59] = 9'b101001001;
assign micromatriz[50][60] = 9'b100000000;
assign micromatriz[50][61] = 9'b100000000;
assign micromatriz[50][62] = 9'b110111111;
assign micromatriz[50][63] = 9'b111111111;
assign micromatriz[50][64] = 9'b110110111;
assign micromatriz[50][65] = 9'b110110111;
assign micromatriz[50][66] = 9'b101101101;
assign micromatriz[50][67] = 9'b100000000;
assign micromatriz[50][68] = 9'b100000000;
assign micromatriz[50][69] = 9'b111111111;
assign micromatriz[50][70] = 9'b111111111;
assign micromatriz[50][71] = 9'b101101101;
assign micromatriz[50][72] = 9'b100000000;
assign micromatriz[50][73] = 9'b100000000;
assign micromatriz[50][74] = 9'b111111111;
assign micromatriz[50][75] = 9'b111111111;
assign micromatriz[50][76] = 9'b110110111;
assign micromatriz[50][77] = 9'b110111111;
assign micromatriz[50][78] = 9'b101101101;
assign micromatriz[50][79] = 9'b100000000;
assign micromatriz[50][80] = 9'b100000000;
assign micromatriz[50][81] = 9'b110010010;
assign micromatriz[50][82] = 9'b111111111;
assign micromatriz[50][83] = 9'b101001001;
assign micromatriz[50][84] = 9'b100000000;
assign micromatriz[50][85] = 9'b100100100;
assign micromatriz[50][86] = 9'b111111111;
assign micromatriz[50][87] = 9'b111111111;
assign micromatriz[50][88] = 9'b111111111;
assign micromatriz[50][89] = 9'b111111111;
assign micromatriz[50][90] = 9'b111111111;
assign micromatriz[50][91] = 9'b111111111;
assign micromatriz[50][92] = 9'b111111111;
assign micromatriz[50][93] = 9'b111111111;
assign micromatriz[50][94] = 9'b111111111;
assign micromatriz[50][95] = 9'b111111111;
assign micromatriz[50][96] = 9'b111111111;
assign micromatriz[50][97] = 9'b111111111;
assign micromatriz[50][98] = 9'b111111111;
assign micromatriz[50][99] = 9'b111111111;
assign micromatriz[51][0] = 9'b111111111;
assign micromatriz[51][1] = 9'b111111111;
assign micromatriz[51][2] = 9'b111111111;
assign micromatriz[51][3] = 9'b111111111;
assign micromatriz[51][4] = 9'b111111111;
assign micromatriz[51][5] = 9'b111111111;
assign micromatriz[51][6] = 9'b111111111;
assign micromatriz[51][7] = 9'b111111111;
assign micromatriz[51][8] = 9'b111111111;
assign micromatriz[51][9] = 9'b111111111;
assign micromatriz[51][10] = 9'b111111111;
assign micromatriz[51][11] = 9'b111111111;
assign micromatriz[51][12] = 9'b111111111;
assign micromatriz[51][13] = 9'b111111111;
assign micromatriz[51][14] = 9'b100100100;
assign micromatriz[51][15] = 9'b100000000;
assign micromatriz[51][16] = 9'b101101101;
assign micromatriz[51][17] = 9'b111111111;
assign micromatriz[51][18] = 9'b111111111;
assign micromatriz[51][19] = 9'b111111111;
assign micromatriz[51][20] = 9'b111111111;
assign micromatriz[51][21] = 9'b100101000;
assign micromatriz[51][22] = 9'b100000000;
assign micromatriz[51][23] = 9'b100100100;
assign micromatriz[51][24] = 9'b101101101;
assign micromatriz[51][25] = 9'b101001101;
assign micromatriz[51][26] = 9'b110001101;
assign micromatriz[51][27] = 9'b111111100;
assign micromatriz[51][28] = 9'b111111100;
assign micromatriz[51][29] = 9'b111111100;
assign micromatriz[51][30] = 9'b111111100;
assign micromatriz[51][31] = 9'b111111100;
assign micromatriz[51][32] = 9'b111111100;
assign micromatriz[51][33] = 9'b111111100;
assign micromatriz[51][34] = 9'b111111100;
assign micromatriz[51][35] = 9'b111111100;
assign micromatriz[51][36] = 9'b111111100;
assign micromatriz[51][37] = 9'b111111100;
assign micromatriz[51][38] = 9'b111111100;
assign micromatriz[51][39] = 9'b111111100;
assign micromatriz[51][40] = 9'b111111100;
assign micromatriz[51][41] = 9'b111111100;
assign micromatriz[51][42] = 9'b111111100;
assign micromatriz[51][43] = 9'b111111100;
assign micromatriz[51][44] = 9'b111111100;
assign micromatriz[51][45] = 9'b111111100;
assign micromatriz[51][46] = 9'b111111100;
assign micromatriz[51][47] = 9'b111111100;
assign micromatriz[51][48] = 9'b111111100;
assign micromatriz[51][49] = 9'b111111100;
assign micromatriz[51][50] = 9'b111111100;
assign micromatriz[51][51] = 9'b111111100;
assign micromatriz[51][52] = 9'b111111100;
assign micromatriz[51][53] = 9'b111111100;
assign micromatriz[51][54] = 9'b111111100;
assign micromatriz[51][55] = 9'b111111100;
assign micromatriz[51][56] = 9'b110010001;
assign micromatriz[51][57] = 9'b110010010;
assign micromatriz[51][58] = 9'b110110110;
assign micromatriz[51][59] = 9'b101001001;
assign micromatriz[51][60] = 9'b100000000;
assign micromatriz[51][61] = 9'b100000000;
assign micromatriz[51][62] = 9'b110111111;
assign micromatriz[51][63] = 9'b111111111;
assign micromatriz[51][64] = 9'b110110111;
assign micromatriz[51][65] = 9'b110110111;
assign micromatriz[51][66] = 9'b101101101;
assign micromatriz[51][67] = 9'b100000000;
assign micromatriz[51][68] = 9'b100000000;
assign micromatriz[51][69] = 9'b111111111;
assign micromatriz[51][70] = 9'b111111111;
assign micromatriz[51][71] = 9'b101101101;
assign micromatriz[51][72] = 9'b100000000;
assign micromatriz[51][73] = 9'b100000000;
assign micromatriz[51][74] = 9'b111111111;
assign micromatriz[51][75] = 9'b111111111;
assign micromatriz[51][76] = 9'b111111111;
assign micromatriz[51][77] = 9'b111111111;
assign micromatriz[51][78] = 9'b101101101;
assign micromatriz[51][79] = 9'b100000000;
assign micromatriz[51][80] = 9'b100000000;
assign micromatriz[51][81] = 9'b110010010;
assign micromatriz[51][82] = 9'b111111111;
assign micromatriz[51][83] = 9'b101001001;
assign micromatriz[51][84] = 9'b100000000;
assign micromatriz[51][85] = 9'b100100100;
assign micromatriz[51][86] = 9'b111111111;
assign micromatriz[51][87] = 9'b111111111;
assign micromatriz[51][88] = 9'b111111111;
assign micromatriz[51][89] = 9'b111111111;
assign micromatriz[51][90] = 9'b111111111;
assign micromatriz[51][91] = 9'b111111111;
assign micromatriz[51][92] = 9'b111111111;
assign micromatriz[51][93] = 9'b111111111;
assign micromatriz[51][94] = 9'b111111111;
assign micromatriz[51][95] = 9'b111111111;
assign micromatriz[51][96] = 9'b111111111;
assign micromatriz[51][97] = 9'b111111111;
assign micromatriz[51][98] = 9'b111111111;
assign micromatriz[51][99] = 9'b111111111;
assign micromatriz[52][0] = 9'b111111111;
assign micromatriz[52][1] = 9'b111111111;
assign micromatriz[52][2] = 9'b111111111;
assign micromatriz[52][3] = 9'b111111111;
assign micromatriz[52][4] = 9'b111111111;
assign micromatriz[52][5] = 9'b111111111;
assign micromatriz[52][6] = 9'b111111111;
assign micromatriz[52][7] = 9'b111111111;
assign micromatriz[52][8] = 9'b111111111;
assign micromatriz[52][9] = 9'b111111111;
assign micromatriz[52][10] = 9'b111111111;
assign micromatriz[52][11] = 9'b111111111;
assign micromatriz[52][12] = 9'b111111111;
assign micromatriz[52][13] = 9'b111111111;
assign micromatriz[52][14] = 9'b100100100;
assign micromatriz[52][15] = 9'b100000000;
assign micromatriz[52][16] = 9'b101101101;
assign micromatriz[52][17] = 9'b111111111;
assign micromatriz[52][18] = 9'b111111111;
assign micromatriz[52][19] = 9'b111111111;
assign micromatriz[52][20] = 9'b111111111;
assign micromatriz[52][21] = 9'b100101000;
assign micromatriz[52][22] = 9'b100000000;
assign micromatriz[52][23] = 9'b100100100;
assign micromatriz[52][24] = 9'b101101101;
assign micromatriz[52][25] = 9'b101001101;
assign micromatriz[52][26] = 9'b110001101;
assign micromatriz[52][27] = 9'b111111100;
assign micromatriz[52][28] = 9'b111111100;
assign micromatriz[52][29] = 9'b111111100;
assign micromatriz[52][30] = 9'b111111100;
assign micromatriz[52][31] = 9'b111111100;
assign micromatriz[52][32] = 9'b111111100;
assign micromatriz[52][33] = 9'b111111100;
assign micromatriz[52][34] = 9'b111111100;
assign micromatriz[52][35] = 9'b111111100;
assign micromatriz[52][36] = 9'b111111100;
assign micromatriz[52][37] = 9'b111111100;
assign micromatriz[52][38] = 9'b111111100;
assign micromatriz[52][39] = 9'b111111100;
assign micromatriz[52][40] = 9'b111111100;
assign micromatriz[52][41] = 9'b111111100;
assign micromatriz[52][42] = 9'b111111100;
assign micromatriz[52][43] = 9'b111111100;
assign micromatriz[52][44] = 9'b111111100;
assign micromatriz[52][45] = 9'b111111100;
assign micromatriz[52][46] = 9'b111111100;
assign micromatriz[52][47] = 9'b111111100;
assign micromatriz[52][48] = 9'b111111100;
assign micromatriz[52][49] = 9'b111111100;
assign micromatriz[52][50] = 9'b111111100;
assign micromatriz[52][51] = 9'b111111100;
assign micromatriz[52][52] = 9'b111111100;
assign micromatriz[52][53] = 9'b111111100;
assign micromatriz[52][54] = 9'b111111100;
assign micromatriz[52][55] = 9'b111111100;
assign micromatriz[52][56] = 9'b110010001;
assign micromatriz[52][57] = 9'b110010010;
assign micromatriz[52][58] = 9'b110110110;
assign micromatriz[52][59] = 9'b101001001;
assign micromatriz[52][60] = 9'b100000000;
assign micromatriz[52][61] = 9'b100000000;
assign micromatriz[52][62] = 9'b110111111;
assign micromatriz[52][63] = 9'b111111111;
assign micromatriz[52][64] = 9'b110110111;
assign micromatriz[52][65] = 9'b110110111;
assign micromatriz[52][66] = 9'b101101101;
assign micromatriz[52][67] = 9'b100000000;
assign micromatriz[52][68] = 9'b100000000;
assign micromatriz[52][69] = 9'b111111111;
assign micromatriz[52][70] = 9'b111111111;
assign micromatriz[52][71] = 9'b110110111;
assign micromatriz[52][72] = 9'b101101101;
assign micromatriz[52][73] = 9'b101101101;
assign micromatriz[52][74] = 9'b101001001;
assign micromatriz[52][75] = 9'b101001001;
assign micromatriz[52][76] = 9'b101001001;
assign micromatriz[52][77] = 9'b101001000;
assign micromatriz[52][78] = 9'b101001001;
assign micromatriz[52][79] = 9'b101101101;
assign micromatriz[52][80] = 9'b101101101;
assign micromatriz[52][81] = 9'b110010110;
assign micromatriz[52][82] = 9'b110111111;
assign micromatriz[52][83] = 9'b101001001;
assign micromatriz[52][84] = 9'b100000000;
assign micromatriz[52][85] = 9'b100100100;
assign micromatriz[52][86] = 9'b111111111;
assign micromatriz[52][87] = 9'b111111111;
assign micromatriz[52][88] = 9'b111111111;
assign micromatriz[52][89] = 9'b111111111;
assign micromatriz[52][90] = 9'b111111111;
assign micromatriz[52][91] = 9'b111111111;
assign micromatriz[52][92] = 9'b111111111;
assign micromatriz[52][93] = 9'b111111111;
assign micromatriz[52][94] = 9'b111111111;
assign micromatriz[52][95] = 9'b111111111;
assign micromatriz[52][96] = 9'b111111111;
assign micromatriz[52][97] = 9'b111111111;
assign micromatriz[52][98] = 9'b111111111;
assign micromatriz[52][99] = 9'b111111111;
assign micromatriz[53][0] = 9'b111111111;
assign micromatriz[53][1] = 9'b111111111;
assign micromatriz[53][2] = 9'b111111111;
assign micromatriz[53][3] = 9'b111111111;
assign micromatriz[53][4] = 9'b111111111;
assign micromatriz[53][5] = 9'b111111111;
assign micromatriz[53][6] = 9'b111111111;
assign micromatriz[53][7] = 9'b111111111;
assign micromatriz[53][8] = 9'b111111111;
assign micromatriz[53][9] = 9'b111111111;
assign micromatriz[53][10] = 9'b111111111;
assign micromatriz[53][11] = 9'b111111111;
assign micromatriz[53][12] = 9'b111111111;
assign micromatriz[53][13] = 9'b111111111;
assign micromatriz[53][14] = 9'b100100100;
assign micromatriz[53][15] = 9'b100000000;
assign micromatriz[53][16] = 9'b101101101;
assign micromatriz[53][17] = 9'b111111111;
assign micromatriz[53][18] = 9'b111111111;
assign micromatriz[53][19] = 9'b111111111;
assign micromatriz[53][20] = 9'b111111111;
assign micromatriz[53][21] = 9'b100101000;
assign micromatriz[53][22] = 9'b100000000;
assign micromatriz[53][23] = 9'b100100100;
assign micromatriz[53][24] = 9'b101101101;
assign micromatriz[53][25] = 9'b101001101;
assign micromatriz[53][26] = 9'b110001101;
assign micromatriz[53][27] = 9'b111111100;
assign micromatriz[53][28] = 9'b111111100;
assign micromatriz[53][29] = 9'b111111100;
assign micromatriz[53][30] = 9'b111111100;
assign micromatriz[53][31] = 9'b111111100;
assign micromatriz[53][32] = 9'b111111100;
assign micromatriz[53][33] = 9'b111111100;
assign micromatriz[53][34] = 9'b111111100;
assign micromatriz[53][35] = 9'b111111100;
assign micromatriz[53][36] = 9'b111111100;
assign micromatriz[53][37] = 9'b111111100;
assign micromatriz[53][38] = 9'b111111100;
assign micromatriz[53][39] = 9'b111111100;
assign micromatriz[53][40] = 9'b111111100;
assign micromatriz[53][41] = 9'b111111100;
assign micromatriz[53][42] = 9'b111111100;
assign micromatriz[53][43] = 9'b111111100;
assign micromatriz[53][44] = 9'b111111100;
assign micromatriz[53][45] = 9'b111111100;
assign micromatriz[53][46] = 9'b111111100;
assign micromatriz[53][47] = 9'b111111100;
assign micromatriz[53][48] = 9'b111111100;
assign micromatriz[53][49] = 9'b111111100;
assign micromatriz[53][50] = 9'b111111100;
assign micromatriz[53][51] = 9'b111111100;
assign micromatriz[53][52] = 9'b111111100;
assign micromatriz[53][53] = 9'b111111100;
assign micromatriz[53][54] = 9'b111111100;
assign micromatriz[53][55] = 9'b111111100;
assign micromatriz[53][56] = 9'b110010001;
assign micromatriz[53][57] = 9'b110010010;
assign micromatriz[53][58] = 9'b110110110;
assign micromatriz[53][59] = 9'b101001001;
assign micromatriz[53][60] = 9'b100000000;
assign micromatriz[53][61] = 9'b100000000;
assign micromatriz[53][62] = 9'b110111111;
assign micromatriz[53][63] = 9'b111111111;
assign micromatriz[53][64] = 9'b110110111;
assign micromatriz[53][65] = 9'b110110111;
assign micromatriz[53][66] = 9'b101101101;
assign micromatriz[53][67] = 9'b100000000;
assign micromatriz[53][68] = 9'b100000000;
assign micromatriz[53][69] = 9'b111111111;
assign micromatriz[53][70] = 9'b111111111;
assign micromatriz[53][71] = 9'b111111111;
assign micromatriz[53][72] = 9'b111111111;
assign micromatriz[53][73] = 9'b110111111;
assign micromatriz[53][74] = 9'b100000000;
assign micromatriz[53][75] = 9'b100000000;
assign micromatriz[53][76] = 9'b100000000;
assign micromatriz[53][77] = 9'b100000000;
assign micromatriz[53][78] = 9'b100100100;
assign micromatriz[53][79] = 9'b111111111;
assign micromatriz[53][80] = 9'b111111111;
assign micromatriz[53][81] = 9'b110110111;
assign micromatriz[53][82] = 9'b110111111;
assign micromatriz[53][83] = 9'b101001001;
assign micromatriz[53][84] = 9'b100000000;
assign micromatriz[53][85] = 9'b100100100;
assign micromatriz[53][86] = 9'b111111111;
assign micromatriz[53][87] = 9'b111111111;
assign micromatriz[53][88] = 9'b111111111;
assign micromatriz[53][89] = 9'b111111111;
assign micromatriz[53][90] = 9'b111111111;
assign micromatriz[53][91] = 9'b111111111;
assign micromatriz[53][92] = 9'b111111111;
assign micromatriz[53][93] = 9'b111111111;
assign micromatriz[53][94] = 9'b111111111;
assign micromatriz[53][95] = 9'b111111111;
assign micromatriz[53][96] = 9'b111111111;
assign micromatriz[53][97] = 9'b111111111;
assign micromatriz[53][98] = 9'b111111111;
assign micromatriz[53][99] = 9'b111111111;
assign micromatriz[54][0] = 9'b111111111;
assign micromatriz[54][1] = 9'b111111111;
assign micromatriz[54][2] = 9'b111111111;
assign micromatriz[54][3] = 9'b111111111;
assign micromatriz[54][4] = 9'b111111111;
assign micromatriz[54][5] = 9'b111111111;
assign micromatriz[54][6] = 9'b111111111;
assign micromatriz[54][7] = 9'b111111111;
assign micromatriz[54][8] = 9'b111111111;
assign micromatriz[54][9] = 9'b111111111;
assign micromatriz[54][10] = 9'b111111111;
assign micromatriz[54][11] = 9'b111111111;
assign micromatriz[54][12] = 9'b111111111;
assign micromatriz[54][13] = 9'b111111111;
assign micromatriz[54][14] = 9'b100100100;
assign micromatriz[54][15] = 9'b100000000;
assign micromatriz[54][16] = 9'b101101101;
assign micromatriz[54][17] = 9'b111111111;
assign micromatriz[54][18] = 9'b111111111;
assign micromatriz[54][19] = 9'b111111111;
assign micromatriz[54][20] = 9'b111111111;
assign micromatriz[54][21] = 9'b100101000;
assign micromatriz[54][22] = 9'b100000000;
assign micromatriz[54][23] = 9'b100100100;
assign micromatriz[54][24] = 9'b101101101;
assign micromatriz[54][25] = 9'b101001101;
assign micromatriz[54][26] = 9'b110001101;
assign micromatriz[54][27] = 9'b111111100;
assign micromatriz[54][28] = 9'b111111100;
assign micromatriz[54][29] = 9'b111111100;
assign micromatriz[54][30] = 9'b111111100;
assign micromatriz[54][31] = 9'b111111100;
assign micromatriz[54][32] = 9'b111111100;
assign micromatriz[54][33] = 9'b111111100;
assign micromatriz[54][34] = 9'b111111100;
assign micromatriz[54][35] = 9'b111111100;
assign micromatriz[54][36] = 9'b111111100;
assign micromatriz[54][37] = 9'b111111100;
assign micromatriz[54][38] = 9'b111111100;
assign micromatriz[54][39] = 9'b111111100;
assign micromatriz[54][40] = 9'b111111100;
assign micromatriz[54][41] = 9'b111111100;
assign micromatriz[54][42] = 9'b111111100;
assign micromatriz[54][43] = 9'b111111100;
assign micromatriz[54][44] = 9'b111111100;
assign micromatriz[54][45] = 9'b111111100;
assign micromatriz[54][46] = 9'b111111100;
assign micromatriz[54][47] = 9'b111111100;
assign micromatriz[54][48] = 9'b111111100;
assign micromatriz[54][49] = 9'b111111100;
assign micromatriz[54][50] = 9'b111111100;
assign micromatriz[54][51] = 9'b111111100;
assign micromatriz[54][52] = 9'b111111100;
assign micromatriz[54][53] = 9'b111111100;
assign micromatriz[54][54] = 9'b111111100;
assign micromatriz[54][55] = 9'b111111100;
assign micromatriz[54][56] = 9'b110010001;
assign micromatriz[54][57] = 9'b110010010;
assign micromatriz[54][58] = 9'b110110110;
assign micromatriz[54][59] = 9'b101001001;
assign micromatriz[54][60] = 9'b100000000;
assign micromatriz[54][61] = 9'b100000000;
assign micromatriz[54][62] = 9'b110111111;
assign micromatriz[54][63] = 9'b111111111;
assign micromatriz[54][64] = 9'b110110111;
assign micromatriz[54][65] = 9'b110110111;
assign micromatriz[54][66] = 9'b101101101;
assign micromatriz[54][67] = 9'b100000000;
assign micromatriz[54][68] = 9'b100000000;
assign micromatriz[54][69] = 9'b111111111;
assign micromatriz[54][70] = 9'b111111111;
assign micromatriz[54][71] = 9'b111111111;
assign micromatriz[54][72] = 9'b111111111;
assign micromatriz[54][73] = 9'b110110111;
assign micromatriz[54][74] = 9'b100100100;
assign micromatriz[54][75] = 9'b100100100;
assign micromatriz[54][76] = 9'b100100100;
assign micromatriz[54][77] = 9'b100100100;
assign micromatriz[54][78] = 9'b101001001;
assign micromatriz[54][79] = 9'b111111111;
assign micromatriz[54][80] = 9'b111111111;
assign micromatriz[54][81] = 9'b110110111;
assign micromatriz[54][82] = 9'b110111111;
assign micromatriz[54][83] = 9'b101001001;
assign micromatriz[54][84] = 9'b100000000;
assign micromatriz[54][85] = 9'b100100100;
assign micromatriz[54][86] = 9'b111111111;
assign micromatriz[54][87] = 9'b111111111;
assign micromatriz[54][88] = 9'b111111111;
assign micromatriz[54][89] = 9'b111111111;
assign micromatriz[54][90] = 9'b111111111;
assign micromatriz[54][91] = 9'b111111111;
assign micromatriz[54][92] = 9'b111111111;
assign micromatriz[54][93] = 9'b111111111;
assign micromatriz[54][94] = 9'b111111111;
assign micromatriz[54][95] = 9'b111111111;
assign micromatriz[54][96] = 9'b111111111;
assign micromatriz[54][97] = 9'b111111111;
assign micromatriz[54][98] = 9'b111111111;
assign micromatriz[54][99] = 9'b111111111;
assign micromatriz[55][0] = 9'b111111111;
assign micromatriz[55][1] = 9'b111111111;
assign micromatriz[55][2] = 9'b111111111;
assign micromatriz[55][3] = 9'b111111111;
assign micromatriz[55][4] = 9'b111111111;
assign micromatriz[55][5] = 9'b111111111;
assign micromatriz[55][6] = 9'b111111111;
assign micromatriz[55][7] = 9'b111111111;
assign micromatriz[55][8] = 9'b111111111;
assign micromatriz[55][9] = 9'b111111111;
assign micromatriz[55][10] = 9'b111111111;
assign micromatriz[55][11] = 9'b111111111;
assign micromatriz[55][12] = 9'b111111111;
assign micromatriz[55][13] = 9'b111111111;
assign micromatriz[55][14] = 9'b100100100;
assign micromatriz[55][15] = 9'b100000000;
assign micromatriz[55][16] = 9'b101101101;
assign micromatriz[55][17] = 9'b111111111;
assign micromatriz[55][18] = 9'b111111111;
assign micromatriz[55][19] = 9'b111111111;
assign micromatriz[55][20] = 9'b111111111;
assign micromatriz[55][21] = 9'b100101000;
assign micromatriz[55][22] = 9'b100000000;
assign micromatriz[55][23] = 9'b100100100;
assign micromatriz[55][24] = 9'b101101101;
assign micromatriz[55][25] = 9'b101001101;
assign micromatriz[55][26] = 9'b110010001;
assign micromatriz[55][27] = 9'b111111100;
assign micromatriz[55][28] = 9'b111111100;
assign micromatriz[55][29] = 9'b111111100;
assign micromatriz[55][30] = 9'b111111100;
assign micromatriz[55][31] = 9'b111111100;
assign micromatriz[55][32] = 9'b111111100;
assign micromatriz[55][33] = 9'b111111100;
assign micromatriz[55][34] = 9'b111111100;
assign micromatriz[55][35] = 9'b111111100;
assign micromatriz[55][36] = 9'b111111100;
assign micromatriz[55][37] = 9'b111111100;
assign micromatriz[55][38] = 9'b111111100;
assign micromatriz[55][39] = 9'b111111100;
assign micromatriz[55][40] = 9'b111111100;
assign micromatriz[55][41] = 9'b111111100;
assign micromatriz[55][42] = 9'b111111100;
assign micromatriz[55][43] = 9'b111111100;
assign micromatriz[55][44] = 9'b111111100;
assign micromatriz[55][45] = 9'b111111100;
assign micromatriz[55][46] = 9'b111111100;
assign micromatriz[55][47] = 9'b111111100;
assign micromatriz[55][48] = 9'b111111100;
assign micromatriz[55][49] = 9'b111111100;
assign micromatriz[55][50] = 9'b111111100;
assign micromatriz[55][51] = 9'b111111100;
assign micromatriz[55][52] = 9'b111111100;
assign micromatriz[55][53] = 9'b111111100;
assign micromatriz[55][54] = 9'b111111100;
assign micromatriz[55][55] = 9'b111111100;
assign micromatriz[55][56] = 9'b110010001;
assign micromatriz[55][57] = 9'b110010010;
assign micromatriz[55][58] = 9'b110110110;
assign micromatriz[55][59] = 9'b101001001;
assign micromatriz[55][60] = 9'b100000000;
assign micromatriz[55][61] = 9'b100000000;
assign micromatriz[55][62] = 9'b110111111;
assign micromatriz[55][63] = 9'b111111111;
assign micromatriz[55][64] = 9'b110110111;
assign micromatriz[55][65] = 9'b110110111;
assign micromatriz[55][66] = 9'b101101101;
assign micromatriz[55][67] = 9'b100000000;
assign micromatriz[55][68] = 9'b100000000;
assign micromatriz[55][69] = 9'b111111111;
assign micromatriz[55][70] = 9'b111111111;
assign micromatriz[55][71] = 9'b111111111;
assign micromatriz[55][72] = 9'b111111111;
assign micromatriz[55][73] = 9'b111111111;
assign micromatriz[55][74] = 9'b111111111;
assign micromatriz[55][75] = 9'b111111111;
assign micromatriz[55][76] = 9'b111111111;
assign micromatriz[55][77] = 9'b111111111;
assign micromatriz[55][78] = 9'b111111111;
assign micromatriz[55][79] = 9'b111111111;
assign micromatriz[55][80] = 9'b111111111;
assign micromatriz[55][81] = 9'b110110111;
assign micromatriz[55][82] = 9'b110111111;
assign micromatriz[55][83] = 9'b101001001;
assign micromatriz[55][84] = 9'b100000000;
assign micromatriz[55][85] = 9'b100100100;
assign micromatriz[55][86] = 9'b111111111;
assign micromatriz[55][87] = 9'b111111111;
assign micromatriz[55][88] = 9'b111111111;
assign micromatriz[55][89] = 9'b111111111;
assign micromatriz[55][90] = 9'b111111111;
assign micromatriz[55][91] = 9'b111111111;
assign micromatriz[55][92] = 9'b111111111;
assign micromatriz[55][93] = 9'b111111111;
assign micromatriz[55][94] = 9'b111111111;
assign micromatriz[55][95] = 9'b111111111;
assign micromatriz[55][96] = 9'b111111111;
assign micromatriz[55][97] = 9'b111111111;
assign micromatriz[55][98] = 9'b111111111;
assign micromatriz[55][99] = 9'b111111111;
assign micromatriz[56][0] = 9'b111111111;
assign micromatriz[56][1] = 9'b111111111;
assign micromatriz[56][2] = 9'b111111111;
assign micromatriz[56][3] = 9'b111111111;
assign micromatriz[56][4] = 9'b111111111;
assign micromatriz[56][5] = 9'b111111111;
assign micromatriz[56][6] = 9'b111111111;
assign micromatriz[56][7] = 9'b111111111;
assign micromatriz[56][8] = 9'b111111111;
assign micromatriz[56][9] = 9'b111111111;
assign micromatriz[56][10] = 9'b111111111;
assign micromatriz[56][11] = 9'b111111111;
assign micromatriz[56][12] = 9'b111111111;
assign micromatriz[56][13] = 9'b111111111;
assign micromatriz[56][14] = 9'b100100100;
assign micromatriz[56][15] = 9'b100000000;
assign micromatriz[56][16] = 9'b101101101;
assign micromatriz[56][17] = 9'b111111111;
assign micromatriz[56][18] = 9'b111111111;
assign micromatriz[56][19] = 9'b111111111;
assign micromatriz[56][20] = 9'b111111111;
assign micromatriz[56][21] = 9'b100101000;
assign micromatriz[56][22] = 9'b100000000;
assign micromatriz[56][23] = 9'b100100100;
assign micromatriz[56][24] = 9'b101101101;
assign micromatriz[56][25] = 9'b101101101;
assign micromatriz[56][26] = 9'b101101101;
assign micromatriz[56][27] = 9'b110010001;
assign micromatriz[56][28] = 9'b110010001;
assign micromatriz[56][29] = 9'b110010001;
assign micromatriz[56][30] = 9'b110010001;
assign micromatriz[56][31] = 9'b110010001;
assign micromatriz[56][32] = 9'b110010001;
assign micromatriz[56][33] = 9'b110010001;
assign micromatriz[56][34] = 9'b110010001;
assign micromatriz[56][35] = 9'b110010001;
assign micromatriz[56][36] = 9'b110010001;
assign micromatriz[56][37] = 9'b110010001;
assign micromatriz[56][38] = 9'b110010001;
assign micromatriz[56][39] = 9'b110010001;
assign micromatriz[56][40] = 9'b110010001;
assign micromatriz[56][41] = 9'b110010001;
assign micromatriz[56][42] = 9'b110010001;
assign micromatriz[56][43] = 9'b110010001;
assign micromatriz[56][44] = 9'b110010001;
assign micromatriz[56][45] = 9'b110010001;
assign micromatriz[56][46] = 9'b110010001;
assign micromatriz[56][47] = 9'b110010001;
assign micromatriz[56][48] = 9'b110010001;
assign micromatriz[56][49] = 9'b110010001;
assign micromatriz[56][50] = 9'b110010001;
assign micromatriz[56][51] = 9'b110010001;
assign micromatriz[56][52] = 9'b110010001;
assign micromatriz[56][53] = 9'b110010001;
assign micromatriz[56][54] = 9'b110010001;
assign micromatriz[56][55] = 9'b110010001;
assign micromatriz[56][56] = 9'b101101101;
assign micromatriz[56][57] = 9'b110010001;
assign micromatriz[56][58] = 9'b110110110;
assign micromatriz[56][59] = 9'b101001001;
assign micromatriz[56][60] = 9'b100000000;
assign micromatriz[56][61] = 9'b100000000;
assign micromatriz[56][62] = 9'b110111111;
assign micromatriz[56][63] = 9'b111111111;
assign micromatriz[56][64] = 9'b110110111;
assign micromatriz[56][65] = 9'b110110111;
assign micromatriz[56][66] = 9'b101101101;
assign micromatriz[56][67] = 9'b100000000;
assign micromatriz[56][68] = 9'b100000000;
assign micromatriz[56][69] = 9'b111111111;
assign micromatriz[56][70] = 9'b111111111;
assign micromatriz[56][71] = 9'b111111111;
assign micromatriz[56][72] = 9'b111111111;
assign micromatriz[56][73] = 9'b111111111;
assign micromatriz[56][74] = 9'b111111111;
assign micromatriz[56][75] = 9'b111111111;
assign micromatriz[56][76] = 9'b111111111;
assign micromatriz[56][77] = 9'b111111111;
assign micromatriz[56][78] = 9'b111111111;
assign micromatriz[56][79] = 9'b111111111;
assign micromatriz[56][80] = 9'b111111111;
assign micromatriz[56][81] = 9'b110110111;
assign micromatriz[56][82] = 9'b110111111;
assign micromatriz[56][83] = 9'b101001001;
assign micromatriz[56][84] = 9'b100000000;
assign micromatriz[56][85] = 9'b100100100;
assign micromatriz[56][86] = 9'b111111111;
assign micromatriz[56][87] = 9'b111111111;
assign micromatriz[56][88] = 9'b111111111;
assign micromatriz[56][89] = 9'b111111111;
assign micromatriz[56][90] = 9'b111111111;
assign micromatriz[56][91] = 9'b111111111;
assign micromatriz[56][92] = 9'b111111111;
assign micromatriz[56][93] = 9'b111111111;
assign micromatriz[56][94] = 9'b111111111;
assign micromatriz[56][95] = 9'b111111111;
assign micromatriz[56][96] = 9'b111111111;
assign micromatriz[56][97] = 9'b111111111;
assign micromatriz[56][98] = 9'b111111111;
assign micromatriz[56][99] = 9'b111111111;
assign micromatriz[57][0] = 9'b111111111;
assign micromatriz[57][1] = 9'b111111111;
assign micromatriz[57][2] = 9'b111111111;
assign micromatriz[57][3] = 9'b111111111;
assign micromatriz[57][4] = 9'b111111111;
assign micromatriz[57][5] = 9'b111111111;
assign micromatriz[57][6] = 9'b111111111;
assign micromatriz[57][7] = 9'b111111111;
assign micromatriz[57][8] = 9'b111111111;
assign micromatriz[57][9] = 9'b111111111;
assign micromatriz[57][10] = 9'b111111111;
assign micromatriz[57][11] = 9'b111111111;
assign micromatriz[57][12] = 9'b111111111;
assign micromatriz[57][13] = 9'b111111111;
assign micromatriz[57][14] = 9'b100100100;
assign micromatriz[57][15] = 9'b100000000;
assign micromatriz[57][16] = 9'b101101101;
assign micromatriz[57][17] = 9'b111111111;
assign micromatriz[57][18] = 9'b111111111;
assign micromatriz[57][19] = 9'b111111111;
assign micromatriz[57][20] = 9'b111111111;
assign micromatriz[57][21] = 9'b100101000;
assign micromatriz[57][22] = 9'b100000000;
assign micromatriz[57][23] = 9'b100100100;
assign micromatriz[57][24] = 9'b101101101;
assign micromatriz[57][25] = 9'b101101101;
assign micromatriz[57][26] = 9'b100100100;
assign micromatriz[57][27] = 9'b100000000;
assign micromatriz[57][28] = 9'b100000000;
assign micromatriz[57][29] = 9'b100000000;
assign micromatriz[57][30] = 9'b100000000;
assign micromatriz[57][31] = 9'b100000000;
assign micromatriz[57][32] = 9'b100000000;
assign micromatriz[57][33] = 9'b100000000;
assign micromatriz[57][34] = 9'b100000000;
assign micromatriz[57][35] = 9'b100000000;
assign micromatriz[57][36] = 9'b100000000;
assign micromatriz[57][37] = 9'b100000000;
assign micromatriz[57][38] = 9'b100000000;
assign micromatriz[57][39] = 9'b100000000;
assign micromatriz[57][40] = 9'b100000000;
assign micromatriz[57][41] = 9'b100000000;
assign micromatriz[57][42] = 9'b100000000;
assign micromatriz[57][43] = 9'b100000000;
assign micromatriz[57][44] = 9'b100000000;
assign micromatriz[57][45] = 9'b100000000;
assign micromatriz[57][46] = 9'b100000000;
assign micromatriz[57][47] = 9'b100000000;
assign micromatriz[57][48] = 9'b100000000;
assign micromatriz[57][49] = 9'b100000000;
assign micromatriz[57][50] = 9'b100000000;
assign micromatriz[57][51] = 9'b100000000;
assign micromatriz[57][52] = 9'b100000000;
assign micromatriz[57][53] = 9'b100000000;
assign micromatriz[57][54] = 9'b100000000;
assign micromatriz[57][55] = 9'b100000000;
assign micromatriz[57][56] = 9'b100000000;
assign micromatriz[57][57] = 9'b101101101;
assign micromatriz[57][58] = 9'b110110110;
assign micromatriz[57][59] = 9'b101001001;
assign micromatriz[57][60] = 9'b100000000;
assign micromatriz[57][61] = 9'b100000000;
assign micromatriz[57][62] = 9'b110111111;
assign micromatriz[57][63] = 9'b111111111;
assign micromatriz[57][64] = 9'b110110111;
assign micromatriz[57][65] = 9'b110110111;
assign micromatriz[57][66] = 9'b101101101;
assign micromatriz[57][67] = 9'b100000000;
assign micromatriz[57][68] = 9'b100000000;
assign micromatriz[57][69] = 9'b111111111;
assign micromatriz[57][70] = 9'b111111111;
assign micromatriz[57][71] = 9'b111111111;
assign micromatriz[57][72] = 9'b111111111;
assign micromatriz[57][73] = 9'b110110111;
assign micromatriz[57][74] = 9'b100100100;
assign micromatriz[57][75] = 9'b100100100;
assign micromatriz[57][76] = 9'b100100100;
assign micromatriz[57][77] = 9'b100100100;
assign micromatriz[57][78] = 9'b101001001;
assign micromatriz[57][79] = 9'b111111111;
assign micromatriz[57][80] = 9'b111111111;
assign micromatriz[57][81] = 9'b110110111;
assign micromatriz[57][82] = 9'b110111111;
assign micromatriz[57][83] = 9'b101001001;
assign micromatriz[57][84] = 9'b100000000;
assign micromatriz[57][85] = 9'b100100100;
assign micromatriz[57][86] = 9'b111111111;
assign micromatriz[57][87] = 9'b111111111;
assign micromatriz[57][88] = 9'b111111111;
assign micromatriz[57][89] = 9'b111111111;
assign micromatriz[57][90] = 9'b111111111;
assign micromatriz[57][91] = 9'b111111111;
assign micromatriz[57][92] = 9'b111111111;
assign micromatriz[57][93] = 9'b111111111;
assign micromatriz[57][94] = 9'b111111111;
assign micromatriz[57][95] = 9'b111111111;
assign micromatriz[57][96] = 9'b111111111;
assign micromatriz[57][97] = 9'b111111111;
assign micromatriz[57][98] = 9'b111111111;
assign micromatriz[57][99] = 9'b111111111;
assign micromatriz[58][0] = 9'b111111111;
assign micromatriz[58][1] = 9'b111111111;
assign micromatriz[58][2] = 9'b111111111;
assign micromatriz[58][3] = 9'b111111111;
assign micromatriz[58][4] = 9'b111111111;
assign micromatriz[58][5] = 9'b111111111;
assign micromatriz[58][6] = 9'b111111111;
assign micromatriz[58][7] = 9'b111111111;
assign micromatriz[58][8] = 9'b111111111;
assign micromatriz[58][9] = 9'b111111111;
assign micromatriz[58][10] = 9'b111111111;
assign micromatriz[58][11] = 9'b111111111;
assign micromatriz[58][12] = 9'b111111111;
assign micromatriz[58][13] = 9'b111111111;
assign micromatriz[58][14] = 9'b100100100;
assign micromatriz[58][15] = 9'b100000000;
assign micromatriz[58][16] = 9'b101101101;
assign micromatriz[58][17] = 9'b111111111;
assign micromatriz[58][18] = 9'b111111111;
assign micromatriz[58][19] = 9'b111111111;
assign micromatriz[58][20] = 9'b111111111;
assign micromatriz[58][21] = 9'b100101000;
assign micromatriz[58][22] = 9'b100000000;
assign micromatriz[58][23] = 9'b100100100;
assign micromatriz[58][24] = 9'b101101101;
assign micromatriz[58][25] = 9'b101101101;
assign micromatriz[58][26] = 9'b100000000;
assign micromatriz[58][27] = 9'b100000000;
assign micromatriz[58][28] = 9'b100000000;
assign micromatriz[58][29] = 9'b100000000;
assign micromatriz[58][30] = 9'b100000000;
assign micromatriz[58][31] = 9'b100000000;
assign micromatriz[58][32] = 9'b100000000;
assign micromatriz[58][33] = 9'b100000000;
assign micromatriz[58][34] = 9'b100000000;
assign micromatriz[58][35] = 9'b100000000;
assign micromatriz[58][36] = 9'b100000000;
assign micromatriz[58][37] = 9'b100000000;
assign micromatriz[58][38] = 9'b100000000;
assign micromatriz[58][39] = 9'b100000000;
assign micromatriz[58][40] = 9'b100000000;
assign micromatriz[58][41] = 9'b100000000;
assign micromatriz[58][42] = 9'b100000000;
assign micromatriz[58][43] = 9'b100000000;
assign micromatriz[58][44] = 9'b100000000;
assign micromatriz[58][45] = 9'b100000000;
assign micromatriz[58][46] = 9'b100000000;
assign micromatriz[58][47] = 9'b100000000;
assign micromatriz[58][48] = 9'b100000000;
assign micromatriz[58][49] = 9'b100000000;
assign micromatriz[58][50] = 9'b100000000;
assign micromatriz[58][51] = 9'b100000000;
assign micromatriz[58][52] = 9'b100000000;
assign micromatriz[58][53] = 9'b100000000;
assign micromatriz[58][54] = 9'b100000000;
assign micromatriz[58][55] = 9'b100000000;
assign micromatriz[58][56] = 9'b100000000;
assign micromatriz[58][57] = 9'b101101101;
assign micromatriz[58][58] = 9'b110110110;
assign micromatriz[58][59] = 9'b101001001;
assign micromatriz[58][60] = 9'b100000000;
assign micromatriz[58][61] = 9'b100000000;
assign micromatriz[58][62] = 9'b110111111;
assign micromatriz[58][63] = 9'b111111111;
assign micromatriz[58][64] = 9'b110110111;
assign micromatriz[58][65] = 9'b110110111;
assign micromatriz[58][66] = 9'b101101101;
assign micromatriz[58][67] = 9'b100000000;
assign micromatriz[58][68] = 9'b100000000;
assign micromatriz[58][69] = 9'b111111111;
assign micromatriz[58][70] = 9'b111111111;
assign micromatriz[58][71] = 9'b111111111;
assign micromatriz[58][72] = 9'b111111111;
assign micromatriz[58][73] = 9'b110111111;
assign micromatriz[58][74] = 9'b100000000;
assign micromatriz[58][75] = 9'b100000000;
assign micromatriz[58][76] = 9'b100000000;
assign micromatriz[58][77] = 9'b100000000;
assign micromatriz[58][78] = 9'b100100100;
assign micromatriz[58][79] = 9'b111111111;
assign micromatriz[58][80] = 9'b111111111;
assign micromatriz[58][81] = 9'b110110111;
assign micromatriz[58][82] = 9'b110111111;
assign micromatriz[58][83] = 9'b101001001;
assign micromatriz[58][84] = 9'b100000000;
assign micromatriz[58][85] = 9'b100100100;
assign micromatriz[58][86] = 9'b111111111;
assign micromatriz[58][87] = 9'b111111111;
assign micromatriz[58][88] = 9'b111111111;
assign micromatriz[58][89] = 9'b111111111;
assign micromatriz[58][90] = 9'b111111111;
assign micromatriz[58][91] = 9'b111111111;
assign micromatriz[58][92] = 9'b111111111;
assign micromatriz[58][93] = 9'b111111111;
assign micromatriz[58][94] = 9'b111111111;
assign micromatriz[58][95] = 9'b111111111;
assign micromatriz[58][96] = 9'b111111111;
assign micromatriz[58][97] = 9'b111111111;
assign micromatriz[58][98] = 9'b111111111;
assign micromatriz[58][99] = 9'b111111111;
assign micromatriz[59][0] = 9'b111111111;
assign micromatriz[59][1] = 9'b111111111;
assign micromatriz[59][2] = 9'b111111111;
assign micromatriz[59][3] = 9'b111111111;
assign micromatriz[59][4] = 9'b111111111;
assign micromatriz[59][5] = 9'b111111111;
assign micromatriz[59][6] = 9'b111111111;
assign micromatriz[59][7] = 9'b111111111;
assign micromatriz[59][8] = 9'b111111111;
assign micromatriz[59][9] = 9'b111111111;
assign micromatriz[59][10] = 9'b111111111;
assign micromatriz[59][11] = 9'b111111111;
assign micromatriz[59][12] = 9'b111111111;
assign micromatriz[59][13] = 9'b111111111;
assign micromatriz[59][14] = 9'b100100100;
assign micromatriz[59][15] = 9'b100000000;
assign micromatriz[59][16] = 9'b101101101;
assign micromatriz[59][17] = 9'b111111111;
assign micromatriz[59][18] = 9'b111111111;
assign micromatriz[59][19] = 9'b111111111;
assign micromatriz[59][20] = 9'b111111111;
assign micromatriz[59][21] = 9'b100101000;
assign micromatriz[59][22] = 9'b100000000;
assign micromatriz[59][23] = 9'b100100100;
assign micromatriz[59][24] = 9'b101101101;
assign micromatriz[59][25] = 9'b101101101;
assign micromatriz[59][26] = 9'b101001001;
assign micromatriz[59][27] = 9'b101001000;
assign micromatriz[59][28] = 9'b101001000;
assign micromatriz[59][29] = 9'b101001000;
assign micromatriz[59][30] = 9'b101001000;
assign micromatriz[59][31] = 9'b101001000;
assign micromatriz[59][32] = 9'b101001000;
assign micromatriz[59][33] = 9'b101001000;
assign micromatriz[59][34] = 9'b101001000;
assign micromatriz[59][35] = 9'b101001000;
assign micromatriz[59][36] = 9'b101001000;
assign micromatriz[59][37] = 9'b101001000;
assign micromatriz[59][38] = 9'b101001000;
assign micromatriz[59][39] = 9'b101001000;
assign micromatriz[59][40] = 9'b101001000;
assign micromatriz[59][41] = 9'b101001000;
assign micromatriz[59][42] = 9'b101001000;
assign micromatriz[59][43] = 9'b101001000;
assign micromatriz[59][44] = 9'b101001000;
assign micromatriz[59][45] = 9'b101001000;
assign micromatriz[59][46] = 9'b101001000;
assign micromatriz[59][47] = 9'b101001000;
assign micromatriz[59][48] = 9'b101001000;
assign micromatriz[59][49] = 9'b101001000;
assign micromatriz[59][50] = 9'b101001000;
assign micromatriz[59][51] = 9'b101001000;
assign micromatriz[59][52] = 9'b101001000;
assign micromatriz[59][53] = 9'b101001000;
assign micromatriz[59][54] = 9'b101001000;
assign micromatriz[59][55] = 9'b101001000;
assign micromatriz[59][56] = 9'b101001000;
assign micromatriz[59][57] = 9'b110010001;
assign micromatriz[59][58] = 9'b110110110;
assign micromatriz[59][59] = 9'b101001001;
assign micromatriz[59][60] = 9'b100000000;
assign micromatriz[59][61] = 9'b100000000;
assign micromatriz[59][62] = 9'b110111111;
assign micromatriz[59][63] = 9'b111111111;
assign micromatriz[59][64] = 9'b110110111;
assign micromatriz[59][65] = 9'b110110111;
assign micromatriz[59][66] = 9'b101101101;
assign micromatriz[59][67] = 9'b100000000;
assign micromatriz[59][68] = 9'b100000000;
assign micromatriz[59][69] = 9'b111111111;
assign micromatriz[59][70] = 9'b111111111;
assign micromatriz[59][71] = 9'b110110110;
assign micromatriz[59][72] = 9'b101101101;
assign micromatriz[59][73] = 9'b101101101;
assign micromatriz[59][74] = 9'b101101101;
assign micromatriz[59][75] = 9'b101101101;
assign micromatriz[59][76] = 9'b101001001;
assign micromatriz[59][77] = 9'b101001001;
assign micromatriz[59][78] = 9'b101001101;
assign micromatriz[59][79] = 9'b101101101;
assign micromatriz[59][80] = 9'b101101101;
assign micromatriz[59][81] = 9'b110010010;
assign micromatriz[59][82] = 9'b110111111;
assign micromatriz[59][83] = 9'b101001001;
assign micromatriz[59][84] = 9'b100000000;
assign micromatriz[59][85] = 9'b100100100;
assign micromatriz[59][86] = 9'b111111111;
assign micromatriz[59][87] = 9'b111111111;
assign micromatriz[59][88] = 9'b111111111;
assign micromatriz[59][89] = 9'b111111111;
assign micromatriz[59][90] = 9'b111111111;
assign micromatriz[59][91] = 9'b111111111;
assign micromatriz[59][92] = 9'b111111111;
assign micromatriz[59][93] = 9'b111111111;
assign micromatriz[59][94] = 9'b111111111;
assign micromatriz[59][95] = 9'b111111111;
assign micromatriz[59][96] = 9'b111111111;
assign micromatriz[59][97] = 9'b111111111;
assign micromatriz[59][98] = 9'b111111111;
assign micromatriz[59][99] = 9'b111111111;
assign micromatriz[60][0] = 9'b111111111;
assign micromatriz[60][1] = 9'b111111111;
assign micromatriz[60][2] = 9'b111111111;
assign micromatriz[60][3] = 9'b111111111;
assign micromatriz[60][4] = 9'b111111111;
assign micromatriz[60][5] = 9'b111111111;
assign micromatriz[60][6] = 9'b111111111;
assign micromatriz[60][7] = 9'b111111111;
assign micromatriz[60][8] = 9'b111111111;
assign micromatriz[60][9] = 9'b111111111;
assign micromatriz[60][10] = 9'b111111111;
assign micromatriz[60][11] = 9'b111111111;
assign micromatriz[60][12] = 9'b111111111;
assign micromatriz[60][13] = 9'b111111111;
assign micromatriz[60][14] = 9'b100100100;
assign micromatriz[60][15] = 9'b100000000;
assign micromatriz[60][16] = 9'b101101101;
assign micromatriz[60][17] = 9'b111111111;
assign micromatriz[60][18] = 9'b111111111;
assign micromatriz[60][19] = 9'b111111111;
assign micromatriz[60][20] = 9'b111111111;
assign micromatriz[60][21] = 9'b100101000;
assign micromatriz[60][22] = 9'b100000000;
assign micromatriz[60][23] = 9'b100100100;
assign micromatriz[60][24] = 9'b101101101;
assign micromatriz[60][25] = 9'b101101101;
assign micromatriz[60][26] = 9'b110010010;
assign micromatriz[60][27] = 9'b110110110;
assign micromatriz[60][28] = 9'b110110110;
assign micromatriz[60][29] = 9'b110110110;
assign micromatriz[60][30] = 9'b110110110;
assign micromatriz[60][31] = 9'b110110110;
assign micromatriz[60][32] = 9'b110110110;
assign micromatriz[60][33] = 9'b110110110;
assign micromatriz[60][34] = 9'b110110110;
assign micromatriz[60][35] = 9'b110110110;
assign micromatriz[60][36] = 9'b110110110;
assign micromatriz[60][37] = 9'b110110110;
assign micromatriz[60][38] = 9'b110110110;
assign micromatriz[60][39] = 9'b110110110;
assign micromatriz[60][40] = 9'b110110110;
assign micromatriz[60][41] = 9'b110110110;
assign micromatriz[60][42] = 9'b110110110;
assign micromatriz[60][43] = 9'b110110110;
assign micromatriz[60][44] = 9'b110110110;
assign micromatriz[60][45] = 9'b110110110;
assign micromatriz[60][46] = 9'b110110110;
assign micromatriz[60][47] = 9'b110110110;
assign micromatriz[60][48] = 9'b110110110;
assign micromatriz[60][49] = 9'b110110110;
assign micromatriz[60][50] = 9'b110110110;
assign micromatriz[60][51] = 9'b110110110;
assign micromatriz[60][52] = 9'b110110110;
assign micromatriz[60][53] = 9'b110110110;
assign micromatriz[60][54] = 9'b110110110;
assign micromatriz[60][55] = 9'b110110110;
assign micromatriz[60][56] = 9'b110110110;
assign micromatriz[60][57] = 9'b110010010;
assign micromatriz[60][58] = 9'b110110110;
assign micromatriz[60][59] = 9'b101001001;
assign micromatriz[60][60] = 9'b100000000;
assign micromatriz[60][61] = 9'b100000000;
assign micromatriz[60][62] = 9'b110111111;
assign micromatriz[60][63] = 9'b111111111;
assign micromatriz[60][64] = 9'b110110111;
assign micromatriz[60][65] = 9'b110110111;
assign micromatriz[60][66] = 9'b101101101;
assign micromatriz[60][67] = 9'b100000000;
assign micromatriz[60][68] = 9'b100000000;
assign micromatriz[60][69] = 9'b111111111;
assign micromatriz[60][70] = 9'b111111111;
assign micromatriz[60][71] = 9'b101101101;
assign micromatriz[60][72] = 9'b100000000;
assign micromatriz[60][73] = 9'b100000000;
assign micromatriz[60][74] = 9'b111111111;
assign micromatriz[60][75] = 9'b111111111;
assign micromatriz[60][76] = 9'b111111111;
assign micromatriz[60][77] = 9'b111111111;
assign micromatriz[60][78] = 9'b110010010;
assign micromatriz[60][79] = 9'b100000000;
assign micromatriz[60][80] = 9'b100000000;
assign micromatriz[60][81] = 9'b110010010;
assign micromatriz[60][82] = 9'b111111111;
assign micromatriz[60][83] = 9'b101001001;
assign micromatriz[60][84] = 9'b100000000;
assign micromatriz[60][85] = 9'b100100100;
assign micromatriz[60][86] = 9'b111111111;
assign micromatriz[60][87] = 9'b111111111;
assign micromatriz[60][88] = 9'b111111111;
assign micromatriz[60][89] = 9'b111111111;
assign micromatriz[60][90] = 9'b111111111;
assign micromatriz[60][91] = 9'b111111111;
assign micromatriz[60][92] = 9'b111111111;
assign micromatriz[60][93] = 9'b111111111;
assign micromatriz[60][94] = 9'b111111111;
assign micromatriz[60][95] = 9'b111111111;
assign micromatriz[60][96] = 9'b111111111;
assign micromatriz[60][97] = 9'b111111111;
assign micromatriz[60][98] = 9'b111111111;
assign micromatriz[60][99] = 9'b111111111;
assign micromatriz[61][0] = 9'b111111111;
assign micromatriz[61][1] = 9'b111111111;
assign micromatriz[61][2] = 9'b111111111;
assign micromatriz[61][3] = 9'b111111111;
assign micromatriz[61][4] = 9'b111111111;
assign micromatriz[61][5] = 9'b111111111;
assign micromatriz[61][6] = 9'b111111111;
assign micromatriz[61][7] = 9'b111111111;
assign micromatriz[61][8] = 9'b111111111;
assign micromatriz[61][9] = 9'b111111111;
assign micromatriz[61][10] = 9'b111111111;
assign micromatriz[61][11] = 9'b111111111;
assign micromatriz[61][12] = 9'b111111111;
assign micromatriz[61][13] = 9'b111111111;
assign micromatriz[61][14] = 9'b100100100;
assign micromatriz[61][15] = 9'b100000000;
assign micromatriz[61][16] = 9'b101101101;
assign micromatriz[61][17] = 9'b111111111;
assign micromatriz[61][18] = 9'b111111111;
assign micromatriz[61][19] = 9'b111111111;
assign micromatriz[61][20] = 9'b111111111;
assign micromatriz[61][21] = 9'b100101000;
assign micromatriz[61][22] = 9'b100000000;
assign micromatriz[61][23] = 9'b100100100;
assign micromatriz[61][24] = 9'b101101101;
assign micromatriz[61][25] = 9'b101101101;
assign micromatriz[61][26] = 9'b110010001;
assign micromatriz[61][27] = 9'b110010001;
assign micromatriz[61][28] = 9'b110010001;
assign micromatriz[61][29] = 9'b110010001;
assign micromatriz[61][30] = 9'b110010001;
assign micromatriz[61][31] = 9'b110010001;
assign micromatriz[61][32] = 9'b110010001;
assign micromatriz[61][33] = 9'b110010001;
assign micromatriz[61][34] = 9'b110010001;
assign micromatriz[61][35] = 9'b110010001;
assign micromatriz[61][36] = 9'b110010001;
assign micromatriz[61][37] = 9'b110010001;
assign micromatriz[61][38] = 9'b110010001;
assign micromatriz[61][39] = 9'b110010001;
assign micromatriz[61][40] = 9'b110010001;
assign micromatriz[61][41] = 9'b110010001;
assign micromatriz[61][42] = 9'b110010001;
assign micromatriz[61][43] = 9'b110010001;
assign micromatriz[61][44] = 9'b110010001;
assign micromatriz[61][45] = 9'b110010001;
assign micromatriz[61][46] = 9'b110010001;
assign micromatriz[61][47] = 9'b110010001;
assign micromatriz[61][48] = 9'b110010001;
assign micromatriz[61][49] = 9'b110010001;
assign micromatriz[61][50] = 9'b110010001;
assign micromatriz[61][51] = 9'b110010001;
assign micromatriz[61][52] = 9'b110010001;
assign micromatriz[61][53] = 9'b110010001;
assign micromatriz[61][54] = 9'b110010001;
assign micromatriz[61][55] = 9'b110010001;
assign micromatriz[61][56] = 9'b110010001;
assign micromatriz[61][57] = 9'b110010001;
assign micromatriz[61][58] = 9'b110010001;
assign micromatriz[61][59] = 9'b101001001;
assign micromatriz[61][60] = 9'b100000000;
assign micromatriz[61][61] = 9'b100000000;
assign micromatriz[61][62] = 9'b110111111;
assign micromatriz[61][63] = 9'b111111111;
assign micromatriz[61][64] = 9'b110110111;
assign micromatriz[61][65] = 9'b110110111;
assign micromatriz[61][66] = 9'b101101101;
assign micromatriz[61][67] = 9'b100000000;
assign micromatriz[61][68] = 9'b100000000;
assign micromatriz[61][69] = 9'b111111111;
assign micromatriz[61][70] = 9'b111111111;
assign micromatriz[61][71] = 9'b101101101;
assign micromatriz[61][72] = 9'b100000000;
assign micromatriz[61][73] = 9'b100000100;
assign micromatriz[61][74] = 9'b111111111;
assign micromatriz[61][75] = 9'b111111111;
assign micromatriz[61][76] = 9'b111111111;
assign micromatriz[61][77] = 9'b111111111;
assign micromatriz[61][78] = 9'b110010001;
assign micromatriz[61][79] = 9'b100000000;
assign micromatriz[61][80] = 9'b100000000;
assign micromatriz[61][81] = 9'b110010010;
assign micromatriz[61][82] = 9'b111111111;
assign micromatriz[61][83] = 9'b101001001;
assign micromatriz[61][84] = 9'b100000000;
assign micromatriz[61][85] = 9'b100100100;
assign micromatriz[61][86] = 9'b111111111;
assign micromatriz[61][87] = 9'b111111111;
assign micromatriz[61][88] = 9'b111111111;
assign micromatriz[61][89] = 9'b111111111;
assign micromatriz[61][90] = 9'b111111111;
assign micromatriz[61][91] = 9'b111111111;
assign micromatriz[61][92] = 9'b111111111;
assign micromatriz[61][93] = 9'b111111111;
assign micromatriz[61][94] = 9'b111111111;
assign micromatriz[61][95] = 9'b111111111;
assign micromatriz[61][96] = 9'b111111111;
assign micromatriz[61][97] = 9'b111111111;
assign micromatriz[61][98] = 9'b111111111;
assign micromatriz[61][99] = 9'b111111111;
assign micromatriz[62][0] = 9'b111111111;
assign micromatriz[62][1] = 9'b111111111;
assign micromatriz[62][2] = 9'b111111111;
assign micromatriz[62][3] = 9'b111111111;
assign micromatriz[62][4] = 9'b111111111;
assign micromatriz[62][5] = 9'b111111111;
assign micromatriz[62][6] = 9'b111111111;
assign micromatriz[62][7] = 9'b111111111;
assign micromatriz[62][8] = 9'b111111111;
assign micromatriz[62][9] = 9'b111111111;
assign micromatriz[62][10] = 9'b111111111;
assign micromatriz[62][11] = 9'b111111111;
assign micromatriz[62][12] = 9'b111111111;
assign micromatriz[62][13] = 9'b111111111;
assign micromatriz[62][14] = 9'b100100100;
assign micromatriz[62][15] = 9'b100000000;
assign micromatriz[62][16] = 9'b101101101;
assign micromatriz[62][17] = 9'b111111111;
assign micromatriz[62][18] = 9'b111111111;
assign micromatriz[62][19] = 9'b111111111;
assign micromatriz[62][20] = 9'b111111111;
assign micromatriz[62][21] = 9'b100101000;
assign micromatriz[62][22] = 9'b100000000;
assign micromatriz[62][23] = 9'b100000000;
assign micromatriz[62][24] = 9'b100000000;
assign micromatriz[62][25] = 9'b100000000;
assign micromatriz[62][26] = 9'b100000000;
assign micromatriz[62][27] = 9'b100000000;
assign micromatriz[62][28] = 9'b100000000;
assign micromatriz[62][29] = 9'b100000000;
assign micromatriz[62][30] = 9'b100000000;
assign micromatriz[62][31] = 9'b100000000;
assign micromatriz[62][32] = 9'b100000000;
assign micromatriz[62][33] = 9'b100000000;
assign micromatriz[62][34] = 9'b100000000;
assign micromatriz[62][35] = 9'b100000000;
assign micromatriz[62][36] = 9'b100000000;
assign micromatriz[62][37] = 9'b100000000;
assign micromatriz[62][38] = 9'b100000000;
assign micromatriz[62][39] = 9'b100000000;
assign micromatriz[62][40] = 9'b100000000;
assign micromatriz[62][41] = 9'b100000000;
assign micromatriz[62][42] = 9'b100000000;
assign micromatriz[62][43] = 9'b100000000;
assign micromatriz[62][44] = 9'b100000000;
assign micromatriz[62][45] = 9'b100000000;
assign micromatriz[62][46] = 9'b100000000;
assign micromatriz[62][47] = 9'b100000000;
assign micromatriz[62][48] = 9'b100000000;
assign micromatriz[62][49] = 9'b100000000;
assign micromatriz[62][50] = 9'b100000000;
assign micromatriz[62][51] = 9'b100000000;
assign micromatriz[62][52] = 9'b100000000;
assign micromatriz[62][53] = 9'b100000000;
assign micromatriz[62][54] = 9'b100000000;
assign micromatriz[62][55] = 9'b100000000;
assign micromatriz[62][56] = 9'b100000000;
assign micromatriz[62][57] = 9'b100000000;
assign micromatriz[62][58] = 9'b100000000;
assign micromatriz[62][59] = 9'b100000000;
assign micromatriz[62][60] = 9'b100000000;
assign micromatriz[62][61] = 9'b100000000;
assign micromatriz[62][62] = 9'b110111111;
assign micromatriz[62][63] = 9'b111111111;
assign micromatriz[62][64] = 9'b110110111;
assign micromatriz[62][65] = 9'b110110111;
assign micromatriz[62][66] = 9'b101101101;
assign micromatriz[62][67] = 9'b100000000;
assign micromatriz[62][68] = 9'b100000000;
assign micromatriz[62][69] = 9'b111111111;
assign micromatriz[62][70] = 9'b111111111;
assign micromatriz[62][71] = 9'b101101101;
assign micromatriz[62][72] = 9'b100000000;
assign micromatriz[62][73] = 9'b100000000;
assign micromatriz[62][74] = 9'b111111111;
assign micromatriz[62][75] = 9'b111111111;
assign micromatriz[62][76] = 9'b110110111;
assign micromatriz[62][77] = 9'b110110111;
assign micromatriz[62][78] = 9'b101101101;
assign micromatriz[62][79] = 9'b100000000;
assign micromatriz[62][80] = 9'b100000000;
assign micromatriz[62][81] = 9'b110010010;
assign micromatriz[62][82] = 9'b111111111;
assign micromatriz[62][83] = 9'b101001001;
assign micromatriz[62][84] = 9'b100000000;
assign micromatriz[62][85] = 9'b100100100;
assign micromatriz[62][86] = 9'b111111111;
assign micromatriz[62][87] = 9'b111111111;
assign micromatriz[62][88] = 9'b111111111;
assign micromatriz[62][89] = 9'b111111111;
assign micromatriz[62][90] = 9'b111111111;
assign micromatriz[62][91] = 9'b111111111;
assign micromatriz[62][92] = 9'b111111111;
assign micromatriz[62][93] = 9'b111111111;
assign micromatriz[62][94] = 9'b111111111;
assign micromatriz[62][95] = 9'b111111111;
assign micromatriz[62][96] = 9'b111111111;
assign micromatriz[62][97] = 9'b111111111;
assign micromatriz[62][98] = 9'b111111111;
assign micromatriz[62][99] = 9'b111111111;
assign micromatriz[63][0] = 9'b111111111;
assign micromatriz[63][1] = 9'b111111111;
assign micromatriz[63][2] = 9'b111111111;
assign micromatriz[63][3] = 9'b111111111;
assign micromatriz[63][4] = 9'b111111111;
assign micromatriz[63][5] = 9'b111111111;
assign micromatriz[63][6] = 9'b111111111;
assign micromatriz[63][7] = 9'b111111111;
assign micromatriz[63][8] = 9'b111111111;
assign micromatriz[63][9] = 9'b111111111;
assign micromatriz[63][10] = 9'b111111111;
assign micromatriz[63][11] = 9'b111111111;
assign micromatriz[63][12] = 9'b111111111;
assign micromatriz[63][13] = 9'b111111111;
assign micromatriz[63][14] = 9'b100100100;
assign micromatriz[63][15] = 9'b100000000;
assign micromatriz[63][16] = 9'b101101101;
assign micromatriz[63][17] = 9'b111111111;
assign micromatriz[63][18] = 9'b111111111;
assign micromatriz[63][19] = 9'b111111111;
assign micromatriz[63][20] = 9'b111111111;
assign micromatriz[63][21] = 9'b100100100;
assign micromatriz[63][22] = 9'b100000000;
assign micromatriz[63][23] = 9'b100000000;
assign micromatriz[63][24] = 9'b100000000;
assign micromatriz[63][25] = 9'b100000000;
assign micromatriz[63][26] = 9'b100000000;
assign micromatriz[63][27] = 9'b100000000;
assign micromatriz[63][28] = 9'b100000000;
assign micromatriz[63][29] = 9'b100000000;
assign micromatriz[63][30] = 9'b100000000;
assign micromatriz[63][31] = 9'b100000000;
assign micromatriz[63][32] = 9'b100000000;
assign micromatriz[63][33] = 9'b100000000;
assign micromatriz[63][34] = 9'b100000000;
assign micromatriz[63][35] = 9'b100000000;
assign micromatriz[63][36] = 9'b100000000;
assign micromatriz[63][37] = 9'b100000000;
assign micromatriz[63][38] = 9'b100000000;
assign micromatriz[63][39] = 9'b100000000;
assign micromatriz[63][40] = 9'b100000000;
assign micromatriz[63][41] = 9'b100000000;
assign micromatriz[63][42] = 9'b100000000;
assign micromatriz[63][43] = 9'b100000000;
assign micromatriz[63][44] = 9'b100000000;
assign micromatriz[63][45] = 9'b100000000;
assign micromatriz[63][46] = 9'b100000000;
assign micromatriz[63][47] = 9'b100000000;
assign micromatriz[63][48] = 9'b100000000;
assign micromatriz[63][49] = 9'b100000000;
assign micromatriz[63][50] = 9'b100000000;
assign micromatriz[63][51] = 9'b100000000;
assign micromatriz[63][52] = 9'b100000000;
assign micromatriz[63][53] = 9'b100000000;
assign micromatriz[63][54] = 9'b100000000;
assign micromatriz[63][55] = 9'b100000000;
assign micromatriz[63][56] = 9'b100000000;
assign micromatriz[63][57] = 9'b100000000;
assign micromatriz[63][58] = 9'b100000000;
assign micromatriz[63][59] = 9'b100000000;
assign micromatriz[63][60] = 9'b100000000;
assign micromatriz[63][61] = 9'b100000000;
assign micromatriz[63][62] = 9'b110111111;
assign micromatriz[63][63] = 9'b111111111;
assign micromatriz[63][64] = 9'b110110111;
assign micromatriz[63][65] = 9'b110110111;
assign micromatriz[63][66] = 9'b101101101;
assign micromatriz[63][67] = 9'b100000000;
assign micromatriz[63][68] = 9'b100000000;
assign micromatriz[63][69] = 9'b111111111;
assign micromatriz[63][70] = 9'b111111111;
assign micromatriz[63][71] = 9'b101101101;
assign micromatriz[63][72] = 9'b100000000;
assign micromatriz[63][73] = 9'b100000000;
assign micromatriz[63][74] = 9'b111111111;
assign micromatriz[63][75] = 9'b111111111;
assign micromatriz[63][76] = 9'b111111111;
assign micromatriz[63][77] = 9'b111111111;
assign micromatriz[63][78] = 9'b101101101;
assign micromatriz[63][79] = 9'b100000000;
assign micromatriz[63][80] = 9'b100000000;
assign micromatriz[63][81] = 9'b110010010;
assign micromatriz[63][82] = 9'b111111111;
assign micromatriz[63][83] = 9'b101001001;
assign micromatriz[63][84] = 9'b100000000;
assign micromatriz[63][85] = 9'b100100100;
assign micromatriz[63][86] = 9'b111111111;
assign micromatriz[63][87] = 9'b111111111;
assign micromatriz[63][88] = 9'b111111111;
assign micromatriz[63][89] = 9'b111111111;
assign micromatriz[63][90] = 9'b111111111;
assign micromatriz[63][91] = 9'b111111111;
assign micromatriz[63][92] = 9'b111111111;
assign micromatriz[63][93] = 9'b111111111;
assign micromatriz[63][94] = 9'b111111111;
assign micromatriz[63][95] = 9'b111111111;
assign micromatriz[63][96] = 9'b111111111;
assign micromatriz[63][97] = 9'b111111111;
assign micromatriz[63][98] = 9'b111111111;
assign micromatriz[63][99] = 9'b111111111;
assign micromatriz[64][0] = 9'b111111111;
assign micromatriz[64][1] = 9'b111111111;
assign micromatriz[64][2] = 9'b111111111;
assign micromatriz[64][3] = 9'b111111111;
assign micromatriz[64][4] = 9'b111111111;
assign micromatriz[64][5] = 9'b111111111;
assign micromatriz[64][6] = 9'b111111111;
assign micromatriz[64][7] = 9'b111111111;
assign micromatriz[64][8] = 9'b111111111;
assign micromatriz[64][9] = 9'b111111111;
assign micromatriz[64][10] = 9'b111111111;
assign micromatriz[64][11] = 9'b111111111;
assign micromatriz[64][12] = 9'b111111111;
assign micromatriz[64][13] = 9'b111111111;
assign micromatriz[64][14] = 9'b100100100;
assign micromatriz[64][15] = 9'b100000000;
assign micromatriz[64][16] = 9'b101101101;
assign micromatriz[64][17] = 9'b111111111;
assign micromatriz[64][18] = 9'b111111111;
assign micromatriz[64][19] = 9'b111111111;
assign micromatriz[64][20] = 9'b111111111;
assign micromatriz[64][21] = 9'b110010010;
assign micromatriz[64][22] = 9'b101101101;
assign micromatriz[64][23] = 9'b101110001;
assign micromatriz[64][24] = 9'b101110001;
assign micromatriz[64][25] = 9'b101110001;
assign micromatriz[64][26] = 9'b101110001;
assign micromatriz[64][27] = 9'b101110001;
assign micromatriz[64][28] = 9'b101110001;
assign micromatriz[64][29] = 9'b101110001;
assign micromatriz[64][30] = 9'b101110001;
assign micromatriz[64][31] = 9'b101110001;
assign micromatriz[64][32] = 9'b101110001;
assign micromatriz[64][33] = 9'b101110001;
assign micromatriz[64][34] = 9'b101110001;
assign micromatriz[64][35] = 9'b101110001;
assign micromatriz[64][36] = 9'b101110001;
assign micromatriz[64][37] = 9'b101110001;
assign micromatriz[64][38] = 9'b101110001;
assign micromatriz[64][39] = 9'b101110001;
assign micromatriz[64][40] = 9'b101110001;
assign micromatriz[64][41] = 9'b101110001;
assign micromatriz[64][42] = 9'b101110001;
assign micromatriz[64][43] = 9'b101110001;
assign micromatriz[64][44] = 9'b101110001;
assign micromatriz[64][45] = 9'b101110001;
assign micromatriz[64][46] = 9'b101110001;
assign micromatriz[64][47] = 9'b101110001;
assign micromatriz[64][48] = 9'b101110001;
assign micromatriz[64][49] = 9'b101110001;
assign micromatriz[64][50] = 9'b101110001;
assign micromatriz[64][51] = 9'b101110001;
assign micromatriz[64][52] = 9'b101110001;
assign micromatriz[64][53] = 9'b101110001;
assign micromatriz[64][54] = 9'b101110001;
assign micromatriz[64][55] = 9'b101110001;
assign micromatriz[64][56] = 9'b101110001;
assign micromatriz[64][57] = 9'b101110001;
assign micromatriz[64][58] = 9'b101110001;
assign micromatriz[64][59] = 9'b101110001;
assign micromatriz[64][60] = 9'b101110001;
assign micromatriz[64][61] = 9'b101110001;
assign micromatriz[64][62] = 9'b111111111;
assign micromatriz[64][63] = 9'b111111111;
assign micromatriz[64][64] = 9'b110110111;
assign micromatriz[64][65] = 9'b110110111;
assign micromatriz[64][66] = 9'b101101101;
assign micromatriz[64][67] = 9'b100000000;
assign micromatriz[64][68] = 9'b100000000;
assign micromatriz[64][69] = 9'b111111111;
assign micromatriz[64][70] = 9'b111111111;
assign micromatriz[64][71] = 9'b110110111;
assign micromatriz[64][72] = 9'b101110001;
assign micromatriz[64][73] = 9'b101101101;
assign micromatriz[64][74] = 9'b101001001;
assign micromatriz[64][75] = 9'b101001001;
assign micromatriz[64][76] = 9'b100101000;
assign micromatriz[64][77] = 9'b100100100;
assign micromatriz[64][78] = 9'b101001001;
assign micromatriz[64][79] = 9'b110010001;
assign micromatriz[64][80] = 9'b101110001;
assign micromatriz[64][81] = 9'b110010110;
assign micromatriz[64][82] = 9'b110111111;
assign micromatriz[64][83] = 9'b101001001;
assign micromatriz[64][84] = 9'b100000000;
assign micromatriz[64][85] = 9'b100100100;
assign micromatriz[64][86] = 9'b111111111;
assign micromatriz[64][87] = 9'b111111111;
assign micromatriz[64][88] = 9'b111111111;
assign micromatriz[64][89] = 9'b111111111;
assign micromatriz[64][90] = 9'b111111111;
assign micromatriz[64][91] = 9'b111111111;
assign micromatriz[64][92] = 9'b111111111;
assign micromatriz[64][93] = 9'b111111111;
assign micromatriz[64][94] = 9'b111111111;
assign micromatriz[64][95] = 9'b111111111;
assign micromatriz[64][96] = 9'b111111111;
assign micromatriz[64][97] = 9'b111111111;
assign micromatriz[64][98] = 9'b111111111;
assign micromatriz[64][99] = 9'b111111111;
assign micromatriz[65][0] = 9'b111111111;
assign micromatriz[65][1] = 9'b111111111;
assign micromatriz[65][2] = 9'b111111111;
assign micromatriz[65][3] = 9'b111111111;
assign micromatriz[65][4] = 9'b111111111;
assign micromatriz[65][5] = 9'b111111111;
assign micromatriz[65][6] = 9'b111111111;
assign micromatriz[65][7] = 9'b111111111;
assign micromatriz[65][8] = 9'b111111111;
assign micromatriz[65][9] = 9'b111111111;
assign micromatriz[65][10] = 9'b111111111;
assign micromatriz[65][11] = 9'b111111111;
assign micromatriz[65][12] = 9'b111111111;
assign micromatriz[65][13] = 9'b111111111;
assign micromatriz[65][14] = 9'b100100100;
assign micromatriz[65][15] = 9'b100000000;
assign micromatriz[65][16] = 9'b101101101;
assign micromatriz[65][17] = 9'b111111111;
assign micromatriz[65][18] = 9'b111111111;
assign micromatriz[65][19] = 9'b111111111;
assign micromatriz[65][20] = 9'b111111111;
assign micromatriz[65][21] = 9'b111111111;
assign micromatriz[65][22] = 9'b111111111;
assign micromatriz[65][23] = 9'b111111111;
assign micromatriz[65][24] = 9'b111111111;
assign micromatriz[65][25] = 9'b111111111;
assign micromatriz[65][26] = 9'b111111111;
assign micromatriz[65][27] = 9'b111111111;
assign micromatriz[65][28] = 9'b111111111;
assign micromatriz[65][29] = 9'b111111111;
assign micromatriz[65][30] = 9'b111111111;
assign micromatriz[65][31] = 9'b111111111;
assign micromatriz[65][32] = 9'b111111111;
assign micromatriz[65][33] = 9'b111111111;
assign micromatriz[65][34] = 9'b111111111;
assign micromatriz[65][35] = 9'b111111111;
assign micromatriz[65][36] = 9'b111111111;
assign micromatriz[65][37] = 9'b111111111;
assign micromatriz[65][38] = 9'b111111111;
assign micromatriz[65][39] = 9'b111111111;
assign micromatriz[65][40] = 9'b111111111;
assign micromatriz[65][41] = 9'b111111111;
assign micromatriz[65][42] = 9'b111111111;
assign micromatriz[65][43] = 9'b111111111;
assign micromatriz[65][44] = 9'b111111111;
assign micromatriz[65][45] = 9'b111111111;
assign micromatriz[65][46] = 9'b111111111;
assign micromatriz[65][47] = 9'b111111111;
assign micromatriz[65][48] = 9'b111111111;
assign micromatriz[65][49] = 9'b111111111;
assign micromatriz[65][50] = 9'b111111111;
assign micromatriz[65][51] = 9'b111111111;
assign micromatriz[65][52] = 9'b111111111;
assign micromatriz[65][53] = 9'b111111111;
assign micromatriz[65][54] = 9'b111111111;
assign micromatriz[65][55] = 9'b111111111;
assign micromatriz[65][56] = 9'b111111111;
assign micromatriz[65][57] = 9'b111111111;
assign micromatriz[65][58] = 9'b111111111;
assign micromatriz[65][59] = 9'b111111111;
assign micromatriz[65][60] = 9'b111111111;
assign micromatriz[65][61] = 9'b111111111;
assign micromatriz[65][62] = 9'b111111111;
assign micromatriz[65][63] = 9'b111111111;
assign micromatriz[65][64] = 9'b110110111;
assign micromatriz[65][65] = 9'b110110111;
assign micromatriz[65][66] = 9'b101101101;
assign micromatriz[65][67] = 9'b100000000;
assign micromatriz[65][68] = 9'b100000000;
assign micromatriz[65][69] = 9'b111111111;
assign micromatriz[65][70] = 9'b111111111;
assign micromatriz[65][71] = 9'b111111111;
assign micromatriz[65][72] = 9'b111111111;
assign micromatriz[65][73] = 9'b110111111;
assign micromatriz[65][74] = 9'b100000000;
assign micromatriz[65][75] = 9'b100000000;
assign micromatriz[65][76] = 9'b100000000;
assign micromatriz[65][77] = 9'b100000000;
assign micromatriz[65][78] = 9'b100100100;
assign micromatriz[65][79] = 9'b111111111;
assign micromatriz[65][80] = 9'b111111111;
assign micromatriz[65][81] = 9'b110110111;
assign micromatriz[65][82] = 9'b110111111;
assign micromatriz[65][83] = 9'b101001001;
assign micromatriz[65][84] = 9'b100000000;
assign micromatriz[65][85] = 9'b100100100;
assign micromatriz[65][86] = 9'b111111111;
assign micromatriz[65][87] = 9'b111111111;
assign micromatriz[65][88] = 9'b111111111;
assign micromatriz[65][89] = 9'b111111111;
assign micromatriz[65][90] = 9'b111111111;
assign micromatriz[65][91] = 9'b111111111;
assign micromatriz[65][92] = 9'b111111111;
assign micromatriz[65][93] = 9'b111111111;
assign micromatriz[65][94] = 9'b111111111;
assign micromatriz[65][95] = 9'b111111111;
assign micromatriz[65][96] = 9'b111111111;
assign micromatriz[65][97] = 9'b111111111;
assign micromatriz[65][98] = 9'b111111111;
assign micromatriz[65][99] = 9'b111111111;
assign micromatriz[66][0] = 9'b111111111;
assign micromatriz[66][1] = 9'b111111111;
assign micromatriz[66][2] = 9'b111111111;
assign micromatriz[66][3] = 9'b111111111;
assign micromatriz[66][4] = 9'b111111111;
assign micromatriz[66][5] = 9'b111111111;
assign micromatriz[66][6] = 9'b111111111;
assign micromatriz[66][7] = 9'b111111111;
assign micromatriz[66][8] = 9'b111111111;
assign micromatriz[66][9] = 9'b111111111;
assign micromatriz[66][10] = 9'b111111111;
assign micromatriz[66][11] = 9'b111111111;
assign micromatriz[66][12] = 9'b111111111;
assign micromatriz[66][13] = 9'b111111111;
assign micromatriz[66][14] = 9'b100100100;
assign micromatriz[66][15] = 9'b100000000;
assign micromatriz[66][16] = 9'b101101101;
assign micromatriz[66][17] = 9'b111111111;
assign micromatriz[66][18] = 9'b111111111;
assign micromatriz[66][19] = 9'b110111111;
assign micromatriz[66][20] = 9'b110111111;
assign micromatriz[66][21] = 9'b110111111;
assign micromatriz[66][22] = 9'b110111111;
assign micromatriz[66][23] = 9'b110111111;
assign micromatriz[66][24] = 9'b110111111;
assign micromatriz[66][25] = 9'b110111111;
assign micromatriz[66][26] = 9'b110111111;
assign micromatriz[66][27] = 9'b110111111;
assign micromatriz[66][28] = 9'b110111111;
assign micromatriz[66][29] = 9'b110111111;
assign micromatriz[66][30] = 9'b110111111;
assign micromatriz[66][31] = 9'b110111111;
assign micromatriz[66][32] = 9'b110111111;
assign micromatriz[66][33] = 9'b110111111;
assign micromatriz[66][34] = 9'b110111111;
assign micromatriz[66][35] = 9'b110111111;
assign micromatriz[66][36] = 9'b110111111;
assign micromatriz[66][37] = 9'b110111111;
assign micromatriz[66][38] = 9'b110111111;
assign micromatriz[66][39] = 9'b110111111;
assign micromatriz[66][40] = 9'b110111111;
assign micromatriz[66][41] = 9'b110111111;
assign micromatriz[66][42] = 9'b110111111;
assign micromatriz[66][43] = 9'b110111111;
assign micromatriz[66][44] = 9'b110111111;
assign micromatriz[66][45] = 9'b110111111;
assign micromatriz[66][46] = 9'b110111111;
assign micromatriz[66][47] = 9'b110111111;
assign micromatriz[66][48] = 9'b110111111;
assign micromatriz[66][49] = 9'b110111111;
assign micromatriz[66][50] = 9'b110111111;
assign micromatriz[66][51] = 9'b110111111;
assign micromatriz[66][52] = 9'b110111111;
assign micromatriz[66][53] = 9'b110111111;
assign micromatriz[66][54] = 9'b110111111;
assign micromatriz[66][55] = 9'b110111111;
assign micromatriz[66][56] = 9'b110111111;
assign micromatriz[66][57] = 9'b110111111;
assign micromatriz[66][58] = 9'b110111111;
assign micromatriz[66][59] = 9'b110111111;
assign micromatriz[66][60] = 9'b110111111;
assign micromatriz[66][61] = 9'b110111111;
assign micromatriz[66][62] = 9'b110111111;
assign micromatriz[66][63] = 9'b110111111;
assign micromatriz[66][64] = 9'b110110111;
assign micromatriz[66][65] = 9'b110110111;
assign micromatriz[66][66] = 9'b101101101;
assign micromatriz[66][67] = 9'b100000000;
assign micromatriz[66][68] = 9'b100000000;
assign micromatriz[66][69] = 9'b110111111;
assign micromatriz[66][70] = 9'b111111111;
assign micromatriz[66][71] = 9'b111111111;
assign micromatriz[66][72] = 9'b111111111;
assign micromatriz[66][73] = 9'b110110111;
assign micromatriz[66][74] = 9'b100100100;
assign micromatriz[66][75] = 9'b100100100;
assign micromatriz[66][76] = 9'b100100100;
assign micromatriz[66][77] = 9'b100100100;
assign micromatriz[66][78] = 9'b101001001;
assign micromatriz[66][79] = 9'b111111111;
assign micromatriz[66][80] = 9'b110111111;
assign micromatriz[66][81] = 9'b110110111;
assign micromatriz[66][82] = 9'b110111111;
assign micromatriz[66][83] = 9'b101001001;
assign micromatriz[66][84] = 9'b100000000;
assign micromatriz[66][85] = 9'b100100100;
assign micromatriz[66][86] = 9'b111111111;
assign micromatriz[66][87] = 9'b111111111;
assign micromatriz[66][88] = 9'b111111111;
assign micromatriz[66][89] = 9'b111111111;
assign micromatriz[66][90] = 9'b111111111;
assign micromatriz[66][91] = 9'b111111111;
assign micromatriz[66][92] = 9'b111111111;
assign micromatriz[66][93] = 9'b111111111;
assign micromatriz[66][94] = 9'b111111111;
assign micromatriz[66][95] = 9'b111111111;
assign micromatriz[66][96] = 9'b111111111;
assign micromatriz[66][97] = 9'b111111111;
assign micromatriz[66][98] = 9'b111111111;
assign micromatriz[66][99] = 9'b111111111;
assign micromatriz[67][0] = 9'b111111111;
assign micromatriz[67][1] = 9'b111111111;
assign micromatriz[67][2] = 9'b111111111;
assign micromatriz[67][3] = 9'b111111111;
assign micromatriz[67][4] = 9'b111111111;
assign micromatriz[67][5] = 9'b111111111;
assign micromatriz[67][6] = 9'b111111111;
assign micromatriz[67][7] = 9'b111111111;
assign micromatriz[67][8] = 9'b111111111;
assign micromatriz[67][9] = 9'b111111111;
assign micromatriz[67][10] = 9'b111111111;
assign micromatriz[67][11] = 9'b111111111;
assign micromatriz[67][12] = 9'b111111111;
assign micromatriz[67][13] = 9'b111111111;
assign micromatriz[67][14] = 9'b100100100;
assign micromatriz[67][15] = 9'b100000000;
assign micromatriz[67][16] = 9'b101001101;
assign micromatriz[67][17] = 9'b111111111;
assign micromatriz[67][18] = 9'b110111111;
assign micromatriz[67][19] = 9'b110110111;
assign micromatriz[67][20] = 9'b110110111;
assign micromatriz[67][21] = 9'b110110111;
assign micromatriz[67][22] = 9'b110110111;
assign micromatriz[67][23] = 9'b110110111;
assign micromatriz[67][24] = 9'b110110111;
assign micromatriz[67][25] = 9'b110110111;
assign micromatriz[67][26] = 9'b110110111;
assign micromatriz[67][27] = 9'b110110111;
assign micromatriz[67][28] = 9'b110110111;
assign micromatriz[67][29] = 9'b110110111;
assign micromatriz[67][30] = 9'b110110111;
assign micromatriz[67][31] = 9'b110110111;
assign micromatriz[67][32] = 9'b110110111;
assign micromatriz[67][33] = 9'b110110111;
assign micromatriz[67][34] = 9'b110110111;
assign micromatriz[67][35] = 9'b110110111;
assign micromatriz[67][36] = 9'b110110111;
assign micromatriz[67][37] = 9'b110110111;
assign micromatriz[67][38] = 9'b110110111;
assign micromatriz[67][39] = 9'b110110111;
assign micromatriz[67][40] = 9'b110110111;
assign micromatriz[67][41] = 9'b110110111;
assign micromatriz[67][42] = 9'b110110111;
assign micromatriz[67][43] = 9'b110110111;
assign micromatriz[67][44] = 9'b110110111;
assign micromatriz[67][45] = 9'b110110111;
assign micromatriz[67][46] = 9'b110110111;
assign micromatriz[67][47] = 9'b110110111;
assign micromatriz[67][48] = 9'b110110111;
assign micromatriz[67][49] = 9'b110110111;
assign micromatriz[67][50] = 9'b110110111;
assign micromatriz[67][51] = 9'b110110111;
assign micromatriz[67][52] = 9'b110110111;
assign micromatriz[67][53] = 9'b110110111;
assign micromatriz[67][54] = 9'b110110111;
assign micromatriz[67][55] = 9'b110110111;
assign micromatriz[67][56] = 9'b110110111;
assign micromatriz[67][57] = 9'b110110111;
assign micromatriz[67][58] = 9'b110110111;
assign micromatriz[67][59] = 9'b110110111;
assign micromatriz[67][60] = 9'b110110111;
assign micromatriz[67][61] = 9'b110110111;
assign micromatriz[67][62] = 9'b110110111;
assign micromatriz[67][63] = 9'b110110111;
assign micromatriz[67][64] = 9'b110110111;
assign micromatriz[67][65] = 9'b110111111;
assign micromatriz[67][66] = 9'b101101101;
assign micromatriz[67][67] = 9'b100000000;
assign micromatriz[67][68] = 9'b100000000;
assign micromatriz[67][69] = 9'b110010110;
assign micromatriz[67][70] = 9'b111111111;
assign micromatriz[67][71] = 9'b110111111;
assign micromatriz[67][72] = 9'b110010110;
assign micromatriz[67][73] = 9'b110110111;
assign micromatriz[67][74] = 9'b110111111;
assign micromatriz[67][75] = 9'b110111111;
assign micromatriz[67][76] = 9'b110111111;
assign micromatriz[67][77] = 9'b110111111;
assign micromatriz[67][78] = 9'b110110111;
assign micromatriz[67][79] = 9'b110010111;
assign micromatriz[67][80] = 9'b110110111;
assign micromatriz[67][81] = 9'b110110111;
assign micromatriz[67][82] = 9'b110111111;
assign micromatriz[67][83] = 9'b101001001;
assign micromatriz[67][84] = 9'b100000000;
assign micromatriz[67][85] = 9'b100100100;
assign micromatriz[67][86] = 9'b111111111;
assign micromatriz[67][87] = 9'b111111111;
assign micromatriz[67][88] = 9'b111111111;
assign micromatriz[67][89] = 9'b111111111;
assign micromatriz[67][90] = 9'b111111111;
assign micromatriz[67][91] = 9'b111111111;
assign micromatriz[67][92] = 9'b111111111;
assign micromatriz[67][93] = 9'b111111111;
assign micromatriz[67][94] = 9'b111111111;
assign micromatriz[67][95] = 9'b111111111;
assign micromatriz[67][96] = 9'b111111111;
assign micromatriz[67][97] = 9'b111111111;
assign micromatriz[67][98] = 9'b111111111;
assign micromatriz[67][99] = 9'b111111111;
assign micromatriz[68][0] = 9'b111111111;
assign micromatriz[68][1] = 9'b111111111;
assign micromatriz[68][2] = 9'b111111111;
assign micromatriz[68][3] = 9'b111111111;
assign micromatriz[68][4] = 9'b111111111;
assign micromatriz[68][5] = 9'b111111111;
assign micromatriz[68][6] = 9'b111111111;
assign micromatriz[68][7] = 9'b111111111;
assign micromatriz[68][8] = 9'b111111111;
assign micromatriz[68][9] = 9'b111111111;
assign micromatriz[68][10] = 9'b111111111;
assign micromatriz[68][11] = 9'b111111111;
assign micromatriz[68][12] = 9'b111111111;
assign micromatriz[68][13] = 9'b111111111;
assign micromatriz[68][14] = 9'b100100100;
assign micromatriz[68][15] = 9'b100000000;
assign micromatriz[68][16] = 9'b101101101;
assign micromatriz[68][17] = 9'b111111111;
assign micromatriz[68][18] = 9'b110111111;
assign micromatriz[68][19] = 9'b110110111;
assign micromatriz[68][20] = 9'b110110111;
assign micromatriz[68][21] = 9'b110110111;
assign micromatriz[68][22] = 9'b110110111;
assign micromatriz[68][23] = 9'b110110111;
assign micromatriz[68][24] = 9'b110110111;
assign micromatriz[68][25] = 9'b110110111;
assign micromatriz[68][26] = 9'b110110111;
assign micromatriz[68][27] = 9'b110110111;
assign micromatriz[68][28] = 9'b110110111;
assign micromatriz[68][29] = 9'b110110111;
assign micromatriz[68][30] = 9'b110110111;
assign micromatriz[68][31] = 9'b110110111;
assign micromatriz[68][32] = 9'b110110111;
assign micromatriz[68][33] = 9'b110110111;
assign micromatriz[68][34] = 9'b110110111;
assign micromatriz[68][35] = 9'b110110111;
assign micromatriz[68][36] = 9'b110110111;
assign micromatriz[68][37] = 9'b110110111;
assign micromatriz[68][38] = 9'b110110111;
assign micromatriz[68][39] = 9'b110110111;
assign micromatriz[68][40] = 9'b110110111;
assign micromatriz[68][41] = 9'b110110111;
assign micromatriz[68][42] = 9'b110110111;
assign micromatriz[68][43] = 9'b110110111;
assign micromatriz[68][44] = 9'b110110111;
assign micromatriz[68][45] = 9'b110110111;
assign micromatriz[68][46] = 9'b110110111;
assign micromatriz[68][47] = 9'b110110111;
assign micromatriz[68][48] = 9'b110110111;
assign micromatriz[68][49] = 9'b110110111;
assign micromatriz[68][50] = 9'b110110111;
assign micromatriz[68][51] = 9'b110110111;
assign micromatriz[68][52] = 9'b110110111;
assign micromatriz[68][53] = 9'b110110111;
assign micromatriz[68][54] = 9'b110110111;
assign micromatriz[68][55] = 9'b110110111;
assign micromatriz[68][56] = 9'b110110111;
assign micromatriz[68][57] = 9'b110110111;
assign micromatriz[68][58] = 9'b110110111;
assign micromatriz[68][59] = 9'b110110111;
assign micromatriz[68][60] = 9'b110110111;
assign micromatriz[68][61] = 9'b110110111;
assign micromatriz[68][62] = 9'b110110111;
assign micromatriz[68][63] = 9'b110110111;
assign micromatriz[68][64] = 9'b110110111;
assign micromatriz[68][65] = 9'b110111111;
assign micromatriz[68][66] = 9'b101101101;
assign micromatriz[68][67] = 9'b100000000;
assign micromatriz[68][68] = 9'b100000000;
assign micromatriz[68][69] = 9'b110010110;
assign micromatriz[68][70] = 9'b111111111;
assign micromatriz[68][71] = 9'b110111111;
assign micromatriz[68][72] = 9'b110110111;
assign micromatriz[68][73] = 9'b110110111;
assign micromatriz[68][74] = 9'b110110111;
assign micromatriz[68][75] = 9'b110110111;
assign micromatriz[68][76] = 9'b110110111;
assign micromatriz[68][77] = 9'b110110111;
assign micromatriz[68][78] = 9'b110110111;
assign micromatriz[68][79] = 9'b110110111;
assign micromatriz[68][80] = 9'b110110111;
assign micromatriz[68][81] = 9'b110110111;
assign micromatriz[68][82] = 9'b110111111;
assign micromatriz[68][83] = 9'b101001001;
assign micromatriz[68][84] = 9'b100000000;
assign micromatriz[68][85] = 9'b100100100;
assign micromatriz[68][86] = 9'b111111111;
assign micromatriz[68][87] = 9'b111111111;
assign micromatriz[68][88] = 9'b111111111;
assign micromatriz[68][89] = 9'b111111111;
assign micromatriz[68][90] = 9'b111111111;
assign micromatriz[68][91] = 9'b111111111;
assign micromatriz[68][92] = 9'b111111111;
assign micromatriz[68][93] = 9'b111111111;
assign micromatriz[68][94] = 9'b111111111;
assign micromatriz[68][95] = 9'b111111111;
assign micromatriz[68][96] = 9'b111111111;
assign micromatriz[68][97] = 9'b111111111;
assign micromatriz[68][98] = 9'b111111111;
assign micromatriz[68][99] = 9'b111111111;
assign micromatriz[69][0] = 9'b111111111;
assign micromatriz[69][1] = 9'b111111111;
assign micromatriz[69][2] = 9'b111111111;
assign micromatriz[69][3] = 9'b111111111;
assign micromatriz[69][4] = 9'b111111111;
assign micromatriz[69][5] = 9'b111111111;
assign micromatriz[69][6] = 9'b111111111;
assign micromatriz[69][7] = 9'b111111111;
assign micromatriz[69][8] = 9'b111111111;
assign micromatriz[69][9] = 9'b111111111;
assign micromatriz[69][10] = 9'b111111111;
assign micromatriz[69][11] = 9'b111111111;
assign micromatriz[69][12] = 9'b111111111;
assign micromatriz[69][13] = 9'b111111111;
assign micromatriz[69][14] = 9'b111111111;
assign micromatriz[69][15] = 9'b111111111;
assign micromatriz[69][16] = 9'b101101101;
assign micromatriz[69][17] = 9'b100100100;
assign micromatriz[69][18] = 9'b100100100;
assign micromatriz[69][19] = 9'b100000000;
assign micromatriz[69][20] = 9'b100000000;
assign micromatriz[69][21] = 9'b100000000;
assign micromatriz[69][22] = 9'b100000000;
assign micromatriz[69][23] = 9'b100000000;
assign micromatriz[69][24] = 9'b100000000;
assign micromatriz[69][25] = 9'b100000000;
assign micromatriz[69][26] = 9'b100000000;
assign micromatriz[69][27] = 9'b100000000;
assign micromatriz[69][28] = 9'b100000000;
assign micromatriz[69][29] = 9'b100000000;
assign micromatriz[69][30] = 9'b100000000;
assign micromatriz[69][31] = 9'b100000000;
assign micromatriz[69][32] = 9'b100000000;
assign micromatriz[69][33] = 9'b100000000;
assign micromatriz[69][34] = 9'b100000000;
assign micromatriz[69][35] = 9'b100000000;
assign micromatriz[69][36] = 9'b100000000;
assign micromatriz[69][37] = 9'b100000000;
assign micromatriz[69][38] = 9'b100000000;
assign micromatriz[69][39] = 9'b100000000;
assign micromatriz[69][40] = 9'b100000000;
assign micromatriz[69][41] = 9'b100000000;
assign micromatriz[69][42] = 9'b100000000;
assign micromatriz[69][43] = 9'b100000000;
assign micromatriz[69][44] = 9'b100000000;
assign micromatriz[69][45] = 9'b100000000;
assign micromatriz[69][46] = 9'b100000000;
assign micromatriz[69][47] = 9'b100000000;
assign micromatriz[69][48] = 9'b100000000;
assign micromatriz[69][49] = 9'b100000000;
assign micromatriz[69][50] = 9'b100000000;
assign micromatriz[69][51] = 9'b100000000;
assign micromatriz[69][52] = 9'b100000000;
assign micromatriz[69][53] = 9'b100000000;
assign micromatriz[69][54] = 9'b100000000;
assign micromatriz[69][55] = 9'b100000000;
assign micromatriz[69][56] = 9'b100000000;
assign micromatriz[69][57] = 9'b100000000;
assign micromatriz[69][58] = 9'b100000000;
assign micromatriz[69][59] = 9'b100000000;
assign micromatriz[69][60] = 9'b100000000;
assign micromatriz[69][61] = 9'b100000000;
assign micromatriz[69][62] = 9'b100000000;
assign micromatriz[69][63] = 9'b100000000;
assign micromatriz[69][64] = 9'b100000000;
assign micromatriz[69][65] = 9'b100100100;
assign micromatriz[69][66] = 9'b100000000;
assign micromatriz[69][67] = 9'b100000000;
assign micromatriz[69][68] = 9'b100000000;
assign micromatriz[69][69] = 9'b100000000;
assign micromatriz[69][70] = 9'b100100100;
assign micromatriz[69][71] = 9'b100100100;
assign micromatriz[69][72] = 9'b100000000;
assign micromatriz[69][73] = 9'b100000000;
assign micromatriz[69][74] = 9'b100000000;
assign micromatriz[69][75] = 9'b100000000;
assign micromatriz[69][76] = 9'b100000000;
assign micromatriz[69][77] = 9'b100000000;
assign micromatriz[69][78] = 9'b100000000;
assign micromatriz[69][79] = 9'b100000000;
assign micromatriz[69][80] = 9'b100000000;
assign micromatriz[69][81] = 9'b100000000;
assign micromatriz[69][82] = 9'b100000000;
assign micromatriz[69][83] = 9'b101101101;
assign micromatriz[69][84] = 9'b111111111;
assign micromatriz[69][85] = 9'b111111111;
assign micromatriz[69][86] = 9'b111111111;
assign micromatriz[69][87] = 9'b111111111;
assign micromatriz[69][88] = 9'b111111111;
assign micromatriz[69][89] = 9'b111111111;
assign micromatriz[69][90] = 9'b111111111;
assign micromatriz[69][91] = 9'b111111111;
assign micromatriz[69][92] = 9'b111111111;
assign micromatriz[69][93] = 9'b111111111;
assign micromatriz[69][94] = 9'b111111111;
assign micromatriz[69][95] = 9'b111111111;
assign micromatriz[69][96] = 9'b111111111;
assign micromatriz[69][97] = 9'b111111111;
assign micromatriz[69][98] = 9'b111111111;
assign micromatriz[69][99] = 9'b111111111;
assign micromatriz[70][0] = 9'b111111111;
assign micromatriz[70][1] = 9'b111111111;
assign micromatriz[70][2] = 9'b111111111;
assign micromatriz[70][3] = 9'b111111111;
assign micromatriz[70][4] = 9'b111111111;
assign micromatriz[70][5] = 9'b111111111;
assign micromatriz[70][6] = 9'b111111111;
assign micromatriz[70][7] = 9'b111111111;
assign micromatriz[70][8] = 9'b111111111;
assign micromatriz[70][9] = 9'b111111111;
assign micromatriz[70][10] = 9'b111111111;
assign micromatriz[70][11] = 9'b111111111;
assign micromatriz[70][12] = 9'b111111111;
assign micromatriz[70][13] = 9'b111111111;
assign micromatriz[70][14] = 9'b111111111;
assign micromatriz[70][15] = 9'b111111111;
assign micromatriz[70][16] = 9'b101101101;
assign micromatriz[70][17] = 9'b100000000;
assign micromatriz[70][18] = 9'b100000000;
assign micromatriz[70][19] = 9'b100000000;
assign micromatriz[70][20] = 9'b100000000;
assign micromatriz[70][21] = 9'b100000000;
assign micromatriz[70][22] = 9'b100000000;
assign micromatriz[70][23] = 9'b100000000;
assign micromatriz[70][24] = 9'b100000000;
assign micromatriz[70][25] = 9'b100000000;
assign micromatriz[70][26] = 9'b100000000;
assign micromatriz[70][27] = 9'b100000000;
assign micromatriz[70][28] = 9'b100000000;
assign micromatriz[70][29] = 9'b100000000;
assign micromatriz[70][30] = 9'b100000000;
assign micromatriz[70][31] = 9'b100000000;
assign micromatriz[70][32] = 9'b100000000;
assign micromatriz[70][33] = 9'b100000000;
assign micromatriz[70][34] = 9'b100000000;
assign micromatriz[70][35] = 9'b100000000;
assign micromatriz[70][36] = 9'b100000000;
assign micromatriz[70][37] = 9'b100000000;
assign micromatriz[70][38] = 9'b100000000;
assign micromatriz[70][39] = 9'b100000000;
assign micromatriz[70][40] = 9'b100000000;
assign micromatriz[70][41] = 9'b100000000;
assign micromatriz[70][42] = 9'b100000000;
assign micromatriz[70][43] = 9'b100000000;
assign micromatriz[70][44] = 9'b100000000;
assign micromatriz[70][45] = 9'b100000000;
assign micromatriz[70][46] = 9'b100000000;
assign micromatriz[70][47] = 9'b100000000;
assign micromatriz[70][48] = 9'b100000000;
assign micromatriz[70][49] = 9'b100000000;
assign micromatriz[70][50] = 9'b100000000;
assign micromatriz[70][51] = 9'b100000000;
assign micromatriz[70][52] = 9'b100000000;
assign micromatriz[70][53] = 9'b100000000;
assign micromatriz[70][54] = 9'b100000000;
assign micromatriz[70][55] = 9'b100000000;
assign micromatriz[70][56] = 9'b100000000;
assign micromatriz[70][57] = 9'b100000000;
assign micromatriz[70][58] = 9'b100000000;
assign micromatriz[70][59] = 9'b100000000;
assign micromatriz[70][60] = 9'b100000000;
assign micromatriz[70][61] = 9'b100000000;
assign micromatriz[70][62] = 9'b100000000;
assign micromatriz[70][63] = 9'b100000000;
assign micromatriz[70][64] = 9'b100000000;
assign micromatriz[70][65] = 9'b100000000;
assign micromatriz[70][66] = 9'b100000000;
assign micromatriz[70][67] = 9'b100000000;
assign micromatriz[70][68] = 9'b100000000;
assign micromatriz[70][69] = 9'b100000000;
assign micromatriz[70][70] = 9'b100000000;
assign micromatriz[70][71] = 9'b100000000;
assign micromatriz[70][72] = 9'b100000000;
assign micromatriz[70][73] = 9'b100000000;
assign micromatriz[70][74] = 9'b100000000;
assign micromatriz[70][75] = 9'b100000000;
assign micromatriz[70][76] = 9'b100000000;
assign micromatriz[70][77] = 9'b100000000;
assign micromatriz[70][78] = 9'b100000000;
assign micromatriz[70][79] = 9'b100000000;
assign micromatriz[70][80] = 9'b100000000;
assign micromatriz[70][81] = 9'b100000000;
assign micromatriz[70][82] = 9'b100000000;
assign micromatriz[70][83] = 9'b101101101;
assign micromatriz[70][84] = 9'b111111111;
assign micromatriz[70][85] = 9'b111111111;
assign micromatriz[70][86] = 9'b111111111;
assign micromatriz[70][87] = 9'b111111111;
assign micromatriz[70][88] = 9'b111111111;
assign micromatriz[70][89] = 9'b111111111;
assign micromatriz[70][90] = 9'b111111111;
assign micromatriz[70][91] = 9'b111111111;
assign micromatriz[70][92] = 9'b111111111;
assign micromatriz[70][93] = 9'b111111111;
assign micromatriz[70][94] = 9'b111111111;
assign micromatriz[70][95] = 9'b111111111;
assign micromatriz[70][96] = 9'b111111111;
assign micromatriz[70][97] = 9'b111111111;
assign micromatriz[70][98] = 9'b111111111;
assign micromatriz[70][99] = 9'b111111111;
assign micromatriz[71][0] = 9'b111111111;
assign micromatriz[71][1] = 9'b111111111;
assign micromatriz[71][2] = 9'b111111111;
assign micromatriz[71][3] = 9'b111111111;
assign micromatriz[71][4] = 9'b111111111;
assign micromatriz[71][5] = 9'b111111111;
assign micromatriz[71][6] = 9'b111111111;
assign micromatriz[71][7] = 9'b111111111;
assign micromatriz[71][8] = 9'b111111111;
assign micromatriz[71][9] = 9'b111111111;
assign micromatriz[71][10] = 9'b111111111;
assign micromatriz[71][11] = 9'b111111111;
assign micromatriz[71][12] = 9'b111111111;
assign micromatriz[71][13] = 9'b111111111;
assign micromatriz[71][14] = 9'b111111111;
assign micromatriz[71][15] = 9'b111111111;
assign micromatriz[71][16] = 9'b110110110;
assign micromatriz[71][17] = 9'b101101101;
assign micromatriz[71][18] = 9'b101101101;
assign micromatriz[71][19] = 9'b101101101;
assign micromatriz[71][20] = 9'b101101101;
assign micromatriz[71][21] = 9'b101101101;
assign micromatriz[71][22] = 9'b101101101;
assign micromatriz[71][23] = 9'b101101101;
assign micromatriz[71][24] = 9'b101101101;
assign micromatriz[71][25] = 9'b101101101;
assign micromatriz[71][26] = 9'b101101101;
assign micromatriz[71][27] = 9'b101101101;
assign micromatriz[71][28] = 9'b101101101;
assign micromatriz[71][29] = 9'b101101101;
assign micromatriz[71][30] = 9'b101101101;
assign micromatriz[71][31] = 9'b101101101;
assign micromatriz[71][32] = 9'b101101101;
assign micromatriz[71][33] = 9'b101101101;
assign micromatriz[71][34] = 9'b101101101;
assign micromatriz[71][35] = 9'b101101101;
assign micromatriz[71][36] = 9'b101101101;
assign micromatriz[71][37] = 9'b101101101;
assign micromatriz[71][38] = 9'b101101101;
assign micromatriz[71][39] = 9'b101101101;
assign micromatriz[71][40] = 9'b101101101;
assign micromatriz[71][41] = 9'b101101101;
assign micromatriz[71][42] = 9'b101101101;
assign micromatriz[71][43] = 9'b101101101;
assign micromatriz[71][44] = 9'b101101101;
assign micromatriz[71][45] = 9'b101101101;
assign micromatriz[71][46] = 9'b101101101;
assign micromatriz[71][47] = 9'b101101101;
assign micromatriz[71][48] = 9'b101101101;
assign micromatriz[71][49] = 9'b101101101;
assign micromatriz[71][50] = 9'b101101101;
assign micromatriz[71][51] = 9'b101101101;
assign micromatriz[71][52] = 9'b101101101;
assign micromatriz[71][53] = 9'b101101101;
assign micromatriz[71][54] = 9'b101101101;
assign micromatriz[71][55] = 9'b101101101;
assign micromatriz[71][56] = 9'b101101101;
assign micromatriz[71][57] = 9'b101101101;
assign micromatriz[71][58] = 9'b101101101;
assign micromatriz[71][59] = 9'b101101101;
assign micromatriz[71][60] = 9'b101101101;
assign micromatriz[71][61] = 9'b101101101;
assign micromatriz[71][62] = 9'b101101101;
assign micromatriz[71][63] = 9'b101101101;
assign micromatriz[71][64] = 9'b101101101;
assign micromatriz[71][65] = 9'b101101101;
assign micromatriz[71][66] = 9'b101101101;
assign micromatriz[71][67] = 9'b101101101;
assign micromatriz[71][68] = 9'b101101101;
assign micromatriz[71][69] = 9'b101101101;
assign micromatriz[71][70] = 9'b101101101;
assign micromatriz[71][71] = 9'b101101101;
assign micromatriz[71][72] = 9'b101101101;
assign micromatriz[71][73] = 9'b101101101;
assign micromatriz[71][74] = 9'b101101101;
assign micromatriz[71][75] = 9'b101101101;
assign micromatriz[71][76] = 9'b101101101;
assign micromatriz[71][77] = 9'b101101101;
assign micromatriz[71][78] = 9'b101101101;
assign micromatriz[71][79] = 9'b101101101;
assign micromatriz[71][80] = 9'b101101101;
assign micromatriz[71][81] = 9'b101101101;
assign micromatriz[71][82] = 9'b101101101;
assign micromatriz[71][83] = 9'b110110110;
assign micromatriz[71][84] = 9'b111111111;
assign micromatriz[71][85] = 9'b111111111;
assign micromatriz[71][86] = 9'b111111111;
assign micromatriz[71][87] = 9'b111111111;
assign micromatriz[71][88] = 9'b111111111;
assign micromatriz[71][89] = 9'b111111111;
assign micromatriz[71][90] = 9'b111111111;
assign micromatriz[71][91] = 9'b111111111;
assign micromatriz[71][92] = 9'b111111111;
assign micromatriz[71][93] = 9'b111111111;
assign micromatriz[71][94] = 9'b111111111;
assign micromatriz[71][95] = 9'b111111111;
assign micromatriz[71][96] = 9'b111111111;
assign micromatriz[71][97] = 9'b111111111;
assign micromatriz[71][98] = 9'b111111111;
assign micromatriz[71][99] = 9'b111111111;
assign micromatriz[72][0] = 9'b111111111;
assign micromatriz[72][1] = 9'b111111111;
assign micromatriz[72][2] = 9'b111111111;
assign micromatriz[72][3] = 9'b111111111;
assign micromatriz[72][4] = 9'b111111111;
assign micromatriz[72][5] = 9'b111111111;
assign micromatriz[72][6] = 9'b111111111;
assign micromatriz[72][7] = 9'b111111111;
assign micromatriz[72][8] = 9'b111111111;
assign micromatriz[72][9] = 9'b111111111;
assign micromatriz[72][10] = 9'b111111111;
assign micromatriz[72][11] = 9'b111111111;
assign micromatriz[72][12] = 9'b111111111;
assign micromatriz[72][13] = 9'b111111111;
assign micromatriz[72][14] = 9'b111111111;
assign micromatriz[72][15] = 9'b111111111;
assign micromatriz[72][16] = 9'b111111111;
assign micromatriz[72][17] = 9'b111111111;
assign micromatriz[72][18] = 9'b111111111;
assign micromatriz[72][19] = 9'b111111111;
assign micromatriz[72][20] = 9'b111111111;
assign micromatriz[72][21] = 9'b111111111;
assign micromatriz[72][22] = 9'b111111111;
assign micromatriz[72][23] = 9'b111111111;
assign micromatriz[72][24] = 9'b111111111;
assign micromatriz[72][25] = 9'b111111111;
assign micromatriz[72][26] = 9'b111111111;
assign micromatriz[72][27] = 9'b111111111;
assign micromatriz[72][28] = 9'b111111111;
assign micromatriz[72][29] = 9'b111111111;
assign micromatriz[72][30] = 9'b111111111;
assign micromatriz[72][31] = 9'b111111111;
assign micromatriz[72][32] = 9'b111111111;
assign micromatriz[72][33] = 9'b111111111;
assign micromatriz[72][34] = 9'b111111111;
assign micromatriz[72][35] = 9'b111111111;
assign micromatriz[72][36] = 9'b111111111;
assign micromatriz[72][37] = 9'b111111111;
assign micromatriz[72][38] = 9'b111111111;
assign micromatriz[72][39] = 9'b111111111;
assign micromatriz[72][40] = 9'b111111111;
assign micromatriz[72][41] = 9'b111111111;
assign micromatriz[72][42] = 9'b111111111;
assign micromatriz[72][43] = 9'b111111111;
assign micromatriz[72][44] = 9'b111111111;
assign micromatriz[72][45] = 9'b111111111;
assign micromatriz[72][46] = 9'b111111111;
assign micromatriz[72][47] = 9'b111111111;
assign micromatriz[72][48] = 9'b111111111;
assign micromatriz[72][49] = 9'b111111111;
assign micromatriz[72][50] = 9'b111111111;
assign micromatriz[72][51] = 9'b111111111;
assign micromatriz[72][52] = 9'b111111111;
assign micromatriz[72][53] = 9'b111111111;
assign micromatriz[72][54] = 9'b111111111;
assign micromatriz[72][55] = 9'b111111111;
assign micromatriz[72][56] = 9'b111111111;
assign micromatriz[72][57] = 9'b111111111;
assign micromatriz[72][58] = 9'b111111111;
assign micromatriz[72][59] = 9'b111111111;
assign micromatriz[72][60] = 9'b111111111;
assign micromatriz[72][61] = 9'b111111111;
assign micromatriz[72][62] = 9'b111111111;
assign micromatriz[72][63] = 9'b111111111;
assign micromatriz[72][64] = 9'b111111111;
assign micromatriz[72][65] = 9'b111111111;
assign micromatriz[72][66] = 9'b111111111;
assign micromatriz[72][67] = 9'b111111111;
assign micromatriz[72][68] = 9'b111111111;
assign micromatriz[72][69] = 9'b111111111;
assign micromatriz[72][70] = 9'b111111111;
assign micromatriz[72][71] = 9'b111111111;
assign micromatriz[72][72] = 9'b111111111;
assign micromatriz[72][73] = 9'b111111111;
assign micromatriz[72][74] = 9'b111111111;
assign micromatriz[72][75] = 9'b111111111;
assign micromatriz[72][76] = 9'b111111111;
assign micromatriz[72][77] = 9'b111111111;
assign micromatriz[72][78] = 9'b111111111;
assign micromatriz[72][79] = 9'b111111111;
assign micromatriz[72][80] = 9'b111111111;
assign micromatriz[72][81] = 9'b111111111;
assign micromatriz[72][82] = 9'b111111111;
assign micromatriz[72][83] = 9'b111111111;
assign micromatriz[72][84] = 9'b111111111;
assign micromatriz[72][85] = 9'b111111111;
assign micromatriz[72][86] = 9'b111111111;
assign micromatriz[72][87] = 9'b111111111;
assign micromatriz[72][88] = 9'b111111111;
assign micromatriz[72][89] = 9'b111111111;
assign micromatriz[72][90] = 9'b111111111;
assign micromatriz[72][91] = 9'b111111111;
assign micromatriz[72][92] = 9'b111111111;
assign micromatriz[72][93] = 9'b111111111;
assign micromatriz[72][94] = 9'b111111111;
assign micromatriz[72][95] = 9'b111111111;
assign micromatriz[72][96] = 9'b111111111;
assign micromatriz[72][97] = 9'b111111111;
assign micromatriz[72][98] = 9'b111111111;
assign micromatriz[72][99] = 9'b111111111;
assign micromatriz[73][0] = 9'b111111111;
assign micromatriz[73][1] = 9'b111111111;
assign micromatriz[73][2] = 9'b111111111;
assign micromatriz[73][3] = 9'b111111111;
assign micromatriz[73][4] = 9'b111111111;
assign micromatriz[73][5] = 9'b111111111;
assign micromatriz[73][6] = 9'b111111111;
assign micromatriz[73][7] = 9'b111111111;
assign micromatriz[73][8] = 9'b111111111;
assign micromatriz[73][9] = 9'b111111111;
assign micromatriz[73][10] = 9'b111111111;
assign micromatriz[73][11] = 9'b111111111;
assign micromatriz[73][12] = 9'b111111111;
assign micromatriz[73][13] = 9'b111111111;
assign micromatriz[73][14] = 9'b111111111;
assign micromatriz[73][15] = 9'b111111111;
assign micromatriz[73][16] = 9'b111111111;
assign micromatriz[73][17] = 9'b111111111;
assign micromatriz[73][18] = 9'b111111111;
assign micromatriz[73][19] = 9'b111111111;
assign micromatriz[73][20] = 9'b111111111;
assign micromatriz[73][21] = 9'b111111111;
assign micromatriz[73][22] = 9'b111111111;
assign micromatriz[73][23] = 9'b111111111;
assign micromatriz[73][24] = 9'b111111111;
assign micromatriz[73][25] = 9'b111111111;
assign micromatriz[73][26] = 9'b111111111;
assign micromatriz[73][27] = 9'b111111111;
assign micromatriz[73][28] = 9'b111111111;
assign micromatriz[73][29] = 9'b111111111;
assign micromatriz[73][30] = 9'b111111111;
assign micromatriz[73][31] = 9'b111111111;
assign micromatriz[73][32] = 9'b111111111;
assign micromatriz[73][33] = 9'b111111111;
assign micromatriz[73][34] = 9'b111111111;
assign micromatriz[73][35] = 9'b111111111;
assign micromatriz[73][36] = 9'b111111111;
assign micromatriz[73][37] = 9'b111111111;
assign micromatriz[73][38] = 9'b111111111;
assign micromatriz[73][39] = 9'b111111111;
assign micromatriz[73][40] = 9'b111111111;
assign micromatriz[73][41] = 9'b111111111;
assign micromatriz[73][42] = 9'b111111111;
assign micromatriz[73][43] = 9'b111111111;
assign micromatriz[73][44] = 9'b111111111;
assign micromatriz[73][45] = 9'b111111111;
assign micromatriz[73][46] = 9'b111111111;
assign micromatriz[73][47] = 9'b111111111;
assign micromatriz[73][48] = 9'b111111111;
assign micromatriz[73][49] = 9'b111111111;
assign micromatriz[73][50] = 9'b111111111;
assign micromatriz[73][51] = 9'b111111111;
assign micromatriz[73][52] = 9'b111111111;
assign micromatriz[73][53] = 9'b111111111;
assign micromatriz[73][54] = 9'b111111111;
assign micromatriz[73][55] = 9'b111111111;
assign micromatriz[73][56] = 9'b111111111;
assign micromatriz[73][57] = 9'b111111111;
assign micromatriz[73][58] = 9'b111111111;
assign micromatriz[73][59] = 9'b111111111;
assign micromatriz[73][60] = 9'b111111111;
assign micromatriz[73][61] = 9'b111111111;
assign micromatriz[73][62] = 9'b111111111;
assign micromatriz[73][63] = 9'b111111111;
assign micromatriz[73][64] = 9'b111111111;
assign micromatriz[73][65] = 9'b111111111;
assign micromatriz[73][66] = 9'b111111111;
assign micromatriz[73][67] = 9'b111111111;
assign micromatriz[73][68] = 9'b111111111;
assign micromatriz[73][69] = 9'b111111111;
assign micromatriz[73][70] = 9'b111111111;
assign micromatriz[73][71] = 9'b111111111;
assign micromatriz[73][72] = 9'b111111111;
assign micromatriz[73][73] = 9'b111111111;
assign micromatriz[73][74] = 9'b111111111;
assign micromatriz[73][75] = 9'b111111111;
assign micromatriz[73][76] = 9'b111111111;
assign micromatriz[73][77] = 9'b111111111;
assign micromatriz[73][78] = 9'b111111111;
assign micromatriz[73][79] = 9'b111111111;
assign micromatriz[73][80] = 9'b111111111;
assign micromatriz[73][81] = 9'b111111111;
assign micromatriz[73][82] = 9'b111111111;
assign micromatriz[73][83] = 9'b111111111;
assign micromatriz[73][84] = 9'b111111111;
assign micromatriz[73][85] = 9'b111111111;
assign micromatriz[73][86] = 9'b111111111;
assign micromatriz[73][87] = 9'b111111111;
assign micromatriz[73][88] = 9'b111111111;
assign micromatriz[73][89] = 9'b111111111;
assign micromatriz[73][90] = 9'b111111111;
assign micromatriz[73][91] = 9'b111111111;
assign micromatriz[73][92] = 9'b111111111;
assign micromatriz[73][93] = 9'b111111111;
assign micromatriz[73][94] = 9'b111111111;
assign micromatriz[73][95] = 9'b111111111;
assign micromatriz[73][96] = 9'b111111111;
assign micromatriz[73][97] = 9'b111111111;
assign micromatriz[73][98] = 9'b111111111;
assign micromatriz[73][99] = 9'b111111111;
assign micromatriz[74][0] = 9'b111111111;
assign micromatriz[74][1] = 9'b111111111;
assign micromatriz[74][2] = 9'b111111111;
assign micromatriz[74][3] = 9'b111111111;
assign micromatriz[74][4] = 9'b111111111;
assign micromatriz[74][5] = 9'b111111111;
assign micromatriz[74][6] = 9'b111111111;
assign micromatriz[74][7] = 9'b111111111;
assign micromatriz[74][8] = 9'b111111111;
assign micromatriz[74][9] = 9'b111111111;
assign micromatriz[74][10] = 9'b111111111;
assign micromatriz[74][11] = 9'b111111111;
assign micromatriz[74][12] = 9'b111111111;
assign micromatriz[74][13] = 9'b111111111;
assign micromatriz[74][14] = 9'b111111111;
assign micromatriz[74][15] = 9'b111111111;
assign micromatriz[74][16] = 9'b111111111;
assign micromatriz[74][17] = 9'b111111111;
assign micromatriz[74][18] = 9'b111111111;
assign micromatriz[74][19] = 9'b111111111;
assign micromatriz[74][20] = 9'b111111111;
assign micromatriz[74][21] = 9'b111111111;
assign micromatriz[74][22] = 9'b111111111;
assign micromatriz[74][23] = 9'b111111111;
assign micromatriz[74][24] = 9'b111111111;
assign micromatriz[74][25] = 9'b111111111;
assign micromatriz[74][26] = 9'b111111111;
assign micromatriz[74][27] = 9'b111111111;
assign micromatriz[74][28] = 9'b111111111;
assign micromatriz[74][29] = 9'b111111111;
assign micromatriz[74][30] = 9'b111111111;
assign micromatriz[74][31] = 9'b111111111;
assign micromatriz[74][32] = 9'b111111111;
assign micromatriz[74][33] = 9'b111111111;
assign micromatriz[74][34] = 9'b111111111;
assign micromatriz[74][35] = 9'b111111111;
assign micromatriz[74][36] = 9'b111111111;
assign micromatriz[74][37] = 9'b111111111;
assign micromatriz[74][38] = 9'b111111111;
assign micromatriz[74][39] = 9'b111111111;
assign micromatriz[74][40] = 9'b111111111;
assign micromatriz[74][41] = 9'b111111111;
assign micromatriz[74][42] = 9'b111111111;
assign micromatriz[74][43] = 9'b111111111;
assign micromatriz[74][44] = 9'b111111111;
assign micromatriz[74][45] = 9'b111111111;
assign micromatriz[74][46] = 9'b111111111;
assign micromatriz[74][47] = 9'b111111111;
assign micromatriz[74][48] = 9'b111111111;
assign micromatriz[74][49] = 9'b111111111;
assign micromatriz[74][50] = 9'b111111111;
assign micromatriz[74][51] = 9'b111111111;
assign micromatriz[74][52] = 9'b111111111;
assign micromatriz[74][53] = 9'b111111111;
assign micromatriz[74][54] = 9'b111111111;
assign micromatriz[74][55] = 9'b111111111;
assign micromatriz[74][56] = 9'b111111111;
assign micromatriz[74][57] = 9'b111111111;
assign micromatriz[74][58] = 9'b111111111;
assign micromatriz[74][59] = 9'b111111111;
assign micromatriz[74][60] = 9'b111111111;
assign micromatriz[74][61] = 9'b111111111;
assign micromatriz[74][62] = 9'b111111111;
assign micromatriz[74][63] = 9'b111111111;
assign micromatriz[74][64] = 9'b111111111;
assign micromatriz[74][65] = 9'b111111111;
assign micromatriz[74][66] = 9'b111111111;
assign micromatriz[74][67] = 9'b111111111;
assign micromatriz[74][68] = 9'b111111111;
assign micromatriz[74][69] = 9'b111111111;
assign micromatriz[74][70] = 9'b111111111;
assign micromatriz[74][71] = 9'b111111111;
assign micromatriz[74][72] = 9'b111111111;
assign micromatriz[74][73] = 9'b111111111;
assign micromatriz[74][74] = 9'b111111111;
assign micromatriz[74][75] = 9'b111111111;
assign micromatriz[74][76] = 9'b111111111;
assign micromatriz[74][77] = 9'b111111111;
assign micromatriz[74][78] = 9'b111111111;
assign micromatriz[74][79] = 9'b111111111;
assign micromatriz[74][80] = 9'b111111111;
assign micromatriz[74][81] = 9'b111111111;
assign micromatriz[74][82] = 9'b111111111;
assign micromatriz[74][83] = 9'b111111111;
assign micromatriz[74][84] = 9'b111111111;
assign micromatriz[74][85] = 9'b111111111;
assign micromatriz[74][86] = 9'b111111111;
assign micromatriz[74][87] = 9'b111111111;
assign micromatriz[74][88] = 9'b111111111;
assign micromatriz[74][89] = 9'b111111111;
assign micromatriz[74][90] = 9'b111111111;
assign micromatriz[74][91] = 9'b111111111;
assign micromatriz[74][92] = 9'b111111111;
assign micromatriz[74][93] = 9'b111111111;
assign micromatriz[74][94] = 9'b111111111;
assign micromatriz[74][95] = 9'b111111111;
assign micromatriz[74][96] = 9'b111111111;
assign micromatriz[74][97] = 9'b111111111;
assign micromatriz[74][98] = 9'b111111111;
assign micromatriz[74][99] = 9'b111111111;
assign micromatriz[75][0] = 9'b111111111;
assign micromatriz[75][1] = 9'b111111111;
assign micromatriz[75][2] = 9'b111111111;
assign micromatriz[75][3] = 9'b111111111;
assign micromatriz[75][4] = 9'b111111111;
assign micromatriz[75][5] = 9'b111111111;
assign micromatriz[75][6] = 9'b111111111;
assign micromatriz[75][7] = 9'b111111111;
assign micromatriz[75][8] = 9'b111111111;
assign micromatriz[75][9] = 9'b111111111;
assign micromatriz[75][10] = 9'b111111111;
assign micromatriz[75][11] = 9'b111111111;
assign micromatriz[75][12] = 9'b111111111;
assign micromatriz[75][13] = 9'b111111111;
assign micromatriz[75][14] = 9'b111111111;
assign micromatriz[75][15] = 9'b111111111;
assign micromatriz[75][16] = 9'b111111111;
assign micromatriz[75][17] = 9'b111111111;
assign micromatriz[75][18] = 9'b111111111;
assign micromatriz[75][19] = 9'b111111111;
assign micromatriz[75][20] = 9'b111111111;
assign micromatriz[75][21] = 9'b111111111;
assign micromatriz[75][22] = 9'b111111111;
assign micromatriz[75][23] = 9'b111111111;
assign micromatriz[75][24] = 9'b111111111;
assign micromatriz[75][25] = 9'b111111111;
assign micromatriz[75][26] = 9'b111111111;
assign micromatriz[75][27] = 9'b111111111;
assign micromatriz[75][28] = 9'b111111111;
assign micromatriz[75][29] = 9'b111111111;
assign micromatriz[75][30] = 9'b111111111;
assign micromatriz[75][31] = 9'b111111111;
assign micromatriz[75][32] = 9'b111111111;
assign micromatriz[75][33] = 9'b111111111;
assign micromatriz[75][34] = 9'b111111111;
assign micromatriz[75][35] = 9'b111111111;
assign micromatriz[75][36] = 9'b111111111;
assign micromatriz[75][37] = 9'b111111111;
assign micromatriz[75][38] = 9'b111111111;
assign micromatriz[75][39] = 9'b111111111;
assign micromatriz[75][40] = 9'b111111111;
assign micromatriz[75][41] = 9'b111111111;
assign micromatriz[75][42] = 9'b111111111;
assign micromatriz[75][43] = 9'b111111111;
assign micromatriz[75][44] = 9'b111111111;
assign micromatriz[75][45] = 9'b111111111;
assign micromatriz[75][46] = 9'b111111111;
assign micromatriz[75][47] = 9'b111111111;
assign micromatriz[75][48] = 9'b111111111;
assign micromatriz[75][49] = 9'b111111111;
assign micromatriz[75][50] = 9'b111111111;
assign micromatriz[75][51] = 9'b111111111;
assign micromatriz[75][52] = 9'b111111111;
assign micromatriz[75][53] = 9'b111111111;
assign micromatriz[75][54] = 9'b111111111;
assign micromatriz[75][55] = 9'b111111111;
assign micromatriz[75][56] = 9'b111111111;
assign micromatriz[75][57] = 9'b111111111;
assign micromatriz[75][58] = 9'b111111111;
assign micromatriz[75][59] = 9'b111111111;
assign micromatriz[75][60] = 9'b111111111;
assign micromatriz[75][61] = 9'b111111111;
assign micromatriz[75][62] = 9'b111111111;
assign micromatriz[75][63] = 9'b111111111;
assign micromatriz[75][64] = 9'b111111111;
assign micromatriz[75][65] = 9'b111111111;
assign micromatriz[75][66] = 9'b111111111;
assign micromatriz[75][67] = 9'b111111111;
assign micromatriz[75][68] = 9'b111111111;
assign micromatriz[75][69] = 9'b111111111;
assign micromatriz[75][70] = 9'b111111111;
assign micromatriz[75][71] = 9'b111111111;
assign micromatriz[75][72] = 9'b111111111;
assign micromatriz[75][73] = 9'b111111111;
assign micromatriz[75][74] = 9'b111111111;
assign micromatriz[75][75] = 9'b111111111;
assign micromatriz[75][76] = 9'b111111111;
assign micromatriz[75][77] = 9'b111111111;
assign micromatriz[75][78] = 9'b111111111;
assign micromatriz[75][79] = 9'b111111111;
assign micromatriz[75][80] = 9'b111111111;
assign micromatriz[75][81] = 9'b111111111;
assign micromatriz[75][82] = 9'b111111111;
assign micromatriz[75][83] = 9'b111111111;
assign micromatriz[75][84] = 9'b111111111;
assign micromatriz[75][85] = 9'b111111111;
assign micromatriz[75][86] = 9'b111111111;
assign micromatriz[75][87] = 9'b111111111;
assign micromatriz[75][88] = 9'b111111111;
assign micromatriz[75][89] = 9'b111111111;
assign micromatriz[75][90] = 9'b111111111;
assign micromatriz[75][91] = 9'b111111111;
assign micromatriz[75][92] = 9'b111111111;
assign micromatriz[75][93] = 9'b111111111;
assign micromatriz[75][94] = 9'b111111111;
assign micromatriz[75][95] = 9'b111111111;
assign micromatriz[75][96] = 9'b111111111;
assign micromatriz[75][97] = 9'b111111111;
assign micromatriz[75][98] = 9'b111111111;
assign micromatriz[75][99] = 9'b111111111;
assign micromatriz[76][0] = 9'b111111111;
assign micromatriz[76][1] = 9'b111111111;
assign micromatriz[76][2] = 9'b111111111;
assign micromatriz[76][3] = 9'b111111111;
assign micromatriz[76][4] = 9'b111111111;
assign micromatriz[76][5] = 9'b111111111;
assign micromatriz[76][6] = 9'b111111111;
assign micromatriz[76][7] = 9'b111111111;
assign micromatriz[76][8] = 9'b111111111;
assign micromatriz[76][9] = 9'b111111111;
assign micromatriz[76][10] = 9'b111111111;
assign micromatriz[76][11] = 9'b111111111;
assign micromatriz[76][12] = 9'b111111111;
assign micromatriz[76][13] = 9'b111111111;
assign micromatriz[76][14] = 9'b111111111;
assign micromatriz[76][15] = 9'b111111111;
assign micromatriz[76][16] = 9'b111111111;
assign micromatriz[76][17] = 9'b111111111;
assign micromatriz[76][18] = 9'b111111111;
assign micromatriz[76][19] = 9'b111111111;
assign micromatriz[76][20] = 9'b111111111;
assign micromatriz[76][21] = 9'b111111111;
assign micromatriz[76][22] = 9'b111111111;
assign micromatriz[76][23] = 9'b111111111;
assign micromatriz[76][24] = 9'b111111111;
assign micromatriz[76][25] = 9'b111111111;
assign micromatriz[76][26] = 9'b111111111;
assign micromatriz[76][27] = 9'b111111111;
assign micromatriz[76][28] = 9'b111111111;
assign micromatriz[76][29] = 9'b111111111;
assign micromatriz[76][30] = 9'b111111111;
assign micromatriz[76][31] = 9'b111111111;
assign micromatriz[76][32] = 9'b111111111;
assign micromatriz[76][33] = 9'b111111111;
assign micromatriz[76][34] = 9'b111111111;
assign micromatriz[76][35] = 9'b111111111;
assign micromatriz[76][36] = 9'b111111111;
assign micromatriz[76][37] = 9'b111111111;
assign micromatriz[76][38] = 9'b111111111;
assign micromatriz[76][39] = 9'b111111111;
assign micromatriz[76][40] = 9'b111111111;
assign micromatriz[76][41] = 9'b111111111;
assign micromatriz[76][42] = 9'b111111111;
assign micromatriz[76][43] = 9'b111111111;
assign micromatriz[76][44] = 9'b111111111;
assign micromatriz[76][45] = 9'b111111111;
assign micromatriz[76][46] = 9'b111111111;
assign micromatriz[76][47] = 9'b111111111;
assign micromatriz[76][48] = 9'b111111111;
assign micromatriz[76][49] = 9'b111111111;
assign micromatriz[76][50] = 9'b111111111;
assign micromatriz[76][51] = 9'b111111111;
assign micromatriz[76][52] = 9'b111111111;
assign micromatriz[76][53] = 9'b111111111;
assign micromatriz[76][54] = 9'b111111111;
assign micromatriz[76][55] = 9'b111111111;
assign micromatriz[76][56] = 9'b111111111;
assign micromatriz[76][57] = 9'b111111111;
assign micromatriz[76][58] = 9'b111111111;
assign micromatriz[76][59] = 9'b111111111;
assign micromatriz[76][60] = 9'b111111111;
assign micromatriz[76][61] = 9'b111111111;
assign micromatriz[76][62] = 9'b111111111;
assign micromatriz[76][63] = 9'b111111111;
assign micromatriz[76][64] = 9'b111111111;
assign micromatriz[76][65] = 9'b111111111;
assign micromatriz[76][66] = 9'b111111111;
assign micromatriz[76][67] = 9'b111111111;
assign micromatriz[76][68] = 9'b111111111;
assign micromatriz[76][69] = 9'b111111111;
assign micromatriz[76][70] = 9'b111111111;
assign micromatriz[76][71] = 9'b111111111;
assign micromatriz[76][72] = 9'b111111111;
assign micromatriz[76][73] = 9'b111111111;
assign micromatriz[76][74] = 9'b111111111;
assign micromatriz[76][75] = 9'b111111111;
assign micromatriz[76][76] = 9'b111111111;
assign micromatriz[76][77] = 9'b111111111;
assign micromatriz[76][78] = 9'b111111111;
assign micromatriz[76][79] = 9'b111111111;
assign micromatriz[76][80] = 9'b111111111;
assign micromatriz[76][81] = 9'b111111111;
assign micromatriz[76][82] = 9'b111111111;
assign micromatriz[76][83] = 9'b111111111;
assign micromatriz[76][84] = 9'b111111111;
assign micromatriz[76][85] = 9'b111111111;
assign micromatriz[76][86] = 9'b111111111;
assign micromatriz[76][87] = 9'b111111111;
assign micromatriz[76][88] = 9'b111111111;
assign micromatriz[76][89] = 9'b111111111;
assign micromatriz[76][90] = 9'b111111111;
assign micromatriz[76][91] = 9'b111111111;
assign micromatriz[76][92] = 9'b111111111;
assign micromatriz[76][93] = 9'b111111111;
assign micromatriz[76][94] = 9'b111111111;
assign micromatriz[76][95] = 9'b111111111;
assign micromatriz[76][96] = 9'b111111111;
assign micromatriz[76][97] = 9'b111111111;
assign micromatriz[76][98] = 9'b111111111;
assign micromatriz[76][99] = 9'b111111111;
assign micromatriz[77][0] = 9'b111111111;
assign micromatriz[77][1] = 9'b111111111;
assign micromatriz[77][2] = 9'b111111111;
assign micromatriz[77][3] = 9'b111111111;
assign micromatriz[77][4] = 9'b111111111;
assign micromatriz[77][5] = 9'b111111111;
assign micromatriz[77][6] = 9'b111111111;
assign micromatriz[77][7] = 9'b111111111;
assign micromatriz[77][8] = 9'b111111111;
assign micromatriz[77][9] = 9'b111111111;
assign micromatriz[77][10] = 9'b111111111;
assign micromatriz[77][11] = 9'b111111111;
assign micromatriz[77][12] = 9'b111111111;
assign micromatriz[77][13] = 9'b111111111;
assign micromatriz[77][14] = 9'b111111111;
assign micromatriz[77][15] = 9'b111111111;
assign micromatriz[77][16] = 9'b111111111;
assign micromatriz[77][17] = 9'b111111111;
assign micromatriz[77][18] = 9'b111111111;
assign micromatriz[77][19] = 9'b111111111;
assign micromatriz[77][20] = 9'b111111111;
assign micromatriz[77][21] = 9'b111111111;
assign micromatriz[77][22] = 9'b111111111;
assign micromatriz[77][23] = 9'b111111111;
assign micromatriz[77][24] = 9'b111111111;
assign micromatriz[77][25] = 9'b111111111;
assign micromatriz[77][26] = 9'b111111111;
assign micromatriz[77][27] = 9'b111111111;
assign micromatriz[77][28] = 9'b111111111;
assign micromatriz[77][29] = 9'b111111111;
assign micromatriz[77][30] = 9'b111111111;
assign micromatriz[77][31] = 9'b111111111;
assign micromatriz[77][32] = 9'b111111111;
assign micromatriz[77][33] = 9'b111111111;
assign micromatriz[77][34] = 9'b111111111;
assign micromatriz[77][35] = 9'b111111111;
assign micromatriz[77][36] = 9'b111111111;
assign micromatriz[77][37] = 9'b111111111;
assign micromatriz[77][38] = 9'b111111111;
assign micromatriz[77][39] = 9'b111111111;
assign micromatriz[77][40] = 9'b111111111;
assign micromatriz[77][41] = 9'b111111111;
assign micromatriz[77][42] = 9'b111111111;
assign micromatriz[77][43] = 9'b111111111;
assign micromatriz[77][44] = 9'b111111111;
assign micromatriz[77][45] = 9'b111111111;
assign micromatriz[77][46] = 9'b111111111;
assign micromatriz[77][47] = 9'b111111111;
assign micromatriz[77][48] = 9'b111111111;
assign micromatriz[77][49] = 9'b111111111;
assign micromatriz[77][50] = 9'b111111111;
assign micromatriz[77][51] = 9'b111111111;
assign micromatriz[77][52] = 9'b111111111;
assign micromatriz[77][53] = 9'b111111111;
assign micromatriz[77][54] = 9'b111111111;
assign micromatriz[77][55] = 9'b111111111;
assign micromatriz[77][56] = 9'b111111111;
assign micromatriz[77][57] = 9'b111111111;
assign micromatriz[77][58] = 9'b111111111;
assign micromatriz[77][59] = 9'b111111111;
assign micromatriz[77][60] = 9'b111111111;
assign micromatriz[77][61] = 9'b111111111;
assign micromatriz[77][62] = 9'b111111111;
assign micromatriz[77][63] = 9'b111111111;
assign micromatriz[77][64] = 9'b111111111;
assign micromatriz[77][65] = 9'b111111111;
assign micromatriz[77][66] = 9'b111111111;
assign micromatriz[77][67] = 9'b111111111;
assign micromatriz[77][68] = 9'b111111111;
assign micromatriz[77][69] = 9'b111111111;
assign micromatriz[77][70] = 9'b111111111;
assign micromatriz[77][71] = 9'b111111111;
assign micromatriz[77][72] = 9'b111111111;
assign micromatriz[77][73] = 9'b111111111;
assign micromatriz[77][74] = 9'b111111111;
assign micromatriz[77][75] = 9'b111111111;
assign micromatriz[77][76] = 9'b111111111;
assign micromatriz[77][77] = 9'b111111111;
assign micromatriz[77][78] = 9'b111111111;
assign micromatriz[77][79] = 9'b111111111;
assign micromatriz[77][80] = 9'b111111111;
assign micromatriz[77][81] = 9'b111111111;
assign micromatriz[77][82] = 9'b111111111;
assign micromatriz[77][83] = 9'b111111111;
assign micromatriz[77][84] = 9'b111111111;
assign micromatriz[77][85] = 9'b111111111;
assign micromatriz[77][86] = 9'b111111111;
assign micromatriz[77][87] = 9'b111111111;
assign micromatriz[77][88] = 9'b111111111;
assign micromatriz[77][89] = 9'b111111111;
assign micromatriz[77][90] = 9'b111111111;
assign micromatriz[77][91] = 9'b111111111;
assign micromatriz[77][92] = 9'b111111111;
assign micromatriz[77][93] = 9'b111111111;
assign micromatriz[77][94] = 9'b111111111;
assign micromatriz[77][95] = 9'b111111111;
assign micromatriz[77][96] = 9'b111111111;
assign micromatriz[77][97] = 9'b111111111;
assign micromatriz[77][98] = 9'b111111111;
assign micromatriz[77][99] = 9'b111111111;
assign micromatriz[78][0] = 9'b111111111;
assign micromatriz[78][1] = 9'b111111111;
assign micromatriz[78][2] = 9'b111111111;
assign micromatriz[78][3] = 9'b111111111;
assign micromatriz[78][4] = 9'b111111111;
assign micromatriz[78][5] = 9'b111111111;
assign micromatriz[78][6] = 9'b111111111;
assign micromatriz[78][7] = 9'b111111111;
assign micromatriz[78][8] = 9'b111111111;
assign micromatriz[78][9] = 9'b111111111;
assign micromatriz[78][10] = 9'b111111111;
assign micromatriz[78][11] = 9'b111111111;
assign micromatriz[78][12] = 9'b111111111;
assign micromatriz[78][13] = 9'b111111111;
assign micromatriz[78][14] = 9'b111111111;
assign micromatriz[78][15] = 9'b111111111;
assign micromatriz[78][16] = 9'b111111111;
assign micromatriz[78][17] = 9'b111111111;
assign micromatriz[78][18] = 9'b111111111;
assign micromatriz[78][19] = 9'b111111111;
assign micromatriz[78][20] = 9'b111111111;
assign micromatriz[78][21] = 9'b111111111;
assign micromatriz[78][22] = 9'b111111111;
assign micromatriz[78][23] = 9'b111111111;
assign micromatriz[78][24] = 9'b111111111;
assign micromatriz[78][25] = 9'b111111111;
assign micromatriz[78][26] = 9'b111111111;
assign micromatriz[78][27] = 9'b111111111;
assign micromatriz[78][28] = 9'b111111111;
assign micromatriz[78][29] = 9'b111111111;
assign micromatriz[78][30] = 9'b111111111;
assign micromatriz[78][31] = 9'b111111111;
assign micromatriz[78][32] = 9'b111111111;
assign micromatriz[78][33] = 9'b111111111;
assign micromatriz[78][34] = 9'b111111111;
assign micromatriz[78][35] = 9'b111111111;
assign micromatriz[78][36] = 9'b111111111;
assign micromatriz[78][37] = 9'b111111111;
assign micromatriz[78][38] = 9'b111111111;
assign micromatriz[78][39] = 9'b111111111;
assign micromatriz[78][40] = 9'b111111111;
assign micromatriz[78][41] = 9'b111111111;
assign micromatriz[78][42] = 9'b111111111;
assign micromatriz[78][43] = 9'b111111111;
assign micromatriz[78][44] = 9'b111111111;
assign micromatriz[78][45] = 9'b111111111;
assign micromatriz[78][46] = 9'b111111111;
assign micromatriz[78][47] = 9'b111111111;
assign micromatriz[78][48] = 9'b111111111;
assign micromatriz[78][49] = 9'b111111111;
assign micromatriz[78][50] = 9'b111111111;
assign micromatriz[78][51] = 9'b111111111;
assign micromatriz[78][52] = 9'b111111111;
assign micromatriz[78][53] = 9'b111111111;
assign micromatriz[78][54] = 9'b111111111;
assign micromatriz[78][55] = 9'b111111111;
assign micromatriz[78][56] = 9'b111111111;
assign micromatriz[78][57] = 9'b111111111;
assign micromatriz[78][58] = 9'b111111111;
assign micromatriz[78][59] = 9'b111111111;
assign micromatriz[78][60] = 9'b111111111;
assign micromatriz[78][61] = 9'b111111111;
assign micromatriz[78][62] = 9'b111111111;
assign micromatriz[78][63] = 9'b111111111;
assign micromatriz[78][64] = 9'b111111111;
assign micromatriz[78][65] = 9'b111111111;
assign micromatriz[78][66] = 9'b111111111;
assign micromatriz[78][67] = 9'b111111111;
assign micromatriz[78][68] = 9'b111111111;
assign micromatriz[78][69] = 9'b111111111;
assign micromatriz[78][70] = 9'b111111111;
assign micromatriz[78][71] = 9'b111111111;
assign micromatriz[78][72] = 9'b111111111;
assign micromatriz[78][73] = 9'b111111111;
assign micromatriz[78][74] = 9'b111111111;
assign micromatriz[78][75] = 9'b111111111;
assign micromatriz[78][76] = 9'b111111111;
assign micromatriz[78][77] = 9'b111111111;
assign micromatriz[78][78] = 9'b111111111;
assign micromatriz[78][79] = 9'b111111111;
assign micromatriz[78][80] = 9'b111111111;
assign micromatriz[78][81] = 9'b111111111;
assign micromatriz[78][82] = 9'b111111111;
assign micromatriz[78][83] = 9'b111111111;
assign micromatriz[78][84] = 9'b111111111;
assign micromatriz[78][85] = 9'b111111111;
assign micromatriz[78][86] = 9'b111111111;
assign micromatriz[78][87] = 9'b111111111;
assign micromatriz[78][88] = 9'b111111111;
assign micromatriz[78][89] = 9'b111111111;
assign micromatriz[78][90] = 9'b111111111;
assign micromatriz[78][91] = 9'b111111111;
assign micromatriz[78][92] = 9'b111111111;
assign micromatriz[78][93] = 9'b111111111;
assign micromatriz[78][94] = 9'b111111111;
assign micromatriz[78][95] = 9'b111111111;
assign micromatriz[78][96] = 9'b111111111;
assign micromatriz[78][97] = 9'b111111111;
assign micromatriz[78][98] = 9'b111111111;
assign micromatriz[78][99] = 9'b111111111;
assign micromatriz[79][0] = 9'b111111111;
assign micromatriz[79][1] = 9'b111111111;
assign micromatriz[79][2] = 9'b111111111;
assign micromatriz[79][3] = 9'b111111111;
assign micromatriz[79][4] = 9'b111111111;
assign micromatriz[79][5] = 9'b111111111;
assign micromatriz[79][6] = 9'b111111111;
assign micromatriz[79][7] = 9'b111111111;
assign micromatriz[79][8] = 9'b111111111;
assign micromatriz[79][9] = 9'b111111111;
assign micromatriz[79][10] = 9'b111111111;
assign micromatriz[79][11] = 9'b111111111;
assign micromatriz[79][12] = 9'b111111111;
assign micromatriz[79][13] = 9'b111111111;
assign micromatriz[79][14] = 9'b111111111;
assign micromatriz[79][15] = 9'b111111111;
assign micromatriz[79][16] = 9'b111111111;
assign micromatriz[79][17] = 9'b111111111;
assign micromatriz[79][18] = 9'b111111111;
assign micromatriz[79][19] = 9'b111111111;
assign micromatriz[79][20] = 9'b111111111;
assign micromatriz[79][21] = 9'b111111111;
assign micromatriz[79][22] = 9'b111111111;
assign micromatriz[79][23] = 9'b111111111;
assign micromatriz[79][24] = 9'b111111111;
assign micromatriz[79][25] = 9'b111111111;
assign micromatriz[79][26] = 9'b111111111;
assign micromatriz[79][27] = 9'b111111111;
assign micromatriz[79][28] = 9'b111111111;
assign micromatriz[79][29] = 9'b111111111;
assign micromatriz[79][30] = 9'b111111111;
assign micromatriz[79][31] = 9'b111111111;
assign micromatriz[79][32] = 9'b111111111;
assign micromatriz[79][33] = 9'b111111111;
assign micromatriz[79][34] = 9'b111111111;
assign micromatriz[79][35] = 9'b111111111;
assign micromatriz[79][36] = 9'b111111111;
assign micromatriz[79][37] = 9'b111111111;
assign micromatriz[79][38] = 9'b111111111;
assign micromatriz[79][39] = 9'b111111111;
assign micromatriz[79][40] = 9'b111111111;
assign micromatriz[79][41] = 9'b111111111;
assign micromatriz[79][42] = 9'b111111111;
assign micromatriz[79][43] = 9'b111111111;
assign micromatriz[79][44] = 9'b111111111;
assign micromatriz[79][45] = 9'b111111111;
assign micromatriz[79][46] = 9'b111111111;
assign micromatriz[79][47] = 9'b111111111;
assign micromatriz[79][48] = 9'b111111111;
assign micromatriz[79][49] = 9'b111111111;
assign micromatriz[79][50] = 9'b111111111;
assign micromatriz[79][51] = 9'b111111111;
assign micromatriz[79][52] = 9'b111111111;
assign micromatriz[79][53] = 9'b111111111;
assign micromatriz[79][54] = 9'b111111111;
assign micromatriz[79][55] = 9'b111111111;
assign micromatriz[79][56] = 9'b111111111;
assign micromatriz[79][57] = 9'b111111111;
assign micromatriz[79][58] = 9'b111111111;
assign micromatriz[79][59] = 9'b111111111;
assign micromatriz[79][60] = 9'b111111111;
assign micromatriz[79][61] = 9'b111111111;
assign micromatriz[79][62] = 9'b111111111;
assign micromatriz[79][63] = 9'b111111111;
assign micromatriz[79][64] = 9'b111111111;
assign micromatriz[79][65] = 9'b111111111;
assign micromatriz[79][66] = 9'b111111111;
assign micromatriz[79][67] = 9'b111111111;
assign micromatriz[79][68] = 9'b111111111;
assign micromatriz[79][69] = 9'b111111111;
assign micromatriz[79][70] = 9'b111111111;
assign micromatriz[79][71] = 9'b111111111;
assign micromatriz[79][72] = 9'b111111111;
assign micromatriz[79][73] = 9'b111111111;
assign micromatriz[79][74] = 9'b111111111;
assign micromatriz[79][75] = 9'b111111111;
assign micromatriz[79][76] = 9'b111111111;
assign micromatriz[79][77] = 9'b111111111;
assign micromatriz[79][78] = 9'b111111111;
assign micromatriz[79][79] = 9'b111111111;
assign micromatriz[79][80] = 9'b111111111;
assign micromatriz[79][81] = 9'b111111111;
assign micromatriz[79][82] = 9'b111111111;
assign micromatriz[79][83] = 9'b111111111;
assign micromatriz[79][84] = 9'b111111111;
assign micromatriz[79][85] = 9'b111111111;
assign micromatriz[79][86] = 9'b111111111;
assign micromatriz[79][87] = 9'b111111111;
assign micromatriz[79][88] = 9'b111111111;
assign micromatriz[79][89] = 9'b111111111;
assign micromatriz[79][90] = 9'b111111111;
assign micromatriz[79][91] = 9'b111111111;
assign micromatriz[79][92] = 9'b111111111;
assign micromatriz[79][93] = 9'b111111111;
assign micromatriz[79][94] = 9'b111111111;
assign micromatriz[79][95] = 9'b111111111;
assign micromatriz[79][96] = 9'b111111111;
assign micromatriz[79][97] = 9'b111111111;
assign micromatriz[79][98] = 9'b111111111;
assign micromatriz[79][99] = 9'b111111111;
assign micromatriz[80][0] = 9'b111111111;
assign micromatriz[80][1] = 9'b111111111;
assign micromatriz[80][2] = 9'b111111111;
assign micromatriz[80][3] = 9'b111111111;
assign micromatriz[80][4] = 9'b111111111;
assign micromatriz[80][5] = 9'b111111111;
assign micromatriz[80][6] = 9'b111111111;
assign micromatriz[80][7] = 9'b111111111;
assign micromatriz[80][8] = 9'b111111111;
assign micromatriz[80][9] = 9'b111111111;
assign micromatriz[80][10] = 9'b111111111;
assign micromatriz[80][11] = 9'b111111111;
assign micromatriz[80][12] = 9'b111111111;
assign micromatriz[80][13] = 9'b111111111;
assign micromatriz[80][14] = 9'b111111111;
assign micromatriz[80][15] = 9'b111111111;
assign micromatriz[80][16] = 9'b111111111;
assign micromatriz[80][17] = 9'b111111111;
assign micromatriz[80][18] = 9'b111111111;
assign micromatriz[80][19] = 9'b111111111;
assign micromatriz[80][20] = 9'b111111111;
assign micromatriz[80][21] = 9'b111111111;
assign micromatriz[80][22] = 9'b111111111;
assign micromatriz[80][23] = 9'b111111111;
assign micromatriz[80][24] = 9'b111111111;
assign micromatriz[80][25] = 9'b111111111;
assign micromatriz[80][26] = 9'b111111111;
assign micromatriz[80][27] = 9'b111111111;
assign micromatriz[80][28] = 9'b111111111;
assign micromatriz[80][29] = 9'b111111111;
assign micromatriz[80][30] = 9'b111111111;
assign micromatriz[80][31] = 9'b111111111;
assign micromatriz[80][32] = 9'b111111111;
assign micromatriz[80][33] = 9'b111111111;
assign micromatriz[80][34] = 9'b111111111;
assign micromatriz[80][35] = 9'b111111111;
assign micromatriz[80][36] = 9'b111111111;
assign micromatriz[80][37] = 9'b111111111;
assign micromatriz[80][38] = 9'b111111111;
assign micromatriz[80][39] = 9'b111111111;
assign micromatriz[80][40] = 9'b111111111;
assign micromatriz[80][41] = 9'b111111111;
assign micromatriz[80][42] = 9'b111111111;
assign micromatriz[80][43] = 9'b111111111;
assign micromatriz[80][44] = 9'b111111111;
assign micromatriz[80][45] = 9'b111111111;
assign micromatriz[80][46] = 9'b111111111;
assign micromatriz[80][47] = 9'b111111111;
assign micromatriz[80][48] = 9'b111111111;
assign micromatriz[80][49] = 9'b111111111;
assign micromatriz[80][50] = 9'b111111111;
assign micromatriz[80][51] = 9'b111111111;
assign micromatriz[80][52] = 9'b111111111;
assign micromatriz[80][53] = 9'b111111111;
assign micromatriz[80][54] = 9'b111111111;
assign micromatriz[80][55] = 9'b111111111;
assign micromatriz[80][56] = 9'b111111111;
assign micromatriz[80][57] = 9'b111111111;
assign micromatriz[80][58] = 9'b111111111;
assign micromatriz[80][59] = 9'b111111111;
assign micromatriz[80][60] = 9'b111111111;
assign micromatriz[80][61] = 9'b111111111;
assign micromatriz[80][62] = 9'b111111111;
assign micromatriz[80][63] = 9'b111111111;
assign micromatriz[80][64] = 9'b111111111;
assign micromatriz[80][65] = 9'b111111111;
assign micromatriz[80][66] = 9'b111111111;
assign micromatriz[80][67] = 9'b111111111;
assign micromatriz[80][68] = 9'b111111111;
assign micromatriz[80][69] = 9'b111111111;
assign micromatriz[80][70] = 9'b111111111;
assign micromatriz[80][71] = 9'b111111111;
assign micromatriz[80][72] = 9'b111111111;
assign micromatriz[80][73] = 9'b111111111;
assign micromatriz[80][74] = 9'b111111111;
assign micromatriz[80][75] = 9'b111111111;
assign micromatriz[80][76] = 9'b111111111;
assign micromatriz[80][77] = 9'b111111111;
assign micromatriz[80][78] = 9'b111111111;
assign micromatriz[80][79] = 9'b111111111;
assign micromatriz[80][80] = 9'b111111111;
assign micromatriz[80][81] = 9'b111111111;
assign micromatriz[80][82] = 9'b111111111;
assign micromatriz[80][83] = 9'b111111111;
assign micromatriz[80][84] = 9'b111111111;
assign micromatriz[80][85] = 9'b111111111;
assign micromatriz[80][86] = 9'b111111111;
assign micromatriz[80][87] = 9'b111111111;
assign micromatriz[80][88] = 9'b111111111;
assign micromatriz[80][89] = 9'b111111111;
assign micromatriz[80][90] = 9'b111111111;
assign micromatriz[80][91] = 9'b111111111;
assign micromatriz[80][92] = 9'b111111111;
assign micromatriz[80][93] = 9'b111111111;
assign micromatriz[80][94] = 9'b111111111;
assign micromatriz[80][95] = 9'b111111111;
assign micromatriz[80][96] = 9'b111111111;
assign micromatriz[80][97] = 9'b111111111;
assign micromatriz[80][98] = 9'b111111111;
assign micromatriz[80][99] = 9'b111111111;
assign micromatriz[81][0] = 9'b111111111;
assign micromatriz[81][1] = 9'b111111111;
assign micromatriz[81][2] = 9'b111111111;
assign micromatriz[81][3] = 9'b111111111;
assign micromatriz[81][4] = 9'b111111111;
assign micromatriz[81][5] = 9'b111111111;
assign micromatriz[81][6] = 9'b111111111;
assign micromatriz[81][7] = 9'b111111111;
assign micromatriz[81][8] = 9'b111111111;
assign micromatriz[81][9] = 9'b111111111;
assign micromatriz[81][10] = 9'b111111111;
assign micromatriz[81][11] = 9'b111111111;
assign micromatriz[81][12] = 9'b111111111;
assign micromatriz[81][13] = 9'b111111111;
assign micromatriz[81][14] = 9'b111111111;
assign micromatriz[81][15] = 9'b111111111;
assign micromatriz[81][16] = 9'b111111111;
assign micromatriz[81][17] = 9'b111111111;
assign micromatriz[81][18] = 9'b111111111;
assign micromatriz[81][19] = 9'b111111111;
assign micromatriz[81][20] = 9'b111111111;
assign micromatriz[81][21] = 9'b111111111;
assign micromatriz[81][22] = 9'b111111111;
assign micromatriz[81][23] = 9'b111111111;
assign micromatriz[81][24] = 9'b111111111;
assign micromatriz[81][25] = 9'b111111111;
assign micromatriz[81][26] = 9'b111111111;
assign micromatriz[81][27] = 9'b111111111;
assign micromatriz[81][28] = 9'b111111111;
assign micromatriz[81][29] = 9'b111111111;
assign micromatriz[81][30] = 9'b111111111;
assign micromatriz[81][31] = 9'b111111111;
assign micromatriz[81][32] = 9'b111111111;
assign micromatriz[81][33] = 9'b111111111;
assign micromatriz[81][34] = 9'b111111111;
assign micromatriz[81][35] = 9'b111111111;
assign micromatriz[81][36] = 9'b111111111;
assign micromatriz[81][37] = 9'b111111111;
assign micromatriz[81][38] = 9'b111111111;
assign micromatriz[81][39] = 9'b111111111;
assign micromatriz[81][40] = 9'b111111111;
assign micromatriz[81][41] = 9'b111111111;
assign micromatriz[81][42] = 9'b111111111;
assign micromatriz[81][43] = 9'b111111111;
assign micromatriz[81][44] = 9'b111111111;
assign micromatriz[81][45] = 9'b111111111;
assign micromatriz[81][46] = 9'b111111111;
assign micromatriz[81][47] = 9'b111111111;
assign micromatriz[81][48] = 9'b111111111;
assign micromatriz[81][49] = 9'b111111111;
assign micromatriz[81][50] = 9'b111111111;
assign micromatriz[81][51] = 9'b111111111;
assign micromatriz[81][52] = 9'b111111111;
assign micromatriz[81][53] = 9'b111111111;
assign micromatriz[81][54] = 9'b111111111;
assign micromatriz[81][55] = 9'b111111111;
assign micromatriz[81][56] = 9'b111111111;
assign micromatriz[81][57] = 9'b111111111;
assign micromatriz[81][58] = 9'b111111111;
assign micromatriz[81][59] = 9'b111111111;
assign micromatriz[81][60] = 9'b111111111;
assign micromatriz[81][61] = 9'b111111111;
assign micromatriz[81][62] = 9'b111111111;
assign micromatriz[81][63] = 9'b111111111;
assign micromatriz[81][64] = 9'b111111111;
assign micromatriz[81][65] = 9'b111111111;
assign micromatriz[81][66] = 9'b111111111;
assign micromatriz[81][67] = 9'b111111111;
assign micromatriz[81][68] = 9'b111111111;
assign micromatriz[81][69] = 9'b111111111;
assign micromatriz[81][70] = 9'b111111111;
assign micromatriz[81][71] = 9'b111111111;
assign micromatriz[81][72] = 9'b111111111;
assign micromatriz[81][73] = 9'b111111111;
assign micromatriz[81][74] = 9'b111111111;
assign micromatriz[81][75] = 9'b111111111;
assign micromatriz[81][76] = 9'b111111111;
assign micromatriz[81][77] = 9'b111111111;
assign micromatriz[81][78] = 9'b111111111;
assign micromatriz[81][79] = 9'b111111111;
assign micromatriz[81][80] = 9'b111111111;
assign micromatriz[81][81] = 9'b111111111;
assign micromatriz[81][82] = 9'b111111111;
assign micromatriz[81][83] = 9'b111111111;
assign micromatriz[81][84] = 9'b111111111;
assign micromatriz[81][85] = 9'b111111111;
assign micromatriz[81][86] = 9'b111111111;
assign micromatriz[81][87] = 9'b111111111;
assign micromatriz[81][88] = 9'b111111111;
assign micromatriz[81][89] = 9'b111111111;
assign micromatriz[81][90] = 9'b111111111;
assign micromatriz[81][91] = 9'b111111111;
assign micromatriz[81][92] = 9'b111111111;
assign micromatriz[81][93] = 9'b111111111;
assign micromatriz[81][94] = 9'b111111111;
assign micromatriz[81][95] = 9'b111111111;
assign micromatriz[81][96] = 9'b111111111;
assign micromatriz[81][97] = 9'b111111111;
assign micromatriz[81][98] = 9'b111111111;
assign micromatriz[81][99] = 9'b111111111;
assign micromatriz[82][0] = 9'b111111111;
assign micromatriz[82][1] = 9'b111111111;
assign micromatriz[82][2] = 9'b111111111;
assign micromatriz[82][3] = 9'b111111111;
assign micromatriz[82][4] = 9'b111111111;
assign micromatriz[82][5] = 9'b111111111;
assign micromatriz[82][6] = 9'b111111111;
assign micromatriz[82][7] = 9'b111111111;
assign micromatriz[82][8] = 9'b111111111;
assign micromatriz[82][9] = 9'b111111111;
assign micromatriz[82][10] = 9'b111111111;
assign micromatriz[82][11] = 9'b111111111;
assign micromatriz[82][12] = 9'b111111111;
assign micromatriz[82][13] = 9'b111111111;
assign micromatriz[82][14] = 9'b111111111;
assign micromatriz[82][15] = 9'b111111111;
assign micromatriz[82][16] = 9'b111111111;
assign micromatriz[82][17] = 9'b111111111;
assign micromatriz[82][18] = 9'b111111111;
assign micromatriz[82][19] = 9'b111111111;
assign micromatriz[82][20] = 9'b111111111;
assign micromatriz[82][21] = 9'b111111111;
assign micromatriz[82][22] = 9'b111111111;
assign micromatriz[82][23] = 9'b111111111;
assign micromatriz[82][24] = 9'b111111111;
assign micromatriz[82][25] = 9'b111111111;
assign micromatriz[82][26] = 9'b111111111;
assign micromatriz[82][27] = 9'b111111111;
assign micromatriz[82][28] = 9'b111111111;
assign micromatriz[82][29] = 9'b111111111;
assign micromatriz[82][30] = 9'b111111111;
assign micromatriz[82][31] = 9'b111111111;
assign micromatriz[82][32] = 9'b111111111;
assign micromatriz[82][33] = 9'b111111111;
assign micromatriz[82][34] = 9'b111111111;
assign micromatriz[82][35] = 9'b111111111;
assign micromatriz[82][36] = 9'b111111111;
assign micromatriz[82][37] = 9'b111111111;
assign micromatriz[82][38] = 9'b111111111;
assign micromatriz[82][39] = 9'b111111111;
assign micromatriz[82][40] = 9'b111111111;
assign micromatriz[82][41] = 9'b111111111;
assign micromatriz[82][42] = 9'b111111111;
assign micromatriz[82][43] = 9'b111111111;
assign micromatriz[82][44] = 9'b111111111;
assign micromatriz[82][45] = 9'b111111111;
assign micromatriz[82][46] = 9'b111111111;
assign micromatriz[82][47] = 9'b111111111;
assign micromatriz[82][48] = 9'b111111111;
assign micromatriz[82][49] = 9'b111111111;
assign micromatriz[82][50] = 9'b111111111;
assign micromatriz[82][51] = 9'b111111111;
assign micromatriz[82][52] = 9'b111111111;
assign micromatriz[82][53] = 9'b111111111;
assign micromatriz[82][54] = 9'b111111111;
assign micromatriz[82][55] = 9'b111111111;
assign micromatriz[82][56] = 9'b111111111;
assign micromatriz[82][57] = 9'b111111111;
assign micromatriz[82][58] = 9'b111111111;
assign micromatriz[82][59] = 9'b111111111;
assign micromatriz[82][60] = 9'b111111111;
assign micromatriz[82][61] = 9'b111111111;
assign micromatriz[82][62] = 9'b111111111;
assign micromatriz[82][63] = 9'b111111111;
assign micromatriz[82][64] = 9'b111111111;
assign micromatriz[82][65] = 9'b111111111;
assign micromatriz[82][66] = 9'b111111111;
assign micromatriz[82][67] = 9'b111111111;
assign micromatriz[82][68] = 9'b111111111;
assign micromatriz[82][69] = 9'b111111111;
assign micromatriz[82][70] = 9'b111111111;
assign micromatriz[82][71] = 9'b111111111;
assign micromatriz[82][72] = 9'b111111111;
assign micromatriz[82][73] = 9'b111111111;
assign micromatriz[82][74] = 9'b111111111;
assign micromatriz[82][75] = 9'b111111111;
assign micromatriz[82][76] = 9'b111111111;
assign micromatriz[82][77] = 9'b111111111;
assign micromatriz[82][78] = 9'b111111111;
assign micromatriz[82][79] = 9'b111111111;
assign micromatriz[82][80] = 9'b111111111;
assign micromatriz[82][81] = 9'b111111111;
assign micromatriz[82][82] = 9'b111111111;
assign micromatriz[82][83] = 9'b111111111;
assign micromatriz[82][84] = 9'b111111111;
assign micromatriz[82][85] = 9'b111111111;
assign micromatriz[82][86] = 9'b111111111;
assign micromatriz[82][87] = 9'b111111111;
assign micromatriz[82][88] = 9'b111111111;
assign micromatriz[82][89] = 9'b111111111;
assign micromatriz[82][90] = 9'b111111111;
assign micromatriz[82][91] = 9'b111111111;
assign micromatriz[82][92] = 9'b111111111;
assign micromatriz[82][93] = 9'b111111111;
assign micromatriz[82][94] = 9'b111111111;
assign micromatriz[82][95] = 9'b111111111;
assign micromatriz[82][96] = 9'b111111111;
assign micromatriz[82][97] = 9'b111111111;
assign micromatriz[82][98] = 9'b111111111;
assign micromatriz[82][99] = 9'b111111111;
assign micromatriz[83][0] = 9'b111111111;
assign micromatriz[83][1] = 9'b111111111;
assign micromatriz[83][2] = 9'b111111111;
assign micromatriz[83][3] = 9'b111111111;
assign micromatriz[83][4] = 9'b111111111;
assign micromatriz[83][5] = 9'b111111111;
assign micromatriz[83][6] = 9'b111111111;
assign micromatriz[83][7] = 9'b111111111;
assign micromatriz[83][8] = 9'b111111111;
assign micromatriz[83][9] = 9'b111111111;
assign micromatriz[83][10] = 9'b111111111;
assign micromatriz[83][11] = 9'b111111111;
assign micromatriz[83][12] = 9'b111111111;
assign micromatriz[83][13] = 9'b111111111;
assign micromatriz[83][14] = 9'b111111111;
assign micromatriz[83][15] = 9'b111111111;
assign micromatriz[83][16] = 9'b111111111;
assign micromatriz[83][17] = 9'b111111111;
assign micromatriz[83][18] = 9'b111111111;
assign micromatriz[83][19] = 9'b111111111;
assign micromatriz[83][20] = 9'b111111111;
assign micromatriz[83][21] = 9'b111111111;
assign micromatriz[83][22] = 9'b111111111;
assign micromatriz[83][23] = 9'b111111111;
assign micromatriz[83][24] = 9'b111111111;
assign micromatriz[83][25] = 9'b111111111;
assign micromatriz[83][26] = 9'b111111111;
assign micromatriz[83][27] = 9'b111111111;
assign micromatriz[83][28] = 9'b111111111;
assign micromatriz[83][29] = 9'b111111111;
assign micromatriz[83][30] = 9'b111111111;
assign micromatriz[83][31] = 9'b111111111;
assign micromatriz[83][32] = 9'b111111111;
assign micromatriz[83][33] = 9'b111111111;
assign micromatriz[83][34] = 9'b111111111;
assign micromatriz[83][35] = 9'b111111111;
assign micromatriz[83][36] = 9'b111111111;
assign micromatriz[83][37] = 9'b111111111;
assign micromatriz[83][38] = 9'b111111111;
assign micromatriz[83][39] = 9'b111111111;
assign micromatriz[83][40] = 9'b111111111;
assign micromatriz[83][41] = 9'b111111111;
assign micromatriz[83][42] = 9'b111111111;
assign micromatriz[83][43] = 9'b111111111;
assign micromatriz[83][44] = 9'b111111111;
assign micromatriz[83][45] = 9'b111111111;
assign micromatriz[83][46] = 9'b111111111;
assign micromatriz[83][47] = 9'b111111111;
assign micromatriz[83][48] = 9'b111111111;
assign micromatriz[83][49] = 9'b111111111;
assign micromatriz[83][50] = 9'b111111111;
assign micromatriz[83][51] = 9'b111111111;
assign micromatriz[83][52] = 9'b111111111;
assign micromatriz[83][53] = 9'b111111111;
assign micromatriz[83][54] = 9'b111111111;
assign micromatriz[83][55] = 9'b111111111;
assign micromatriz[83][56] = 9'b111111111;
assign micromatriz[83][57] = 9'b111111111;
assign micromatriz[83][58] = 9'b111111111;
assign micromatriz[83][59] = 9'b111111111;
assign micromatriz[83][60] = 9'b111111111;
assign micromatriz[83][61] = 9'b111111111;
assign micromatriz[83][62] = 9'b111111111;
assign micromatriz[83][63] = 9'b111111111;
assign micromatriz[83][64] = 9'b111111111;
assign micromatriz[83][65] = 9'b111111111;
assign micromatriz[83][66] = 9'b111111111;
assign micromatriz[83][67] = 9'b111111111;
assign micromatriz[83][68] = 9'b111111111;
assign micromatriz[83][69] = 9'b111111111;
assign micromatriz[83][70] = 9'b111111111;
assign micromatriz[83][71] = 9'b111111111;
assign micromatriz[83][72] = 9'b111111111;
assign micromatriz[83][73] = 9'b111111111;
assign micromatriz[83][74] = 9'b111111111;
assign micromatriz[83][75] = 9'b111111111;
assign micromatriz[83][76] = 9'b111111111;
assign micromatriz[83][77] = 9'b111111111;
assign micromatriz[83][78] = 9'b111111111;
assign micromatriz[83][79] = 9'b111111111;
assign micromatriz[83][80] = 9'b111111111;
assign micromatriz[83][81] = 9'b111111111;
assign micromatriz[83][82] = 9'b111111111;
assign micromatriz[83][83] = 9'b111111111;
assign micromatriz[83][84] = 9'b111111111;
assign micromatriz[83][85] = 9'b111111111;
assign micromatriz[83][86] = 9'b111111111;
assign micromatriz[83][87] = 9'b111111111;
assign micromatriz[83][88] = 9'b111111111;
assign micromatriz[83][89] = 9'b111111111;
assign micromatriz[83][90] = 9'b111111111;
assign micromatriz[83][91] = 9'b111111111;
assign micromatriz[83][92] = 9'b111111111;
assign micromatriz[83][93] = 9'b111111111;
assign micromatriz[83][94] = 9'b111111111;
assign micromatriz[83][95] = 9'b111111111;
assign micromatriz[83][96] = 9'b111111111;
assign micromatriz[83][97] = 9'b111111111;
assign micromatriz[83][98] = 9'b111111111;
assign micromatriz[83][99] = 9'b111111111;
assign micromatriz[84][0] = 9'b111111111;
assign micromatriz[84][1] = 9'b111111111;
assign micromatriz[84][2] = 9'b111111111;
assign micromatriz[84][3] = 9'b111111111;
assign micromatriz[84][4] = 9'b111111111;
assign micromatriz[84][5] = 9'b111111111;
assign micromatriz[84][6] = 9'b111111111;
assign micromatriz[84][7] = 9'b111111111;
assign micromatriz[84][8] = 9'b111111111;
assign micromatriz[84][9] = 9'b111111111;
assign micromatriz[84][10] = 9'b111111111;
assign micromatriz[84][11] = 9'b111111111;
assign micromatriz[84][12] = 9'b111111111;
assign micromatriz[84][13] = 9'b111111111;
assign micromatriz[84][14] = 9'b111111111;
assign micromatriz[84][15] = 9'b111111111;
assign micromatriz[84][16] = 9'b111111111;
assign micromatriz[84][17] = 9'b111111111;
assign micromatriz[84][18] = 9'b111111111;
assign micromatriz[84][19] = 9'b111111111;
assign micromatriz[84][20] = 9'b111111111;
assign micromatriz[84][21] = 9'b111111111;
assign micromatriz[84][22] = 9'b111111111;
assign micromatriz[84][23] = 9'b111111111;
assign micromatriz[84][24] = 9'b111111111;
assign micromatriz[84][25] = 9'b111111111;
assign micromatriz[84][26] = 9'b111111111;
assign micromatriz[84][27] = 9'b111111111;
assign micromatriz[84][28] = 9'b111111111;
assign micromatriz[84][29] = 9'b111111111;
assign micromatriz[84][30] = 9'b111111111;
assign micromatriz[84][31] = 9'b111111111;
assign micromatriz[84][32] = 9'b111111111;
assign micromatriz[84][33] = 9'b111111111;
assign micromatriz[84][34] = 9'b111111111;
assign micromatriz[84][35] = 9'b111111111;
assign micromatriz[84][36] = 9'b111111111;
assign micromatriz[84][37] = 9'b111111111;
assign micromatriz[84][38] = 9'b111111111;
assign micromatriz[84][39] = 9'b111111111;
assign micromatriz[84][40] = 9'b111111111;
assign micromatriz[84][41] = 9'b111111111;
assign micromatriz[84][42] = 9'b111111111;
assign micromatriz[84][43] = 9'b111111111;
assign micromatriz[84][44] = 9'b111111111;
assign micromatriz[84][45] = 9'b111111111;
assign micromatriz[84][46] = 9'b111111111;
assign micromatriz[84][47] = 9'b111111111;
assign micromatriz[84][48] = 9'b111111111;
assign micromatriz[84][49] = 9'b111111111;
assign micromatriz[84][50] = 9'b111111111;
assign micromatriz[84][51] = 9'b111111111;
assign micromatriz[84][52] = 9'b111111111;
assign micromatriz[84][53] = 9'b111111111;
assign micromatriz[84][54] = 9'b111111111;
assign micromatriz[84][55] = 9'b111111111;
assign micromatriz[84][56] = 9'b111111111;
assign micromatriz[84][57] = 9'b111111111;
assign micromatriz[84][58] = 9'b111111111;
assign micromatriz[84][59] = 9'b111111111;
assign micromatriz[84][60] = 9'b111111111;
assign micromatriz[84][61] = 9'b111111111;
assign micromatriz[84][62] = 9'b111111111;
assign micromatriz[84][63] = 9'b111111111;
assign micromatriz[84][64] = 9'b111111111;
assign micromatriz[84][65] = 9'b111111111;
assign micromatriz[84][66] = 9'b111111111;
assign micromatriz[84][67] = 9'b111111111;
assign micromatriz[84][68] = 9'b111111111;
assign micromatriz[84][69] = 9'b111111111;
assign micromatriz[84][70] = 9'b111111111;
assign micromatriz[84][71] = 9'b111111111;
assign micromatriz[84][72] = 9'b111111111;
assign micromatriz[84][73] = 9'b111111111;
assign micromatriz[84][74] = 9'b111111111;
assign micromatriz[84][75] = 9'b111111111;
assign micromatriz[84][76] = 9'b111111111;
assign micromatriz[84][77] = 9'b111111111;
assign micromatriz[84][78] = 9'b111111111;
assign micromatriz[84][79] = 9'b111111111;
assign micromatriz[84][80] = 9'b111111111;
assign micromatriz[84][81] = 9'b111111111;
assign micromatriz[84][82] = 9'b111111111;
assign micromatriz[84][83] = 9'b111111111;
assign micromatriz[84][84] = 9'b111111111;
assign micromatriz[84][85] = 9'b111111111;
assign micromatriz[84][86] = 9'b111111111;
assign micromatriz[84][87] = 9'b111111111;
assign micromatriz[84][88] = 9'b111111111;
assign micromatriz[84][89] = 9'b111111111;
assign micromatriz[84][90] = 9'b111111111;
assign micromatriz[84][91] = 9'b111111111;
assign micromatriz[84][92] = 9'b111111111;
assign micromatriz[84][93] = 9'b111111111;
assign micromatriz[84][94] = 9'b111111111;
assign micromatriz[84][95] = 9'b111111111;
assign micromatriz[84][96] = 9'b111111111;
assign micromatriz[84][97] = 9'b111111111;
assign micromatriz[84][98] = 9'b111111111;
assign micromatriz[84][99] = 9'b111111111;
assign micromatriz[85][0] = 9'b111111111;
assign micromatriz[85][1] = 9'b111111111;
assign micromatriz[85][2] = 9'b111111111;
assign micromatriz[85][3] = 9'b111111111;
assign micromatriz[85][4] = 9'b111111111;
assign micromatriz[85][5] = 9'b111111111;
assign micromatriz[85][6] = 9'b111111111;
assign micromatriz[85][7] = 9'b111111111;
assign micromatriz[85][8] = 9'b111111111;
assign micromatriz[85][9] = 9'b111111111;
assign micromatriz[85][10] = 9'b111111111;
assign micromatriz[85][11] = 9'b111111111;
assign micromatriz[85][12] = 9'b111111111;
assign micromatriz[85][13] = 9'b111111111;
assign micromatriz[85][14] = 9'b111111111;
assign micromatriz[85][15] = 9'b111111111;
assign micromatriz[85][16] = 9'b111111111;
assign micromatriz[85][17] = 9'b111111111;
assign micromatriz[85][18] = 9'b111111111;
assign micromatriz[85][19] = 9'b111111111;
assign micromatriz[85][20] = 9'b111111111;
assign micromatriz[85][21] = 9'b111111111;
assign micromatriz[85][22] = 9'b111111111;
assign micromatriz[85][23] = 9'b111111111;
assign micromatriz[85][24] = 9'b111111111;
assign micromatriz[85][25] = 9'b111111111;
assign micromatriz[85][26] = 9'b111111111;
assign micromatriz[85][27] = 9'b111111111;
assign micromatriz[85][28] = 9'b111111111;
assign micromatriz[85][29] = 9'b111111111;
assign micromatriz[85][30] = 9'b111111111;
assign micromatriz[85][31] = 9'b111111111;
assign micromatriz[85][32] = 9'b111111111;
assign micromatriz[85][33] = 9'b111111111;
assign micromatriz[85][34] = 9'b111111111;
assign micromatriz[85][35] = 9'b111111111;
assign micromatriz[85][36] = 9'b111111111;
assign micromatriz[85][37] = 9'b111111111;
assign micromatriz[85][38] = 9'b111111111;
assign micromatriz[85][39] = 9'b111111111;
assign micromatriz[85][40] = 9'b111111111;
assign micromatriz[85][41] = 9'b111111111;
assign micromatriz[85][42] = 9'b111111111;
assign micromatriz[85][43] = 9'b111111111;
assign micromatriz[85][44] = 9'b111111111;
assign micromatriz[85][45] = 9'b111111111;
assign micromatriz[85][46] = 9'b111111111;
assign micromatriz[85][47] = 9'b111111111;
assign micromatriz[85][48] = 9'b111111111;
assign micromatriz[85][49] = 9'b111111111;
assign micromatriz[85][50] = 9'b111111111;
assign micromatriz[85][51] = 9'b111111111;
assign micromatriz[85][52] = 9'b111111111;
assign micromatriz[85][53] = 9'b111111111;
assign micromatriz[85][54] = 9'b111111111;
assign micromatriz[85][55] = 9'b111111111;
assign micromatriz[85][56] = 9'b111111111;
assign micromatriz[85][57] = 9'b111111111;
assign micromatriz[85][58] = 9'b111111111;
assign micromatriz[85][59] = 9'b111111111;
assign micromatriz[85][60] = 9'b111111111;
assign micromatriz[85][61] = 9'b111111111;
assign micromatriz[85][62] = 9'b111111111;
assign micromatriz[85][63] = 9'b111111111;
assign micromatriz[85][64] = 9'b111111111;
assign micromatriz[85][65] = 9'b111111111;
assign micromatriz[85][66] = 9'b111111111;
assign micromatriz[85][67] = 9'b111111111;
assign micromatriz[85][68] = 9'b111111111;
assign micromatriz[85][69] = 9'b111111111;
assign micromatriz[85][70] = 9'b111111111;
assign micromatriz[85][71] = 9'b111111111;
assign micromatriz[85][72] = 9'b111111111;
assign micromatriz[85][73] = 9'b111111111;
assign micromatriz[85][74] = 9'b111111111;
assign micromatriz[85][75] = 9'b111111111;
assign micromatriz[85][76] = 9'b111111111;
assign micromatriz[85][77] = 9'b111111111;
assign micromatriz[85][78] = 9'b111111111;
assign micromatriz[85][79] = 9'b111111111;
assign micromatriz[85][80] = 9'b111111111;
assign micromatriz[85][81] = 9'b111111111;
assign micromatriz[85][82] = 9'b111111111;
assign micromatriz[85][83] = 9'b111111111;
assign micromatriz[85][84] = 9'b111111111;
assign micromatriz[85][85] = 9'b111111111;
assign micromatriz[85][86] = 9'b111111111;
assign micromatriz[85][87] = 9'b111111111;
assign micromatriz[85][88] = 9'b111111111;
assign micromatriz[85][89] = 9'b111111111;
assign micromatriz[85][90] = 9'b111111111;
assign micromatriz[85][91] = 9'b111111111;
assign micromatriz[85][92] = 9'b111111111;
assign micromatriz[85][93] = 9'b111111111;
assign micromatriz[85][94] = 9'b111111111;
assign micromatriz[85][95] = 9'b111111111;
assign micromatriz[85][96] = 9'b111111111;
assign micromatriz[85][97] = 9'b111111111;
assign micromatriz[85][98] = 9'b111111111;
assign micromatriz[85][99] = 9'b111111111;
assign micromatriz[86][0] = 9'b111111111;
assign micromatriz[86][1] = 9'b111111111;
assign micromatriz[86][2] = 9'b111111111;
assign micromatriz[86][3] = 9'b111111111;
assign micromatriz[86][4] = 9'b111111111;
assign micromatriz[86][5] = 9'b111111111;
assign micromatriz[86][6] = 9'b111111111;
assign micromatriz[86][7] = 9'b111111111;
assign micromatriz[86][8] = 9'b111111111;
assign micromatriz[86][9] = 9'b111111111;
assign micromatriz[86][10] = 9'b111111111;
assign micromatriz[86][11] = 9'b111111111;
assign micromatriz[86][12] = 9'b111111111;
assign micromatriz[86][13] = 9'b111111111;
assign micromatriz[86][14] = 9'b111111111;
assign micromatriz[86][15] = 9'b111111111;
assign micromatriz[86][16] = 9'b111111111;
assign micromatriz[86][17] = 9'b111111111;
assign micromatriz[86][18] = 9'b111111111;
assign micromatriz[86][19] = 9'b111111111;
assign micromatriz[86][20] = 9'b111111111;
assign micromatriz[86][21] = 9'b111111111;
assign micromatriz[86][22] = 9'b111111111;
assign micromatriz[86][23] = 9'b111111111;
assign micromatriz[86][24] = 9'b111111111;
assign micromatriz[86][25] = 9'b111111111;
assign micromatriz[86][26] = 9'b111111111;
assign micromatriz[86][27] = 9'b111111111;
assign micromatriz[86][28] = 9'b111111111;
assign micromatriz[86][29] = 9'b111111111;
assign micromatriz[86][30] = 9'b111111111;
assign micromatriz[86][31] = 9'b111111111;
assign micromatriz[86][32] = 9'b111111111;
assign micromatriz[86][33] = 9'b111111111;
assign micromatriz[86][34] = 9'b111111111;
assign micromatriz[86][35] = 9'b111111111;
assign micromatriz[86][36] = 9'b111111111;
assign micromatriz[86][37] = 9'b111111111;
assign micromatriz[86][38] = 9'b111111111;
assign micromatriz[86][39] = 9'b111111111;
assign micromatriz[86][40] = 9'b111111111;
assign micromatriz[86][41] = 9'b111111111;
assign micromatriz[86][42] = 9'b111111111;
assign micromatriz[86][43] = 9'b111111111;
assign micromatriz[86][44] = 9'b111111111;
assign micromatriz[86][45] = 9'b111111111;
assign micromatriz[86][46] = 9'b111111111;
assign micromatriz[86][47] = 9'b111111111;
assign micromatriz[86][48] = 9'b111111111;
assign micromatriz[86][49] = 9'b111111111;
assign micromatriz[86][50] = 9'b111111111;
assign micromatriz[86][51] = 9'b111111111;
assign micromatriz[86][52] = 9'b111111111;
assign micromatriz[86][53] = 9'b111111111;
assign micromatriz[86][54] = 9'b111111111;
assign micromatriz[86][55] = 9'b111111111;
assign micromatriz[86][56] = 9'b111111111;
assign micromatriz[86][57] = 9'b111111111;
assign micromatriz[86][58] = 9'b111111111;
assign micromatriz[86][59] = 9'b111111111;
assign micromatriz[86][60] = 9'b111111111;
assign micromatriz[86][61] = 9'b111111111;
assign micromatriz[86][62] = 9'b111111111;
assign micromatriz[86][63] = 9'b111111111;
assign micromatriz[86][64] = 9'b111111111;
assign micromatriz[86][65] = 9'b111111111;
assign micromatriz[86][66] = 9'b111111111;
assign micromatriz[86][67] = 9'b111111111;
assign micromatriz[86][68] = 9'b111111111;
assign micromatriz[86][69] = 9'b111111111;
assign micromatriz[86][70] = 9'b111111111;
assign micromatriz[86][71] = 9'b111111111;
assign micromatriz[86][72] = 9'b111111111;
assign micromatriz[86][73] = 9'b111111111;
assign micromatriz[86][74] = 9'b111111111;
assign micromatriz[86][75] = 9'b111111111;
assign micromatriz[86][76] = 9'b111111111;
assign micromatriz[86][77] = 9'b111111111;
assign micromatriz[86][78] = 9'b111111111;
assign micromatriz[86][79] = 9'b111111111;
assign micromatriz[86][80] = 9'b111111111;
assign micromatriz[86][81] = 9'b111111111;
assign micromatriz[86][82] = 9'b111111111;
assign micromatriz[86][83] = 9'b111111111;
assign micromatriz[86][84] = 9'b111111111;
assign micromatriz[86][85] = 9'b111111111;
assign micromatriz[86][86] = 9'b111111111;
assign micromatriz[86][87] = 9'b111111111;
assign micromatriz[86][88] = 9'b111111111;
assign micromatriz[86][89] = 9'b111111111;
assign micromatriz[86][90] = 9'b111111111;
assign micromatriz[86][91] = 9'b111111111;
assign micromatriz[86][92] = 9'b111111111;
assign micromatriz[86][93] = 9'b111111111;
assign micromatriz[86][94] = 9'b111111111;
assign micromatriz[86][95] = 9'b111111111;
assign micromatriz[86][96] = 9'b111111111;
assign micromatriz[86][97] = 9'b111111111;
assign micromatriz[86][98] = 9'b111111111;
assign micromatriz[86][99] = 9'b111111111;
assign micromatriz[87][0] = 9'b111111111;
assign micromatriz[87][1] = 9'b111111111;
assign micromatriz[87][2] = 9'b111111111;
assign micromatriz[87][3] = 9'b111111111;
assign micromatriz[87][4] = 9'b111111111;
assign micromatriz[87][5] = 9'b111111111;
assign micromatriz[87][6] = 9'b111111111;
assign micromatriz[87][7] = 9'b111111111;
assign micromatriz[87][8] = 9'b111111111;
assign micromatriz[87][9] = 9'b111111111;
assign micromatriz[87][10] = 9'b111111111;
assign micromatriz[87][11] = 9'b111111111;
assign micromatriz[87][12] = 9'b111111111;
assign micromatriz[87][13] = 9'b111111111;
assign micromatriz[87][14] = 9'b111111111;
assign micromatriz[87][15] = 9'b111111111;
assign micromatriz[87][16] = 9'b111111111;
assign micromatriz[87][17] = 9'b111111111;
assign micromatriz[87][18] = 9'b111111111;
assign micromatriz[87][19] = 9'b111111111;
assign micromatriz[87][20] = 9'b111111111;
assign micromatriz[87][21] = 9'b111111111;
assign micromatriz[87][22] = 9'b111111111;
assign micromatriz[87][23] = 9'b111111111;
assign micromatriz[87][24] = 9'b111111111;
assign micromatriz[87][25] = 9'b111111111;
assign micromatriz[87][26] = 9'b111111111;
assign micromatriz[87][27] = 9'b111111111;
assign micromatriz[87][28] = 9'b111111111;
assign micromatriz[87][29] = 9'b111111111;
assign micromatriz[87][30] = 9'b111111111;
assign micromatriz[87][31] = 9'b111111111;
assign micromatriz[87][32] = 9'b111111111;
assign micromatriz[87][33] = 9'b111111111;
assign micromatriz[87][34] = 9'b111111111;
assign micromatriz[87][35] = 9'b111111111;
assign micromatriz[87][36] = 9'b111111111;
assign micromatriz[87][37] = 9'b111111111;
assign micromatriz[87][38] = 9'b111111111;
assign micromatriz[87][39] = 9'b111111111;
assign micromatriz[87][40] = 9'b111111111;
assign micromatriz[87][41] = 9'b111111111;
assign micromatriz[87][42] = 9'b111111111;
assign micromatriz[87][43] = 9'b111111111;
assign micromatriz[87][44] = 9'b111111111;
assign micromatriz[87][45] = 9'b111111111;
assign micromatriz[87][46] = 9'b111111111;
assign micromatriz[87][47] = 9'b111111111;
assign micromatriz[87][48] = 9'b111111111;
assign micromatriz[87][49] = 9'b111111111;
assign micromatriz[87][50] = 9'b111111111;
assign micromatriz[87][51] = 9'b111111111;
assign micromatriz[87][52] = 9'b111111111;
assign micromatriz[87][53] = 9'b111111111;
assign micromatriz[87][54] = 9'b111111111;
assign micromatriz[87][55] = 9'b111111111;
assign micromatriz[87][56] = 9'b111111111;
assign micromatriz[87][57] = 9'b111111111;
assign micromatriz[87][58] = 9'b111111111;
assign micromatriz[87][59] = 9'b111111111;
assign micromatriz[87][60] = 9'b111111111;
assign micromatriz[87][61] = 9'b111111111;
assign micromatriz[87][62] = 9'b111111111;
assign micromatriz[87][63] = 9'b111111111;
assign micromatriz[87][64] = 9'b111111111;
assign micromatriz[87][65] = 9'b111111111;
assign micromatriz[87][66] = 9'b111111111;
assign micromatriz[87][67] = 9'b111111111;
assign micromatriz[87][68] = 9'b111111111;
assign micromatriz[87][69] = 9'b111111111;
assign micromatriz[87][70] = 9'b111111111;
assign micromatriz[87][71] = 9'b111111111;
assign micromatriz[87][72] = 9'b111111111;
assign micromatriz[87][73] = 9'b111111111;
assign micromatriz[87][74] = 9'b111111111;
assign micromatriz[87][75] = 9'b111111111;
assign micromatriz[87][76] = 9'b111111111;
assign micromatriz[87][77] = 9'b111111111;
assign micromatriz[87][78] = 9'b111111111;
assign micromatriz[87][79] = 9'b111111111;
assign micromatriz[87][80] = 9'b111111111;
assign micromatriz[87][81] = 9'b111111111;
assign micromatriz[87][82] = 9'b111111111;
assign micromatriz[87][83] = 9'b111111111;
assign micromatriz[87][84] = 9'b111111111;
assign micromatriz[87][85] = 9'b111111111;
assign micromatriz[87][86] = 9'b111111111;
assign micromatriz[87][87] = 9'b111111111;
assign micromatriz[87][88] = 9'b111111111;
assign micromatriz[87][89] = 9'b111111111;
assign micromatriz[87][90] = 9'b111111111;
assign micromatriz[87][91] = 9'b111111111;
assign micromatriz[87][92] = 9'b111111111;
assign micromatriz[87][93] = 9'b111111111;
assign micromatriz[87][94] = 9'b111111111;
assign micromatriz[87][95] = 9'b111111111;
assign micromatriz[87][96] = 9'b111111111;
assign micromatriz[87][97] = 9'b111111111;
assign micromatriz[87][98] = 9'b111111111;
assign micromatriz[87][99] = 9'b111111111;
assign micromatriz[88][0] = 9'b111111111;
assign micromatriz[88][1] = 9'b111111111;
assign micromatriz[88][2] = 9'b111111111;
assign micromatriz[88][3] = 9'b111111111;
assign micromatriz[88][4] = 9'b111111111;
assign micromatriz[88][5] = 9'b111111111;
assign micromatriz[88][6] = 9'b111111111;
assign micromatriz[88][7] = 9'b111111111;
assign micromatriz[88][8] = 9'b111111111;
assign micromatriz[88][9] = 9'b111111111;
assign micromatriz[88][10] = 9'b111111111;
assign micromatriz[88][11] = 9'b111111111;
assign micromatriz[88][12] = 9'b111111111;
assign micromatriz[88][13] = 9'b111111111;
assign micromatriz[88][14] = 9'b111111111;
assign micromatriz[88][15] = 9'b111111111;
assign micromatriz[88][16] = 9'b111111111;
assign micromatriz[88][17] = 9'b111111111;
assign micromatriz[88][18] = 9'b111111111;
assign micromatriz[88][19] = 9'b111111111;
assign micromatriz[88][20] = 9'b111111111;
assign micromatriz[88][21] = 9'b111111111;
assign micromatriz[88][22] = 9'b111111111;
assign micromatriz[88][23] = 9'b111111111;
assign micromatriz[88][24] = 9'b111111111;
assign micromatriz[88][25] = 9'b111111111;
assign micromatriz[88][26] = 9'b111111111;
assign micromatriz[88][27] = 9'b111111111;
assign micromatriz[88][28] = 9'b111111111;
assign micromatriz[88][29] = 9'b111111111;
assign micromatriz[88][30] = 9'b111111111;
assign micromatriz[88][31] = 9'b111111111;
assign micromatriz[88][32] = 9'b111111111;
assign micromatriz[88][33] = 9'b111111111;
assign micromatriz[88][34] = 9'b111111111;
assign micromatriz[88][35] = 9'b111111111;
assign micromatriz[88][36] = 9'b111111111;
assign micromatriz[88][37] = 9'b111111111;
assign micromatriz[88][38] = 9'b111111111;
assign micromatriz[88][39] = 9'b111111111;
assign micromatriz[88][40] = 9'b111111111;
assign micromatriz[88][41] = 9'b111111111;
assign micromatriz[88][42] = 9'b111111111;
assign micromatriz[88][43] = 9'b111111111;
assign micromatriz[88][44] = 9'b111111111;
assign micromatriz[88][45] = 9'b111111111;
assign micromatriz[88][46] = 9'b111111111;
assign micromatriz[88][47] = 9'b111111111;
assign micromatriz[88][48] = 9'b111111111;
assign micromatriz[88][49] = 9'b111111111;
assign micromatriz[88][50] = 9'b111111111;
assign micromatriz[88][51] = 9'b111111111;
assign micromatriz[88][52] = 9'b111111111;
assign micromatriz[88][53] = 9'b111111111;
assign micromatriz[88][54] = 9'b111111111;
assign micromatriz[88][55] = 9'b111111111;
assign micromatriz[88][56] = 9'b111111111;
assign micromatriz[88][57] = 9'b111111111;
assign micromatriz[88][58] = 9'b111111111;
assign micromatriz[88][59] = 9'b111111111;
assign micromatriz[88][60] = 9'b111111111;
assign micromatriz[88][61] = 9'b111111111;
assign micromatriz[88][62] = 9'b111111111;
assign micromatriz[88][63] = 9'b111111111;
assign micromatriz[88][64] = 9'b111111111;
assign micromatriz[88][65] = 9'b111111111;
assign micromatriz[88][66] = 9'b111111111;
assign micromatriz[88][67] = 9'b111111111;
assign micromatriz[88][68] = 9'b111111111;
assign micromatriz[88][69] = 9'b111111111;
assign micromatriz[88][70] = 9'b111111111;
assign micromatriz[88][71] = 9'b111111111;
assign micromatriz[88][72] = 9'b111111111;
assign micromatriz[88][73] = 9'b111111111;
assign micromatriz[88][74] = 9'b111111111;
assign micromatriz[88][75] = 9'b111111111;
assign micromatriz[88][76] = 9'b111111111;
assign micromatriz[88][77] = 9'b111111111;
assign micromatriz[88][78] = 9'b111111111;
assign micromatriz[88][79] = 9'b111111111;
assign micromatriz[88][80] = 9'b111111111;
assign micromatriz[88][81] = 9'b111111111;
assign micromatriz[88][82] = 9'b111111111;
assign micromatriz[88][83] = 9'b111111111;
assign micromatriz[88][84] = 9'b111111111;
assign micromatriz[88][85] = 9'b111111111;
assign micromatriz[88][86] = 9'b111111111;
assign micromatriz[88][87] = 9'b111111111;
assign micromatriz[88][88] = 9'b111111111;
assign micromatriz[88][89] = 9'b111111111;
assign micromatriz[88][90] = 9'b111111111;
assign micromatriz[88][91] = 9'b111111111;
assign micromatriz[88][92] = 9'b111111111;
assign micromatriz[88][93] = 9'b111111111;
assign micromatriz[88][94] = 9'b111111111;
assign micromatriz[88][95] = 9'b111111111;
assign micromatriz[88][96] = 9'b111111111;
assign micromatriz[88][97] = 9'b111111111;
assign micromatriz[88][98] = 9'b111111111;
assign micromatriz[88][99] = 9'b111111111;
assign micromatriz[89][0] = 9'b111111111;
assign micromatriz[89][1] = 9'b111111111;
assign micromatriz[89][2] = 9'b111111111;
assign micromatriz[89][3] = 9'b111111111;
assign micromatriz[89][4] = 9'b111111111;
assign micromatriz[89][5] = 9'b111111111;
assign micromatriz[89][6] = 9'b111111111;
assign micromatriz[89][7] = 9'b111111111;
assign micromatriz[89][8] = 9'b111111111;
assign micromatriz[89][9] = 9'b111111111;
assign micromatriz[89][10] = 9'b111111111;
assign micromatriz[89][11] = 9'b111111111;
assign micromatriz[89][12] = 9'b111111111;
assign micromatriz[89][13] = 9'b111111111;
assign micromatriz[89][14] = 9'b111111111;
assign micromatriz[89][15] = 9'b111111111;
assign micromatriz[89][16] = 9'b111111111;
assign micromatriz[89][17] = 9'b111111111;
assign micromatriz[89][18] = 9'b111111111;
assign micromatriz[89][19] = 9'b111111111;
assign micromatriz[89][20] = 9'b111111111;
assign micromatriz[89][21] = 9'b111111111;
assign micromatriz[89][22] = 9'b111111111;
assign micromatriz[89][23] = 9'b111111111;
assign micromatriz[89][24] = 9'b111111111;
assign micromatriz[89][25] = 9'b111111111;
assign micromatriz[89][26] = 9'b111111111;
assign micromatriz[89][27] = 9'b111111111;
assign micromatriz[89][28] = 9'b111111111;
assign micromatriz[89][29] = 9'b111111111;
assign micromatriz[89][30] = 9'b111111111;
assign micromatriz[89][31] = 9'b111111111;
assign micromatriz[89][32] = 9'b111111111;
assign micromatriz[89][33] = 9'b111111111;
assign micromatriz[89][34] = 9'b111111111;
assign micromatriz[89][35] = 9'b111111111;
assign micromatriz[89][36] = 9'b111111111;
assign micromatriz[89][37] = 9'b111111111;
assign micromatriz[89][38] = 9'b111111111;
assign micromatriz[89][39] = 9'b111111111;
assign micromatriz[89][40] = 9'b111111111;
assign micromatriz[89][41] = 9'b111111111;
assign micromatriz[89][42] = 9'b111111111;
assign micromatriz[89][43] = 9'b111111111;
assign micromatriz[89][44] = 9'b111111111;
assign micromatriz[89][45] = 9'b111111111;
assign micromatriz[89][46] = 9'b111111111;
assign micromatriz[89][47] = 9'b111111111;
assign micromatriz[89][48] = 9'b111111111;
assign micromatriz[89][49] = 9'b111111111;
assign micromatriz[89][50] = 9'b111111111;
assign micromatriz[89][51] = 9'b111111111;
assign micromatriz[89][52] = 9'b111111111;
assign micromatriz[89][53] = 9'b111111111;
assign micromatriz[89][54] = 9'b111111111;
assign micromatriz[89][55] = 9'b111111111;
assign micromatriz[89][56] = 9'b111111111;
assign micromatriz[89][57] = 9'b111111111;
assign micromatriz[89][58] = 9'b111111111;
assign micromatriz[89][59] = 9'b111111111;
assign micromatriz[89][60] = 9'b111111111;
assign micromatriz[89][61] = 9'b111111111;
assign micromatriz[89][62] = 9'b111111111;
assign micromatriz[89][63] = 9'b111111111;
assign micromatriz[89][64] = 9'b111111111;
assign micromatriz[89][65] = 9'b111111111;
assign micromatriz[89][66] = 9'b111111111;
assign micromatriz[89][67] = 9'b111111111;
assign micromatriz[89][68] = 9'b111111111;
assign micromatriz[89][69] = 9'b111111111;
assign micromatriz[89][70] = 9'b111111111;
assign micromatriz[89][71] = 9'b111111111;
assign micromatriz[89][72] = 9'b111111111;
assign micromatriz[89][73] = 9'b111111111;
assign micromatriz[89][74] = 9'b111111111;
assign micromatriz[89][75] = 9'b111111111;
assign micromatriz[89][76] = 9'b111111111;
assign micromatriz[89][77] = 9'b111111111;
assign micromatriz[89][78] = 9'b111111111;
assign micromatriz[89][79] = 9'b111111111;
assign micromatriz[89][80] = 9'b111111111;
assign micromatriz[89][81] = 9'b111111111;
assign micromatriz[89][82] = 9'b111111111;
assign micromatriz[89][83] = 9'b111111111;
assign micromatriz[89][84] = 9'b111111111;
assign micromatriz[89][85] = 9'b111111111;
assign micromatriz[89][86] = 9'b111111111;
assign micromatriz[89][87] = 9'b111111111;
assign micromatriz[89][88] = 9'b111111111;
assign micromatriz[89][89] = 9'b111111111;
assign micromatriz[89][90] = 9'b111111111;
assign micromatriz[89][91] = 9'b111111111;
assign micromatriz[89][92] = 9'b111111111;
assign micromatriz[89][93] = 9'b111111111;
assign micromatriz[89][94] = 9'b111111111;
assign micromatriz[89][95] = 9'b111111111;
assign micromatriz[89][96] = 9'b111111111;
assign micromatriz[89][97] = 9'b111111111;
assign micromatriz[89][98] = 9'b111111111;
assign micromatriz[89][99] = 9'b111111111;
assign micromatriz[90][0] = 9'b111111111;
assign micromatriz[90][1] = 9'b111111111;
assign micromatriz[90][2] = 9'b111111111;
assign micromatriz[90][3] = 9'b111111111;
assign micromatriz[90][4] = 9'b111111111;
assign micromatriz[90][5] = 9'b111111111;
assign micromatriz[90][6] = 9'b111111111;
assign micromatriz[90][7] = 9'b111111111;
assign micromatriz[90][8] = 9'b111111111;
assign micromatriz[90][9] = 9'b111111111;
assign micromatriz[90][10] = 9'b111111111;
assign micromatriz[90][11] = 9'b111111111;
assign micromatriz[90][12] = 9'b111111111;
assign micromatriz[90][13] = 9'b111111111;
assign micromatriz[90][14] = 9'b111111111;
assign micromatriz[90][15] = 9'b111111111;
assign micromatriz[90][16] = 9'b111111111;
assign micromatriz[90][17] = 9'b111111111;
assign micromatriz[90][18] = 9'b111111111;
assign micromatriz[90][19] = 9'b111111111;
assign micromatriz[90][20] = 9'b111111111;
assign micromatriz[90][21] = 9'b111111111;
assign micromatriz[90][22] = 9'b111111111;
assign micromatriz[90][23] = 9'b111111111;
assign micromatriz[90][24] = 9'b111111111;
assign micromatriz[90][25] = 9'b111111111;
assign micromatriz[90][26] = 9'b111111111;
assign micromatriz[90][27] = 9'b111111111;
assign micromatriz[90][28] = 9'b111111111;
assign micromatriz[90][29] = 9'b111111111;
assign micromatriz[90][30] = 9'b111111111;
assign micromatriz[90][31] = 9'b111111111;
assign micromatriz[90][32] = 9'b111111111;
assign micromatriz[90][33] = 9'b111111111;
assign micromatriz[90][34] = 9'b111111111;
assign micromatriz[90][35] = 9'b111111111;
assign micromatriz[90][36] = 9'b111111111;
assign micromatriz[90][37] = 9'b111111111;
assign micromatriz[90][38] = 9'b111111111;
assign micromatriz[90][39] = 9'b111111111;
assign micromatriz[90][40] = 9'b111111111;
assign micromatriz[90][41] = 9'b111111111;
assign micromatriz[90][42] = 9'b111111111;
assign micromatriz[90][43] = 9'b111111111;
assign micromatriz[90][44] = 9'b111111111;
assign micromatriz[90][45] = 9'b111111111;
assign micromatriz[90][46] = 9'b111111111;
assign micromatriz[90][47] = 9'b111111111;
assign micromatriz[90][48] = 9'b111111111;
assign micromatriz[90][49] = 9'b111111111;
assign micromatriz[90][50] = 9'b111111111;
assign micromatriz[90][51] = 9'b111111111;
assign micromatriz[90][52] = 9'b111111111;
assign micromatriz[90][53] = 9'b111111111;
assign micromatriz[90][54] = 9'b111111111;
assign micromatriz[90][55] = 9'b111111111;
assign micromatriz[90][56] = 9'b111111111;
assign micromatriz[90][57] = 9'b111111111;
assign micromatriz[90][58] = 9'b111111111;
assign micromatriz[90][59] = 9'b111111111;
assign micromatriz[90][60] = 9'b111111111;
assign micromatriz[90][61] = 9'b111111111;
assign micromatriz[90][62] = 9'b111111111;
assign micromatriz[90][63] = 9'b111111111;
assign micromatriz[90][64] = 9'b111111111;
assign micromatriz[90][65] = 9'b111111111;
assign micromatriz[90][66] = 9'b111111111;
assign micromatriz[90][67] = 9'b111111111;
assign micromatriz[90][68] = 9'b111111111;
assign micromatriz[90][69] = 9'b111111111;
assign micromatriz[90][70] = 9'b111111111;
assign micromatriz[90][71] = 9'b111111111;
assign micromatriz[90][72] = 9'b111111111;
assign micromatriz[90][73] = 9'b111111111;
assign micromatriz[90][74] = 9'b111111111;
assign micromatriz[90][75] = 9'b111111111;
assign micromatriz[90][76] = 9'b111111111;
assign micromatriz[90][77] = 9'b111111111;
assign micromatriz[90][78] = 9'b111111111;
assign micromatriz[90][79] = 9'b111111111;
assign micromatriz[90][80] = 9'b111111111;
assign micromatriz[90][81] = 9'b111111111;
assign micromatriz[90][82] = 9'b111111111;
assign micromatriz[90][83] = 9'b111111111;
assign micromatriz[90][84] = 9'b111111111;
assign micromatriz[90][85] = 9'b111111111;
assign micromatriz[90][86] = 9'b111111111;
assign micromatriz[90][87] = 9'b111111111;
assign micromatriz[90][88] = 9'b111111111;
assign micromatriz[90][89] = 9'b111111111;
assign micromatriz[90][90] = 9'b111111111;
assign micromatriz[90][91] = 9'b111111111;
assign micromatriz[90][92] = 9'b111111111;
assign micromatriz[90][93] = 9'b111111111;
assign micromatriz[90][94] = 9'b111111111;
assign micromatriz[90][95] = 9'b111111111;
assign micromatriz[90][96] = 9'b111111111;
assign micromatriz[90][97] = 9'b111111111;
assign micromatriz[90][98] = 9'b111111111;
assign micromatriz[90][99] = 9'b111111111;
assign micromatriz[91][0] = 9'b111111111;
assign micromatriz[91][1] = 9'b111111111;
assign micromatriz[91][2] = 9'b111111111;
assign micromatriz[91][3] = 9'b111111111;
assign micromatriz[91][4] = 9'b111111111;
assign micromatriz[91][5] = 9'b111111111;
assign micromatriz[91][6] = 9'b111111111;
assign micromatriz[91][7] = 9'b111111111;
assign micromatriz[91][8] = 9'b111111111;
assign micromatriz[91][9] = 9'b111111111;
assign micromatriz[91][10] = 9'b111111111;
assign micromatriz[91][11] = 9'b111111111;
assign micromatriz[91][12] = 9'b111111111;
assign micromatriz[91][13] = 9'b111111111;
assign micromatriz[91][14] = 9'b111111111;
assign micromatriz[91][15] = 9'b111111111;
assign micromatriz[91][16] = 9'b111111111;
assign micromatriz[91][17] = 9'b111111111;
assign micromatriz[91][18] = 9'b111111111;
assign micromatriz[91][19] = 9'b111111111;
assign micromatriz[91][20] = 9'b111111111;
assign micromatriz[91][21] = 9'b111111111;
assign micromatriz[91][22] = 9'b111111111;
assign micromatriz[91][23] = 9'b111111111;
assign micromatriz[91][24] = 9'b111111111;
assign micromatriz[91][25] = 9'b111111111;
assign micromatriz[91][26] = 9'b111111111;
assign micromatriz[91][27] = 9'b111111111;
assign micromatriz[91][28] = 9'b111111111;
assign micromatriz[91][29] = 9'b111111111;
assign micromatriz[91][30] = 9'b111111111;
assign micromatriz[91][31] = 9'b111111111;
assign micromatriz[91][32] = 9'b111111111;
assign micromatriz[91][33] = 9'b111111111;
assign micromatriz[91][34] = 9'b111111111;
assign micromatriz[91][35] = 9'b111111111;
assign micromatriz[91][36] = 9'b111111111;
assign micromatriz[91][37] = 9'b111111111;
assign micromatriz[91][38] = 9'b111111111;
assign micromatriz[91][39] = 9'b111111111;
assign micromatriz[91][40] = 9'b111111111;
assign micromatriz[91][41] = 9'b111111111;
assign micromatriz[91][42] = 9'b111111111;
assign micromatriz[91][43] = 9'b111111111;
assign micromatriz[91][44] = 9'b111111111;
assign micromatriz[91][45] = 9'b111111111;
assign micromatriz[91][46] = 9'b111111111;
assign micromatriz[91][47] = 9'b111111111;
assign micromatriz[91][48] = 9'b111111111;
assign micromatriz[91][49] = 9'b111111111;
assign micromatriz[91][50] = 9'b111111111;
assign micromatriz[91][51] = 9'b111111111;
assign micromatriz[91][52] = 9'b111111111;
assign micromatriz[91][53] = 9'b111111111;
assign micromatriz[91][54] = 9'b111111111;
assign micromatriz[91][55] = 9'b111111111;
assign micromatriz[91][56] = 9'b111111111;
assign micromatriz[91][57] = 9'b111111111;
assign micromatriz[91][58] = 9'b111111111;
assign micromatriz[91][59] = 9'b111111111;
assign micromatriz[91][60] = 9'b111111111;
assign micromatriz[91][61] = 9'b111111111;
assign micromatriz[91][62] = 9'b111111111;
assign micromatriz[91][63] = 9'b111111111;
assign micromatriz[91][64] = 9'b111111111;
assign micromatriz[91][65] = 9'b111111111;
assign micromatriz[91][66] = 9'b111111111;
assign micromatriz[91][67] = 9'b111111111;
assign micromatriz[91][68] = 9'b111111111;
assign micromatriz[91][69] = 9'b111111111;
assign micromatriz[91][70] = 9'b111111111;
assign micromatriz[91][71] = 9'b111111111;
assign micromatriz[91][72] = 9'b111111111;
assign micromatriz[91][73] = 9'b111111111;
assign micromatriz[91][74] = 9'b111111111;
assign micromatriz[91][75] = 9'b111111111;
assign micromatriz[91][76] = 9'b111111111;
assign micromatriz[91][77] = 9'b111111111;
assign micromatriz[91][78] = 9'b111111111;
assign micromatriz[91][79] = 9'b111111111;
assign micromatriz[91][80] = 9'b111111111;
assign micromatriz[91][81] = 9'b111111111;
assign micromatriz[91][82] = 9'b111111111;
assign micromatriz[91][83] = 9'b111111111;
assign micromatriz[91][84] = 9'b111111111;
assign micromatriz[91][85] = 9'b111111111;
assign micromatriz[91][86] = 9'b111111111;
assign micromatriz[91][87] = 9'b111111111;
assign micromatriz[91][88] = 9'b111111111;
assign micromatriz[91][89] = 9'b111111111;
assign micromatriz[91][90] = 9'b111111111;
assign micromatriz[91][91] = 9'b111111111;
assign micromatriz[91][92] = 9'b111111111;
assign micromatriz[91][93] = 9'b111111111;
assign micromatriz[91][94] = 9'b111111111;
assign micromatriz[91][95] = 9'b111111111;
assign micromatriz[91][96] = 9'b111111111;
assign micromatriz[91][97] = 9'b111111111;
assign micromatriz[91][98] = 9'b111111111;
assign micromatriz[91][99] = 9'b111111111;
assign micromatriz[92][0] = 9'b111111111;
assign micromatriz[92][1] = 9'b111111111;
assign micromatriz[92][2] = 9'b111111111;
assign micromatriz[92][3] = 9'b111111111;
assign micromatriz[92][4] = 9'b111111111;
assign micromatriz[92][5] = 9'b111111111;
assign micromatriz[92][6] = 9'b111111111;
assign micromatriz[92][7] = 9'b111111111;
assign micromatriz[92][8] = 9'b111111111;
assign micromatriz[92][9] = 9'b111111111;
assign micromatriz[92][10] = 9'b111111111;
assign micromatriz[92][11] = 9'b111111111;
assign micromatriz[92][12] = 9'b111111111;
assign micromatriz[92][13] = 9'b111111111;
assign micromatriz[92][14] = 9'b111111111;
assign micromatriz[92][15] = 9'b111111111;
assign micromatriz[92][16] = 9'b111111111;
assign micromatriz[92][17] = 9'b111111111;
assign micromatriz[92][18] = 9'b111111111;
assign micromatriz[92][19] = 9'b111111111;
assign micromatriz[92][20] = 9'b111111111;
assign micromatriz[92][21] = 9'b111111111;
assign micromatriz[92][22] = 9'b111111111;
assign micromatriz[92][23] = 9'b111111111;
assign micromatriz[92][24] = 9'b111111111;
assign micromatriz[92][25] = 9'b111111111;
assign micromatriz[92][26] = 9'b111111111;
assign micromatriz[92][27] = 9'b111111111;
assign micromatriz[92][28] = 9'b111111111;
assign micromatriz[92][29] = 9'b111111111;
assign micromatriz[92][30] = 9'b111111111;
assign micromatriz[92][31] = 9'b111111111;
assign micromatriz[92][32] = 9'b111111111;
assign micromatriz[92][33] = 9'b111111111;
assign micromatriz[92][34] = 9'b111111111;
assign micromatriz[92][35] = 9'b111111111;
assign micromatriz[92][36] = 9'b111111111;
assign micromatriz[92][37] = 9'b111111111;
assign micromatriz[92][38] = 9'b111111111;
assign micromatriz[92][39] = 9'b111111111;
assign micromatriz[92][40] = 9'b111111111;
assign micromatriz[92][41] = 9'b111111111;
assign micromatriz[92][42] = 9'b111111111;
assign micromatriz[92][43] = 9'b111111111;
assign micromatriz[92][44] = 9'b111111111;
assign micromatriz[92][45] = 9'b111111111;
assign micromatriz[92][46] = 9'b111111111;
assign micromatriz[92][47] = 9'b111111111;
assign micromatriz[92][48] = 9'b111111111;
assign micromatriz[92][49] = 9'b111111111;
assign micromatriz[92][50] = 9'b111111111;
assign micromatriz[92][51] = 9'b111111111;
assign micromatriz[92][52] = 9'b111111111;
assign micromatriz[92][53] = 9'b111111111;
assign micromatriz[92][54] = 9'b111111111;
assign micromatriz[92][55] = 9'b111111111;
assign micromatriz[92][56] = 9'b111111111;
assign micromatriz[92][57] = 9'b111111111;
assign micromatriz[92][58] = 9'b111111111;
assign micromatriz[92][59] = 9'b111111111;
assign micromatriz[92][60] = 9'b111111111;
assign micromatriz[92][61] = 9'b111111111;
assign micromatriz[92][62] = 9'b111111111;
assign micromatriz[92][63] = 9'b111111111;
assign micromatriz[92][64] = 9'b111111111;
assign micromatriz[92][65] = 9'b111111111;
assign micromatriz[92][66] = 9'b111111111;
assign micromatriz[92][67] = 9'b111111111;
assign micromatriz[92][68] = 9'b111111111;
assign micromatriz[92][69] = 9'b111111111;
assign micromatriz[92][70] = 9'b111111111;
assign micromatriz[92][71] = 9'b111111111;
assign micromatriz[92][72] = 9'b111111111;
assign micromatriz[92][73] = 9'b111111111;
assign micromatriz[92][74] = 9'b111111111;
assign micromatriz[92][75] = 9'b111111111;
assign micromatriz[92][76] = 9'b111111111;
assign micromatriz[92][77] = 9'b111111111;
assign micromatriz[92][78] = 9'b111111111;
assign micromatriz[92][79] = 9'b111111111;
assign micromatriz[92][80] = 9'b111111111;
assign micromatriz[92][81] = 9'b111111111;
assign micromatriz[92][82] = 9'b111111111;
assign micromatriz[92][83] = 9'b111111111;
assign micromatriz[92][84] = 9'b111111111;
assign micromatriz[92][85] = 9'b111111111;
assign micromatriz[92][86] = 9'b111111111;
assign micromatriz[92][87] = 9'b111111111;
assign micromatriz[92][88] = 9'b111111111;
assign micromatriz[92][89] = 9'b111111111;
assign micromatriz[92][90] = 9'b111111111;
assign micromatriz[92][91] = 9'b111111111;
assign micromatriz[92][92] = 9'b111111111;
assign micromatriz[92][93] = 9'b111111111;
assign micromatriz[92][94] = 9'b111111111;
assign micromatriz[92][95] = 9'b111111111;
assign micromatriz[92][96] = 9'b111111111;
assign micromatriz[92][97] = 9'b111111111;
assign micromatriz[92][98] = 9'b111111111;
assign micromatriz[92][99] = 9'b111111111;
assign micromatriz[93][0] = 9'b111111111;
assign micromatriz[93][1] = 9'b111111111;
assign micromatriz[93][2] = 9'b111111111;
assign micromatriz[93][3] = 9'b111111111;
assign micromatriz[93][4] = 9'b111111111;
assign micromatriz[93][5] = 9'b111111111;
assign micromatriz[93][6] = 9'b111111111;
assign micromatriz[93][7] = 9'b111111111;
assign micromatriz[93][8] = 9'b111111111;
assign micromatriz[93][9] = 9'b111111111;
assign micromatriz[93][10] = 9'b111111111;
assign micromatriz[93][11] = 9'b111111111;
assign micromatriz[93][12] = 9'b111111111;
assign micromatriz[93][13] = 9'b111111111;
assign micromatriz[93][14] = 9'b111111111;
assign micromatriz[93][15] = 9'b111111111;
assign micromatriz[93][16] = 9'b111111111;
assign micromatriz[93][17] = 9'b111111111;
assign micromatriz[93][18] = 9'b111111111;
assign micromatriz[93][19] = 9'b111111111;
assign micromatriz[93][20] = 9'b111111111;
assign micromatriz[93][21] = 9'b111111111;
assign micromatriz[93][22] = 9'b111111111;
assign micromatriz[93][23] = 9'b111111111;
assign micromatriz[93][24] = 9'b111111111;
assign micromatriz[93][25] = 9'b111111111;
assign micromatriz[93][26] = 9'b111111111;
assign micromatriz[93][27] = 9'b111111111;
assign micromatriz[93][28] = 9'b111111111;
assign micromatriz[93][29] = 9'b111111111;
assign micromatriz[93][30] = 9'b111111111;
assign micromatriz[93][31] = 9'b111111111;
assign micromatriz[93][32] = 9'b111111111;
assign micromatriz[93][33] = 9'b111111111;
assign micromatriz[93][34] = 9'b111111111;
assign micromatriz[93][35] = 9'b111111111;
assign micromatriz[93][36] = 9'b111111111;
assign micromatriz[93][37] = 9'b111111111;
assign micromatriz[93][38] = 9'b111111111;
assign micromatriz[93][39] = 9'b111111111;
assign micromatriz[93][40] = 9'b111111111;
assign micromatriz[93][41] = 9'b111111111;
assign micromatriz[93][42] = 9'b111111111;
assign micromatriz[93][43] = 9'b111111111;
assign micromatriz[93][44] = 9'b111111111;
assign micromatriz[93][45] = 9'b111111111;
assign micromatriz[93][46] = 9'b111111111;
assign micromatriz[93][47] = 9'b111111111;
assign micromatriz[93][48] = 9'b111111111;
assign micromatriz[93][49] = 9'b111111111;
assign micromatriz[93][50] = 9'b111111111;
assign micromatriz[93][51] = 9'b111111111;
assign micromatriz[93][52] = 9'b111111111;
assign micromatriz[93][53] = 9'b111111111;
assign micromatriz[93][54] = 9'b111111111;
assign micromatriz[93][55] = 9'b111111111;
assign micromatriz[93][56] = 9'b111111111;
assign micromatriz[93][57] = 9'b111111111;
assign micromatriz[93][58] = 9'b111111111;
assign micromatriz[93][59] = 9'b111111111;
assign micromatriz[93][60] = 9'b111111111;
assign micromatriz[93][61] = 9'b111111111;
assign micromatriz[93][62] = 9'b111111111;
assign micromatriz[93][63] = 9'b111111111;
assign micromatriz[93][64] = 9'b111111111;
assign micromatriz[93][65] = 9'b111111111;
assign micromatriz[93][66] = 9'b111111111;
assign micromatriz[93][67] = 9'b111111111;
assign micromatriz[93][68] = 9'b111111111;
assign micromatriz[93][69] = 9'b111111111;
assign micromatriz[93][70] = 9'b111111111;
assign micromatriz[93][71] = 9'b111111111;
assign micromatriz[93][72] = 9'b111111111;
assign micromatriz[93][73] = 9'b111111111;
assign micromatriz[93][74] = 9'b111111111;
assign micromatriz[93][75] = 9'b111111111;
assign micromatriz[93][76] = 9'b111111111;
assign micromatriz[93][77] = 9'b111111111;
assign micromatriz[93][78] = 9'b111111111;
assign micromatriz[93][79] = 9'b111111111;
assign micromatriz[93][80] = 9'b111111111;
assign micromatriz[93][81] = 9'b111111111;
assign micromatriz[93][82] = 9'b111111111;
assign micromatriz[93][83] = 9'b111111111;
assign micromatriz[93][84] = 9'b111111111;
assign micromatriz[93][85] = 9'b111111111;
assign micromatriz[93][86] = 9'b111111111;
assign micromatriz[93][87] = 9'b111111111;
assign micromatriz[93][88] = 9'b111111111;
assign micromatriz[93][89] = 9'b111111111;
assign micromatriz[93][90] = 9'b111111111;
assign micromatriz[93][91] = 9'b111111111;
assign micromatriz[93][92] = 9'b111111111;
assign micromatriz[93][93] = 9'b111111111;
assign micromatriz[93][94] = 9'b111111111;
assign micromatriz[93][95] = 9'b111111111;
assign micromatriz[93][96] = 9'b111111111;
assign micromatriz[93][97] = 9'b111111111;
assign micromatriz[93][98] = 9'b111111111;
assign micromatriz[93][99] = 9'b111111111;
assign micromatriz[94][0] = 9'b111111111;
assign micromatriz[94][1] = 9'b111111111;
assign micromatriz[94][2] = 9'b111111111;
assign micromatriz[94][3] = 9'b111111111;
assign micromatriz[94][4] = 9'b111111111;
assign micromatriz[94][5] = 9'b111111111;
assign micromatriz[94][6] = 9'b111111111;
assign micromatriz[94][7] = 9'b111111111;
assign micromatriz[94][8] = 9'b111111111;
assign micromatriz[94][9] = 9'b111111111;
assign micromatriz[94][10] = 9'b111111111;
assign micromatriz[94][11] = 9'b111111111;
assign micromatriz[94][12] = 9'b111111111;
assign micromatriz[94][13] = 9'b111111111;
assign micromatriz[94][14] = 9'b111111111;
assign micromatriz[94][15] = 9'b111111111;
assign micromatriz[94][16] = 9'b111111111;
assign micromatriz[94][17] = 9'b111111111;
assign micromatriz[94][18] = 9'b111111111;
assign micromatriz[94][19] = 9'b111111111;
assign micromatriz[94][20] = 9'b111111111;
assign micromatriz[94][21] = 9'b111111111;
assign micromatriz[94][22] = 9'b111111111;
assign micromatriz[94][23] = 9'b111111111;
assign micromatriz[94][24] = 9'b111111111;
assign micromatriz[94][25] = 9'b111111111;
assign micromatriz[94][26] = 9'b111111111;
assign micromatriz[94][27] = 9'b111111111;
assign micromatriz[94][28] = 9'b111111111;
assign micromatriz[94][29] = 9'b111111111;
assign micromatriz[94][30] = 9'b111111111;
assign micromatriz[94][31] = 9'b111111111;
assign micromatriz[94][32] = 9'b111111111;
assign micromatriz[94][33] = 9'b111111111;
assign micromatriz[94][34] = 9'b111111111;
assign micromatriz[94][35] = 9'b111111111;
assign micromatriz[94][36] = 9'b111111111;
assign micromatriz[94][37] = 9'b111111111;
assign micromatriz[94][38] = 9'b111111111;
assign micromatriz[94][39] = 9'b111111111;
assign micromatriz[94][40] = 9'b111111111;
assign micromatriz[94][41] = 9'b111111111;
assign micromatriz[94][42] = 9'b111111111;
assign micromatriz[94][43] = 9'b111111111;
assign micromatriz[94][44] = 9'b111111111;
assign micromatriz[94][45] = 9'b111111111;
assign micromatriz[94][46] = 9'b111111111;
assign micromatriz[94][47] = 9'b111111111;
assign micromatriz[94][48] = 9'b111111111;
assign micromatriz[94][49] = 9'b111111111;
assign micromatriz[94][50] = 9'b111111111;
assign micromatriz[94][51] = 9'b111111111;
assign micromatriz[94][52] = 9'b111111111;
assign micromatriz[94][53] = 9'b111111111;
assign micromatriz[94][54] = 9'b111111111;
assign micromatriz[94][55] = 9'b111111111;
assign micromatriz[94][56] = 9'b111111111;
assign micromatriz[94][57] = 9'b111111111;
assign micromatriz[94][58] = 9'b111111111;
assign micromatriz[94][59] = 9'b111111111;
assign micromatriz[94][60] = 9'b111111111;
assign micromatriz[94][61] = 9'b111111111;
assign micromatriz[94][62] = 9'b111111111;
assign micromatriz[94][63] = 9'b111111111;
assign micromatriz[94][64] = 9'b111111111;
assign micromatriz[94][65] = 9'b111111111;
assign micromatriz[94][66] = 9'b111111111;
assign micromatriz[94][67] = 9'b111111111;
assign micromatriz[94][68] = 9'b111111111;
assign micromatriz[94][69] = 9'b111111111;
assign micromatriz[94][70] = 9'b111111111;
assign micromatriz[94][71] = 9'b111111111;
assign micromatriz[94][72] = 9'b111111111;
assign micromatriz[94][73] = 9'b111111111;
assign micromatriz[94][74] = 9'b111111111;
assign micromatriz[94][75] = 9'b111111111;
assign micromatriz[94][76] = 9'b111111111;
assign micromatriz[94][77] = 9'b111111111;
assign micromatriz[94][78] = 9'b111111111;
assign micromatriz[94][79] = 9'b111111111;
assign micromatriz[94][80] = 9'b111111111;
assign micromatriz[94][81] = 9'b111111111;
assign micromatriz[94][82] = 9'b111111111;
assign micromatriz[94][83] = 9'b111111111;
assign micromatriz[94][84] = 9'b111111111;
assign micromatriz[94][85] = 9'b111111111;
assign micromatriz[94][86] = 9'b111111111;
assign micromatriz[94][87] = 9'b111111111;
assign micromatriz[94][88] = 9'b111111111;
assign micromatriz[94][89] = 9'b111111111;
assign micromatriz[94][90] = 9'b111111111;
assign micromatriz[94][91] = 9'b111111111;
assign micromatriz[94][92] = 9'b111111111;
assign micromatriz[94][93] = 9'b111111111;
assign micromatriz[94][94] = 9'b111111111;
assign micromatriz[94][95] = 9'b111111111;
assign micromatriz[94][96] = 9'b111111111;
assign micromatriz[94][97] = 9'b111111111;
assign micromatriz[94][98] = 9'b111111111;
assign micromatriz[94][99] = 9'b111111111;
assign micromatriz[95][0] = 9'b111111111;
assign micromatriz[95][1] = 9'b111111111;
assign micromatriz[95][2] = 9'b111111111;
assign micromatriz[95][3] = 9'b111111111;
assign micromatriz[95][4] = 9'b111111111;
assign micromatriz[95][5] = 9'b111111111;
assign micromatriz[95][6] = 9'b111111111;
assign micromatriz[95][7] = 9'b111111111;
assign micromatriz[95][8] = 9'b111111111;
assign micromatriz[95][9] = 9'b111111111;
assign micromatriz[95][10] = 9'b111111111;
assign micromatriz[95][11] = 9'b111111111;
assign micromatriz[95][12] = 9'b111111111;
assign micromatriz[95][13] = 9'b111111111;
assign micromatriz[95][14] = 9'b111111111;
assign micromatriz[95][15] = 9'b111111111;
assign micromatriz[95][16] = 9'b111111111;
assign micromatriz[95][17] = 9'b111111111;
assign micromatriz[95][18] = 9'b111111111;
assign micromatriz[95][19] = 9'b111111111;
assign micromatriz[95][20] = 9'b111111111;
assign micromatriz[95][21] = 9'b111111111;
assign micromatriz[95][22] = 9'b111111111;
assign micromatriz[95][23] = 9'b111111111;
assign micromatriz[95][24] = 9'b111111111;
assign micromatriz[95][25] = 9'b111111111;
assign micromatriz[95][26] = 9'b111111111;
assign micromatriz[95][27] = 9'b111111111;
assign micromatriz[95][28] = 9'b111111111;
assign micromatriz[95][29] = 9'b111111111;
assign micromatriz[95][30] = 9'b111111111;
assign micromatriz[95][31] = 9'b111111111;
assign micromatriz[95][32] = 9'b111111111;
assign micromatriz[95][33] = 9'b111111111;
assign micromatriz[95][34] = 9'b111111111;
assign micromatriz[95][35] = 9'b111111111;
assign micromatriz[95][36] = 9'b111111111;
assign micromatriz[95][37] = 9'b111111111;
assign micromatriz[95][38] = 9'b111111111;
assign micromatriz[95][39] = 9'b111111111;
assign micromatriz[95][40] = 9'b111111111;
assign micromatriz[95][41] = 9'b111111111;
assign micromatriz[95][42] = 9'b111111111;
assign micromatriz[95][43] = 9'b111111111;
assign micromatriz[95][44] = 9'b111111111;
assign micromatriz[95][45] = 9'b111111111;
assign micromatriz[95][46] = 9'b111111111;
assign micromatriz[95][47] = 9'b111111111;
assign micromatriz[95][48] = 9'b111111111;
assign micromatriz[95][49] = 9'b111111111;
assign micromatriz[95][50] = 9'b111111111;
assign micromatriz[95][51] = 9'b111111111;
assign micromatriz[95][52] = 9'b111111111;
assign micromatriz[95][53] = 9'b111111111;
assign micromatriz[95][54] = 9'b111111111;
assign micromatriz[95][55] = 9'b111111111;
assign micromatriz[95][56] = 9'b111111111;
assign micromatriz[95][57] = 9'b111111111;
assign micromatriz[95][58] = 9'b111111111;
assign micromatriz[95][59] = 9'b111111111;
assign micromatriz[95][60] = 9'b111111111;
assign micromatriz[95][61] = 9'b111111111;
assign micromatriz[95][62] = 9'b111111111;
assign micromatriz[95][63] = 9'b111111111;
assign micromatriz[95][64] = 9'b111111111;
assign micromatriz[95][65] = 9'b111111111;
assign micromatriz[95][66] = 9'b111111111;
assign micromatriz[95][67] = 9'b111111111;
assign micromatriz[95][68] = 9'b111111111;
assign micromatriz[95][69] = 9'b111111111;
assign micromatriz[95][70] = 9'b111111111;
assign micromatriz[95][71] = 9'b111111111;
assign micromatriz[95][72] = 9'b111111111;
assign micromatriz[95][73] = 9'b111111111;
assign micromatriz[95][74] = 9'b111111111;
assign micromatriz[95][75] = 9'b111111111;
assign micromatriz[95][76] = 9'b111111111;
assign micromatriz[95][77] = 9'b111111111;
assign micromatriz[95][78] = 9'b111111111;
assign micromatriz[95][79] = 9'b111111111;
assign micromatriz[95][80] = 9'b111111111;
assign micromatriz[95][81] = 9'b111111111;
assign micromatriz[95][82] = 9'b111111111;
assign micromatriz[95][83] = 9'b111111111;
assign micromatriz[95][84] = 9'b111111111;
assign micromatriz[95][85] = 9'b111111111;
assign micromatriz[95][86] = 9'b111111111;
assign micromatriz[95][87] = 9'b111111111;
assign micromatriz[95][88] = 9'b111111111;
assign micromatriz[95][89] = 9'b111111111;
assign micromatriz[95][90] = 9'b111111111;
assign micromatriz[95][91] = 9'b111111111;
assign micromatriz[95][92] = 9'b111111111;
assign micromatriz[95][93] = 9'b111111111;
assign micromatriz[95][94] = 9'b111111111;
assign micromatriz[95][95] = 9'b111111111;
assign micromatriz[95][96] = 9'b111111111;
assign micromatriz[95][97] = 9'b111111111;
assign micromatriz[95][98] = 9'b111111111;
assign micromatriz[95][99] = 9'b111111111;
assign micromatriz[96][0] = 9'b111111111;
assign micromatriz[96][1] = 9'b111111111;
assign micromatriz[96][2] = 9'b111111111;
assign micromatriz[96][3] = 9'b111111111;
assign micromatriz[96][4] = 9'b111111111;
assign micromatriz[96][5] = 9'b111111111;
assign micromatriz[96][6] = 9'b111111111;
assign micromatriz[96][7] = 9'b111111111;
assign micromatriz[96][8] = 9'b111111111;
assign micromatriz[96][9] = 9'b111111111;
assign micromatriz[96][10] = 9'b111111111;
assign micromatriz[96][11] = 9'b111111111;
assign micromatriz[96][12] = 9'b111111111;
assign micromatriz[96][13] = 9'b111111111;
assign micromatriz[96][14] = 9'b111111111;
assign micromatriz[96][15] = 9'b111111111;
assign micromatriz[96][16] = 9'b111111111;
assign micromatriz[96][17] = 9'b111111111;
assign micromatriz[96][18] = 9'b111111111;
assign micromatriz[96][19] = 9'b111111111;
assign micromatriz[96][20] = 9'b111111111;
assign micromatriz[96][21] = 9'b111111111;
assign micromatriz[96][22] = 9'b111111111;
assign micromatriz[96][23] = 9'b111111111;
assign micromatriz[96][24] = 9'b111111111;
assign micromatriz[96][25] = 9'b111111111;
assign micromatriz[96][26] = 9'b111111111;
assign micromatriz[96][27] = 9'b111111111;
assign micromatriz[96][28] = 9'b111111111;
assign micromatriz[96][29] = 9'b111111111;
assign micromatriz[96][30] = 9'b111111111;
assign micromatriz[96][31] = 9'b111111111;
assign micromatriz[96][32] = 9'b111111111;
assign micromatriz[96][33] = 9'b111111111;
assign micromatriz[96][34] = 9'b111111111;
assign micromatriz[96][35] = 9'b111111111;
assign micromatriz[96][36] = 9'b111111111;
assign micromatriz[96][37] = 9'b111111111;
assign micromatriz[96][38] = 9'b111111111;
assign micromatriz[96][39] = 9'b111111111;
assign micromatriz[96][40] = 9'b111111111;
assign micromatriz[96][41] = 9'b111111111;
assign micromatriz[96][42] = 9'b111111111;
assign micromatriz[96][43] = 9'b111111111;
assign micromatriz[96][44] = 9'b111111111;
assign micromatriz[96][45] = 9'b111111111;
assign micromatriz[96][46] = 9'b111111111;
assign micromatriz[96][47] = 9'b111111111;
assign micromatriz[96][48] = 9'b111111111;
assign micromatriz[96][49] = 9'b111111111;
assign micromatriz[96][50] = 9'b111111111;
assign micromatriz[96][51] = 9'b111111111;
assign micromatriz[96][52] = 9'b111111111;
assign micromatriz[96][53] = 9'b111111111;
assign micromatriz[96][54] = 9'b111111111;
assign micromatriz[96][55] = 9'b111111111;
assign micromatriz[96][56] = 9'b111111111;
assign micromatriz[96][57] = 9'b111111111;
assign micromatriz[96][58] = 9'b111111111;
assign micromatriz[96][59] = 9'b111111111;
assign micromatriz[96][60] = 9'b111111111;
assign micromatriz[96][61] = 9'b111111111;
assign micromatriz[96][62] = 9'b111111111;
assign micromatriz[96][63] = 9'b111111111;
assign micromatriz[96][64] = 9'b111111111;
assign micromatriz[96][65] = 9'b111111111;
assign micromatriz[96][66] = 9'b111111111;
assign micromatriz[96][67] = 9'b111111111;
assign micromatriz[96][68] = 9'b111111111;
assign micromatriz[96][69] = 9'b111111111;
assign micromatriz[96][70] = 9'b111111111;
assign micromatriz[96][71] = 9'b111111111;
assign micromatriz[96][72] = 9'b111111111;
assign micromatriz[96][73] = 9'b111111111;
assign micromatriz[96][74] = 9'b111111111;
assign micromatriz[96][75] = 9'b111111111;
assign micromatriz[96][76] = 9'b111111111;
assign micromatriz[96][77] = 9'b111111111;
assign micromatriz[96][78] = 9'b111111111;
assign micromatriz[96][79] = 9'b111111111;
assign micromatriz[96][80] = 9'b111111111;
assign micromatriz[96][81] = 9'b111111111;
assign micromatriz[96][82] = 9'b111111111;
assign micromatriz[96][83] = 9'b111111111;
assign micromatriz[96][84] = 9'b111111111;
assign micromatriz[96][85] = 9'b111111111;
assign micromatriz[96][86] = 9'b111111111;
assign micromatriz[96][87] = 9'b111111111;
assign micromatriz[96][88] = 9'b111111111;
assign micromatriz[96][89] = 9'b111111111;
assign micromatriz[96][90] = 9'b111111111;
assign micromatriz[96][91] = 9'b111111111;
assign micromatriz[96][92] = 9'b111111111;
assign micromatriz[96][93] = 9'b111111111;
assign micromatriz[96][94] = 9'b111111111;
assign micromatriz[96][95] = 9'b111111111;
assign micromatriz[96][96] = 9'b111111111;
assign micromatriz[96][97] = 9'b111111111;
assign micromatriz[96][98] = 9'b111111111;
assign micromatriz[96][99] = 9'b111111111;
assign micromatriz[97][0] = 9'b111111111;
assign micromatriz[97][1] = 9'b111111111;
assign micromatriz[97][2] = 9'b111111111;
assign micromatriz[97][3] = 9'b111111111;
assign micromatriz[97][4] = 9'b111111111;
assign micromatriz[97][5] = 9'b111111111;
assign micromatriz[97][6] = 9'b111111111;
assign micromatriz[97][7] = 9'b111111111;
assign micromatriz[97][8] = 9'b111111111;
assign micromatriz[97][9] = 9'b111111111;
assign micromatriz[97][10] = 9'b111111111;
assign micromatriz[97][11] = 9'b111111111;
assign micromatriz[97][12] = 9'b111111111;
assign micromatriz[97][13] = 9'b111111111;
assign micromatriz[97][14] = 9'b111111111;
assign micromatriz[97][15] = 9'b111111111;
assign micromatriz[97][16] = 9'b111111111;
assign micromatriz[97][17] = 9'b111111111;
assign micromatriz[97][18] = 9'b111111111;
assign micromatriz[97][19] = 9'b111111111;
assign micromatriz[97][20] = 9'b111111111;
assign micromatriz[97][21] = 9'b111111111;
assign micromatriz[97][22] = 9'b111111111;
assign micromatriz[97][23] = 9'b111111111;
assign micromatriz[97][24] = 9'b111111111;
assign micromatriz[97][25] = 9'b111111111;
assign micromatriz[97][26] = 9'b111111111;
assign micromatriz[97][27] = 9'b111111111;
assign micromatriz[97][28] = 9'b111111111;
assign micromatriz[97][29] = 9'b111111111;
assign micromatriz[97][30] = 9'b111111111;
assign micromatriz[97][31] = 9'b111111111;
assign micromatriz[97][32] = 9'b111111111;
assign micromatriz[97][33] = 9'b111111111;
assign micromatriz[97][34] = 9'b111111111;
assign micromatriz[97][35] = 9'b111111111;
assign micromatriz[97][36] = 9'b111111111;
assign micromatriz[97][37] = 9'b111111111;
assign micromatriz[97][38] = 9'b111111111;
assign micromatriz[97][39] = 9'b111111111;
assign micromatriz[97][40] = 9'b111111111;
assign micromatriz[97][41] = 9'b111111111;
assign micromatriz[97][42] = 9'b111111111;
assign micromatriz[97][43] = 9'b111111111;
assign micromatriz[97][44] = 9'b111111111;
assign micromatriz[97][45] = 9'b111111111;
assign micromatriz[97][46] = 9'b111111111;
assign micromatriz[97][47] = 9'b111111111;
assign micromatriz[97][48] = 9'b111111111;
assign micromatriz[97][49] = 9'b111111111;
assign micromatriz[97][50] = 9'b111111111;
assign micromatriz[97][51] = 9'b111111111;
assign micromatriz[97][52] = 9'b111111111;
assign micromatriz[97][53] = 9'b111111111;
assign micromatriz[97][54] = 9'b111111111;
assign micromatriz[97][55] = 9'b111111111;
assign micromatriz[97][56] = 9'b111111111;
assign micromatriz[97][57] = 9'b111111111;
assign micromatriz[97][58] = 9'b111111111;
assign micromatriz[97][59] = 9'b111111111;
assign micromatriz[97][60] = 9'b111111111;
assign micromatriz[97][61] = 9'b111111111;
assign micromatriz[97][62] = 9'b111111111;
assign micromatriz[97][63] = 9'b111111111;
assign micromatriz[97][64] = 9'b111111111;
assign micromatriz[97][65] = 9'b111111111;
assign micromatriz[97][66] = 9'b111111111;
assign micromatriz[97][67] = 9'b111111111;
assign micromatriz[97][68] = 9'b111111111;
assign micromatriz[97][69] = 9'b111111111;
assign micromatriz[97][70] = 9'b111111111;
assign micromatriz[97][71] = 9'b111111111;
assign micromatriz[97][72] = 9'b111111111;
assign micromatriz[97][73] = 9'b111111111;
assign micromatriz[97][74] = 9'b111111111;
assign micromatriz[97][75] = 9'b111111111;
assign micromatriz[97][76] = 9'b111111111;
assign micromatriz[97][77] = 9'b111111111;
assign micromatriz[97][78] = 9'b111111111;
assign micromatriz[97][79] = 9'b111111111;
assign micromatriz[97][80] = 9'b111111111;
assign micromatriz[97][81] = 9'b111111111;
assign micromatriz[97][82] = 9'b111111111;
assign micromatriz[97][83] = 9'b111111111;
assign micromatriz[97][84] = 9'b111111111;
assign micromatriz[97][85] = 9'b111111111;
assign micromatriz[97][86] = 9'b111111111;
assign micromatriz[97][87] = 9'b111111111;
assign micromatriz[97][88] = 9'b111111111;
assign micromatriz[97][89] = 9'b111111111;
assign micromatriz[97][90] = 9'b111111111;
assign micromatriz[97][91] = 9'b111111111;
assign micromatriz[97][92] = 9'b111111111;
assign micromatriz[97][93] = 9'b111111111;
assign micromatriz[97][94] = 9'b111111111;
assign micromatriz[97][95] = 9'b111111111;
assign micromatriz[97][96] = 9'b111111111;
assign micromatriz[97][97] = 9'b111111111;
assign micromatriz[97][98] = 9'b111111111;
assign micromatriz[97][99] = 9'b111111111;
assign micromatriz[98][0] = 9'b111111111;
assign micromatriz[98][1] = 9'b111111111;
assign micromatriz[98][2] = 9'b111111111;
assign micromatriz[98][3] = 9'b111111111;
assign micromatriz[98][4] = 9'b111111111;
assign micromatriz[98][5] = 9'b111111111;
assign micromatriz[98][6] = 9'b111111111;
assign micromatriz[98][7] = 9'b111111111;
assign micromatriz[98][8] = 9'b111111111;
assign micromatriz[98][9] = 9'b111111111;
assign micromatriz[98][10] = 9'b111111111;
assign micromatriz[98][11] = 9'b111111111;
assign micromatriz[98][12] = 9'b111111111;
assign micromatriz[98][13] = 9'b111111111;
assign micromatriz[98][14] = 9'b111111111;
assign micromatriz[98][15] = 9'b111111111;
assign micromatriz[98][16] = 9'b111111111;
assign micromatriz[98][17] = 9'b111111111;
assign micromatriz[98][18] = 9'b111111111;
assign micromatriz[98][19] = 9'b111111111;
assign micromatriz[98][20] = 9'b111111111;
assign micromatriz[98][21] = 9'b111111111;
assign micromatriz[98][22] = 9'b111111111;
assign micromatriz[98][23] = 9'b111111111;
assign micromatriz[98][24] = 9'b111111111;
assign micromatriz[98][25] = 9'b111111111;
assign micromatriz[98][26] = 9'b111111111;
assign micromatriz[98][27] = 9'b111111111;
assign micromatriz[98][28] = 9'b111111111;
assign micromatriz[98][29] = 9'b111111111;
assign micromatriz[98][30] = 9'b111111111;
assign micromatriz[98][31] = 9'b111111111;
assign micromatriz[98][32] = 9'b111111111;
assign micromatriz[98][33] = 9'b111111111;
assign micromatriz[98][34] = 9'b111111111;
assign micromatriz[98][35] = 9'b111111111;
assign micromatriz[98][36] = 9'b111111111;
assign micromatriz[98][37] = 9'b111111111;
assign micromatriz[98][38] = 9'b111111111;
assign micromatriz[98][39] = 9'b111111111;
assign micromatriz[98][40] = 9'b111111111;
assign micromatriz[98][41] = 9'b111111111;
assign micromatriz[98][42] = 9'b111111111;
assign micromatriz[98][43] = 9'b111111111;
assign micromatriz[98][44] = 9'b111111111;
assign micromatriz[98][45] = 9'b111111111;
assign micromatriz[98][46] = 9'b111111111;
assign micromatriz[98][47] = 9'b111111111;
assign micromatriz[98][48] = 9'b111111111;
assign micromatriz[98][49] = 9'b111111111;
assign micromatriz[98][50] = 9'b111111111;
assign micromatriz[98][51] = 9'b111111111;
assign micromatriz[98][52] = 9'b111111111;
assign micromatriz[98][53] = 9'b111111111;
assign micromatriz[98][54] = 9'b111111111;
assign micromatriz[98][55] = 9'b111111111;
assign micromatriz[98][56] = 9'b111111111;
assign micromatriz[98][57] = 9'b111111111;
assign micromatriz[98][58] = 9'b111111111;
assign micromatriz[98][59] = 9'b111111111;
assign micromatriz[98][60] = 9'b111111111;
assign micromatriz[98][61] = 9'b111111111;
assign micromatriz[98][62] = 9'b111111111;
assign micromatriz[98][63] = 9'b111111111;
assign micromatriz[98][64] = 9'b111111111;
assign micromatriz[98][65] = 9'b111111111;
assign micromatriz[98][66] = 9'b111111111;
assign micromatriz[98][67] = 9'b111111111;
assign micromatriz[98][68] = 9'b111111111;
assign micromatriz[98][69] = 9'b111111111;
assign micromatriz[98][70] = 9'b111111111;
assign micromatriz[98][71] = 9'b111111111;
assign micromatriz[98][72] = 9'b111111111;
assign micromatriz[98][73] = 9'b111111111;
assign micromatriz[98][74] = 9'b111111111;
assign micromatriz[98][75] = 9'b111111111;
assign micromatriz[98][76] = 9'b111111111;
assign micromatriz[98][77] = 9'b111111111;
assign micromatriz[98][78] = 9'b111111111;
assign micromatriz[98][79] = 9'b111111111;
assign micromatriz[98][80] = 9'b111111111;
assign micromatriz[98][81] = 9'b111111111;
assign micromatriz[98][82] = 9'b111111111;
assign micromatriz[98][83] = 9'b111111111;
assign micromatriz[98][84] = 9'b111111111;
assign micromatriz[98][85] = 9'b111111111;
assign micromatriz[98][86] = 9'b111111111;
assign micromatriz[98][87] = 9'b111111111;
assign micromatriz[98][88] = 9'b111111111;
assign micromatriz[98][89] = 9'b111111111;
assign micromatriz[98][90] = 9'b111111111;
assign micromatriz[98][91] = 9'b111111111;
assign micromatriz[98][92] = 9'b111111111;
assign micromatriz[98][93] = 9'b111111111;
assign micromatriz[98][94] = 9'b111111111;
assign micromatriz[98][95] = 9'b111111111;
assign micromatriz[98][96] = 9'b111111111;
assign micromatriz[98][97] = 9'b111111111;
assign micromatriz[98][98] = 9'b111111111;
assign micromatriz[98][99] = 9'b111111111;
assign micromatriz[99][0] = 9'b111111111;
assign micromatriz[99][1] = 9'b111111111;
assign micromatriz[99][2] = 9'b111111111;
assign micromatriz[99][3] = 9'b111111111;
assign micromatriz[99][4] = 9'b111111111;
assign micromatriz[99][5] = 9'b111111111;
assign micromatriz[99][6] = 9'b111111111;
assign micromatriz[99][7] = 9'b111111111;
assign micromatriz[99][8] = 9'b111111111;
assign micromatriz[99][9] = 9'b111111111;
assign micromatriz[99][10] = 9'b111111111;
assign micromatriz[99][11] = 9'b111111111;
assign micromatriz[99][12] = 9'b111111111;
assign micromatriz[99][13] = 9'b111111111;
assign micromatriz[99][14] = 9'b111111111;
assign micromatriz[99][15] = 9'b111111111;
assign micromatriz[99][16] = 9'b111111111;
assign micromatriz[99][17] = 9'b111111111;
assign micromatriz[99][18] = 9'b111111111;
assign micromatriz[99][19] = 9'b111111111;
assign micromatriz[99][20] = 9'b111111111;
assign micromatriz[99][21] = 9'b111111111;
assign micromatriz[99][22] = 9'b111111111;
assign micromatriz[99][23] = 9'b111111111;
assign micromatriz[99][24] = 9'b111111111;
assign micromatriz[99][25] = 9'b111111111;
assign micromatriz[99][26] = 9'b111111111;
assign micromatriz[99][27] = 9'b111111111;
assign micromatriz[99][28] = 9'b111111111;
assign micromatriz[99][29] = 9'b111111111;
assign micromatriz[99][30] = 9'b111111111;
assign micromatriz[99][31] = 9'b111111111;
assign micromatriz[99][32] = 9'b111111111;
assign micromatriz[99][33] = 9'b111111111;
assign micromatriz[99][34] = 9'b111111111;
assign micromatriz[99][35] = 9'b111111111;
assign micromatriz[99][36] = 9'b111111111;
assign micromatriz[99][37] = 9'b111111111;
assign micromatriz[99][38] = 9'b111111111;
assign micromatriz[99][39] = 9'b111111111;
assign micromatriz[99][40] = 9'b111111111;
assign micromatriz[99][41] = 9'b111111111;
assign micromatriz[99][42] = 9'b111111111;
assign micromatriz[99][43] = 9'b111111111;
assign micromatriz[99][44] = 9'b111111111;
assign micromatriz[99][45] = 9'b111111111;
assign micromatriz[99][46] = 9'b111111111;
assign micromatriz[99][47] = 9'b111111111;
assign micromatriz[99][48] = 9'b111111111;
assign micromatriz[99][49] = 9'b111111111;
assign micromatriz[99][50] = 9'b111111111;
assign micromatriz[99][51] = 9'b111111111;
assign micromatriz[99][52] = 9'b111111111;
assign micromatriz[99][53] = 9'b111111111;
assign micromatriz[99][54] = 9'b111111111;
assign micromatriz[99][55] = 9'b111111111;
assign micromatriz[99][56] = 9'b111111111;
assign micromatriz[99][57] = 9'b111111111;
assign micromatriz[99][58] = 9'b111111111;
assign micromatriz[99][59] = 9'b111111111;
assign micromatriz[99][60] = 9'b111111111;
assign micromatriz[99][61] = 9'b111111111;
assign micromatriz[99][62] = 9'b111111111;
assign micromatriz[99][63] = 9'b111111111;
assign micromatriz[99][64] = 9'b111111111;
assign micromatriz[99][65] = 9'b111111111;
assign micromatriz[99][66] = 9'b111111111;
assign micromatriz[99][67] = 9'b111111111;
assign micromatriz[99][68] = 9'b111111111;
assign micromatriz[99][69] = 9'b111111111;
assign micromatriz[99][70] = 9'b111111111;
assign micromatriz[99][71] = 9'b111111111;
assign micromatriz[99][72] = 9'b111111111;
assign micromatriz[99][73] = 9'b111111111;
assign micromatriz[99][74] = 9'b111111111;
assign micromatriz[99][75] = 9'b111111111;
assign micromatriz[99][76] = 9'b111111111;
assign micromatriz[99][77] = 9'b111111111;
assign micromatriz[99][78] = 9'b111111111;
assign micromatriz[99][79] = 9'b111111111;
assign micromatriz[99][80] = 9'b111111111;
assign micromatriz[99][81] = 9'b111111111;
assign micromatriz[99][82] = 9'b111111111;
assign micromatriz[99][83] = 9'b111111111;
assign micromatriz[99][84] = 9'b111111111;
assign micromatriz[99][85] = 9'b111111111;
assign micromatriz[99][86] = 9'b111111111;
assign micromatriz[99][87] = 9'b111111111;
assign micromatriz[99][88] = 9'b111111111;
assign micromatriz[99][89] = 9'b111111111;
assign micromatriz[99][90] = 9'b111111111;
assign micromatriz[99][91] = 9'b111111111;
assign micromatriz[99][92] = 9'b111111111;
assign micromatriz[99][93] = 9'b111111111;
assign micromatriz[99][94] = 9'b111111111;
assign micromatriz[99][95] = 9'b111111111;
assign micromatriz[99][96] = 9'b111111111;
assign micromatriz[99][97] = 9'b111111111;
assign micromatriz[99][98] = 9'b111111111;
assign micromatriz[99][99] = 9'b111111111;
//Total de Lineas = 10000
endmodule




