`timescale 1ns / 1ps
module prueba_2 (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (micromatr[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= micromatr[vcount- posy][hcount- posx][7:5];
				green <= micromatr[vcount- posy][hcount- posx][4:2];
            blue 	<= micromatr[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 100;
parameter RESOLUCION_Y = 50;
wire [8:0] micromatr[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign micromatr[0][0] = 9'b111111111;
assign micromatr[0][1] = 9'b111111111;
assign micromatr[0][2] = 9'b111111111;
assign micromatr[0][3] = 9'b111111111;
assign micromatr[0][4] = 9'b111111111;
assign micromatr[0][5] = 9'b111111111;
assign micromatr[0][6] = 9'b111111111;
assign micromatr[0][7] = 9'b111111111;
assign micromatr[0][8] = 9'b111111111;
assign micromatr[0][9] = 9'b111111111;
assign micromatr[0][10] = 9'b111111111;
assign micromatr[0][11] = 9'b111111111;
assign micromatr[0][12] = 9'b111111111;
assign micromatr[0][13] = 9'b111111111;
assign micromatr[0][14] = 9'b111111111;
assign micromatr[0][15] = 9'b111111111;
assign micromatr[0][16] = 9'b111111111;
assign micromatr[0][17] = 9'b111111111;
assign micromatr[0][18] = 9'b111111111;
assign micromatr[0][19] = 9'b111111111;
assign micromatr[0][20] = 9'b111111111;
assign micromatr[0][21] = 9'b111111111;
assign micromatr[0][22] = 9'b111111111;
assign micromatr[0][23] = 9'b111111111;
assign micromatr[0][24] = 9'b111111111;
assign micromatr[0][25] = 9'b111111111;
assign micromatr[0][26] = 9'b111111111;
assign micromatr[0][27] = 9'b111111111;
assign micromatr[0][28] = 9'b111111111;
assign micromatr[0][29] = 9'b111111111;
assign micromatr[0][30] = 9'b111111111;
assign micromatr[0][31] = 9'b111111111;
assign micromatr[0][32] = 9'b111111111;
assign micromatr[0][33] = 9'b111111111;
assign micromatr[0][34] = 9'b111111111;
assign micromatr[0][35] = 9'b111111111;
assign micromatr[0][36] = 9'b111111111;
assign micromatr[0][37] = 9'b111111111;
assign micromatr[0][38] = 9'b111111111;
assign micromatr[0][39] = 9'b111111111;
assign micromatr[0][40] = 9'b111111111;
assign micromatr[0][41] = 9'b111111111;
assign micromatr[0][42] = 9'b111111111;
assign micromatr[0][43] = 9'b111111111;
assign micromatr[0][44] = 9'b111111111;
assign micromatr[0][45] = 9'b111111111;
assign micromatr[0][46] = 9'b111111111;
assign micromatr[0][47] = 9'b111111111;
assign micromatr[0][48] = 9'b111111111;
assign micromatr[0][49] = 9'b111111111;
assign micromatr[0][50] = 9'b111111111;
assign micromatr[0][51] = 9'b111111111;
assign micromatr[0][52] = 9'b111111111;
assign micromatr[0][53] = 9'b111111111;
assign micromatr[0][54] = 9'b111111111;
assign micromatr[0][55] = 9'b111111111;
assign micromatr[0][56] = 9'b111111111;
assign micromatr[0][57] = 9'b111111111;
assign micromatr[0][58] = 9'b111111111;
assign micromatr[0][59] = 9'b111111111;
assign micromatr[0][60] = 9'b111111111;
assign micromatr[0][61] = 9'b111111111;
assign micromatr[0][62] = 9'b111111111;
assign micromatr[0][63] = 9'b111111111;
assign micromatr[0][64] = 9'b111111111;
assign micromatr[0][65] = 9'b111111111;
assign micromatr[0][66] = 9'b111111111;
assign micromatr[0][67] = 9'b111111111;
assign micromatr[0][68] = 9'b111111111;
assign micromatr[0][69] = 9'b111111111;
assign micromatr[0][70] = 9'b111111111;
assign micromatr[0][71] = 9'b111111111;
assign micromatr[0][72] = 9'b111111111;
assign micromatr[0][73] = 9'b111111111;
assign micromatr[0][74] = 9'b111111111;
assign micromatr[0][75] = 9'b111111111;
assign micromatr[0][76] = 9'b111111111;
assign micromatr[0][77] = 9'b111111111;
assign micromatr[0][78] = 9'b111111111;
assign micromatr[0][79] = 9'b111111111;
assign micromatr[0][80] = 9'b111111111;
assign micromatr[0][81] = 9'b111111111;
assign micromatr[0][82] = 9'b111111111;
assign micromatr[0][83] = 9'b111111111;
assign micromatr[0][84] = 9'b111111111;
assign micromatr[0][85] = 9'b111111111;
assign micromatr[0][86] = 9'b111111111;
assign micromatr[0][87] = 9'b111111111;
assign micromatr[0][88] = 9'b111111111;
assign micromatr[0][89] = 9'b111111111;
assign micromatr[0][90] = 9'b111111111;
assign micromatr[0][91] = 9'b111111111;
assign micromatr[0][92] = 9'b111111111;
assign micromatr[0][93] = 9'b111111111;
assign micromatr[0][94] = 9'b111111111;
assign micromatr[0][95] = 9'b111111111;
assign micromatr[0][96] = 9'b111111111;
assign micromatr[0][97] = 9'b111111111;
assign micromatr[0][98] = 9'b111111111;
assign micromatr[0][99] = 9'b111111111;
assign micromatr[1][0] = 9'b111111111;
assign micromatr[1][1] = 9'b111111111;
assign micromatr[1][2] = 9'b111111111;
assign micromatr[1][3] = 9'b111111111;
assign micromatr[1][4] = 9'b111111111;
assign micromatr[1][5] = 9'b111111111;
assign micromatr[1][6] = 9'b111111111;
assign micromatr[1][7] = 9'b111111111;
assign micromatr[1][8] = 9'b111111111;
assign micromatr[1][9] = 9'b111111111;
assign micromatr[1][10] = 9'b111111111;
assign micromatr[1][11] = 9'b111111111;
assign micromatr[1][12] = 9'b111111111;
assign micromatr[1][13] = 9'b111111111;
assign micromatr[1][14] = 9'b111111111;
assign micromatr[1][15] = 9'b111111111;
assign micromatr[1][16] = 9'b111111111;
assign micromatr[1][17] = 9'b111111111;
assign micromatr[1][18] = 9'b111111111;
assign micromatr[1][19] = 9'b111111111;
assign micromatr[1][20] = 9'b111111111;
assign micromatr[1][21] = 9'b111111111;
assign micromatr[1][22] = 9'b111111111;
assign micromatr[1][23] = 9'b111111111;
assign micromatr[1][24] = 9'b111111111;
assign micromatr[1][25] = 9'b111111111;
assign micromatr[1][26] = 9'b111111111;
assign micromatr[1][27] = 9'b111111111;
assign micromatr[1][28] = 9'b111111111;
assign micromatr[1][29] = 9'b111111111;
assign micromatr[1][30] = 9'b111111111;
assign micromatr[1][31] = 9'b111111111;
assign micromatr[1][32] = 9'b111111111;
assign micromatr[1][33] = 9'b111111111;
assign micromatr[1][34] = 9'b111111111;
assign micromatr[1][35] = 9'b111111111;
assign micromatr[1][36] = 9'b111111111;
assign micromatr[1][37] = 9'b111111111;
assign micromatr[1][38] = 9'b111111111;
assign micromatr[1][39] = 9'b111111111;
assign micromatr[1][40] = 9'b111111111;
assign micromatr[1][41] = 9'b111111111;
assign micromatr[1][42] = 9'b111111111;
assign micromatr[1][43] = 9'b111111111;
assign micromatr[1][44] = 9'b111111111;
assign micromatr[1][45] = 9'b111111111;
assign micromatr[1][46] = 9'b111111111;
assign micromatr[1][47] = 9'b111111111;
assign micromatr[1][48] = 9'b111111111;
assign micromatr[1][49] = 9'b111111111;
assign micromatr[1][50] = 9'b111111111;
assign micromatr[1][51] = 9'b111111111;
assign micromatr[1][52] = 9'b111111111;
assign micromatr[1][53] = 9'b111111111;
assign micromatr[1][54] = 9'b111111111;
assign micromatr[1][55] = 9'b111111111;
assign micromatr[1][56] = 9'b111111111;
assign micromatr[1][57] = 9'b111111111;
assign micromatr[1][58] = 9'b111111111;
assign micromatr[1][59] = 9'b111111111;
assign micromatr[1][60] = 9'b111111111;
assign micromatr[1][61] = 9'b111111111;
assign micromatr[1][62] = 9'b111111111;
assign micromatr[1][63] = 9'b111111111;
assign micromatr[1][64] = 9'b111111111;
assign micromatr[1][65] = 9'b111111111;
assign micromatr[1][66] = 9'b111111111;
assign micromatr[1][67] = 9'b111111111;
assign micromatr[1][68] = 9'b111111111;
assign micromatr[1][69] = 9'b111111111;
assign micromatr[1][70] = 9'b111111111;
assign micromatr[1][71] = 9'b111111111;
assign micromatr[1][72] = 9'b111111111;
assign micromatr[1][73] = 9'b111111111;
assign micromatr[1][74] = 9'b111111111;
assign micromatr[1][75] = 9'b111111111;
assign micromatr[1][76] = 9'b111111111;
assign micromatr[1][77] = 9'b111111111;
assign micromatr[1][78] = 9'b111111111;
assign micromatr[1][79] = 9'b111111111;
assign micromatr[1][80] = 9'b111111111;
assign micromatr[1][81] = 9'b111111111;
assign micromatr[1][82] = 9'b111111111;
assign micromatr[1][83] = 9'b111111111;
assign micromatr[1][84] = 9'b111111111;
assign micromatr[1][85] = 9'b111111111;
assign micromatr[1][86] = 9'b111111111;
assign micromatr[1][87] = 9'b111111111;
assign micromatr[1][88] = 9'b111111111;
assign micromatr[1][89] = 9'b111111111;
assign micromatr[1][90] = 9'b111111111;
assign micromatr[1][91] = 9'b111111111;
assign micromatr[1][92] = 9'b111111111;
assign micromatr[1][93] = 9'b111111111;
assign micromatr[1][94] = 9'b111111111;
assign micromatr[1][95] = 9'b111111111;
assign micromatr[1][96] = 9'b111111111;
assign micromatr[1][97] = 9'b111111111;
assign micromatr[1][98] = 9'b111111111;
assign micromatr[1][99] = 9'b111111111;
assign micromatr[2][0] = 9'b111111111;
assign micromatr[2][1] = 9'b111111111;
assign micromatr[2][2] = 9'b111111111;
assign micromatr[2][3] = 9'b111111111;
assign micromatr[2][4] = 9'b111111111;
assign micromatr[2][5] = 9'b111111111;
assign micromatr[2][6] = 9'b111111111;
assign micromatr[2][7] = 9'b111111111;
assign micromatr[2][8] = 9'b111111111;
assign micromatr[2][9] = 9'b111111111;
assign micromatr[2][10] = 9'b111111111;
assign micromatr[2][11] = 9'b111111111;
assign micromatr[2][12] = 9'b111111111;
assign micromatr[2][13] = 9'b111111111;
assign micromatr[2][14] = 9'b111111111;
assign micromatr[2][15] = 9'b111111111;
assign micromatr[2][16] = 9'b111111111;
assign micromatr[2][17] = 9'b111111111;
assign micromatr[2][18] = 9'b111111111;
assign micromatr[2][19] = 9'b111111111;
assign micromatr[2][20] = 9'b111111111;
assign micromatr[2][21] = 9'b111111111;
assign micromatr[2][22] = 9'b111111111;
assign micromatr[2][23] = 9'b111111111;
assign micromatr[2][24] = 9'b111111111;
assign micromatr[2][25] = 9'b111111111;
assign micromatr[2][26] = 9'b111111111;
assign micromatr[2][27] = 9'b111111111;
assign micromatr[2][28] = 9'b111111111;
assign micromatr[2][29] = 9'b111111111;
assign micromatr[2][30] = 9'b111111111;
assign micromatr[2][31] = 9'b111111111;
assign micromatr[2][32] = 9'b111111111;
assign micromatr[2][33] = 9'b111111111;
assign micromatr[2][34] = 9'b111111111;
assign micromatr[2][35] = 9'b111111111;
assign micromatr[2][36] = 9'b111111111;
assign micromatr[2][37] = 9'b111111111;
assign micromatr[2][38] = 9'b111111111;
assign micromatr[2][39] = 9'b111111111;
assign micromatr[2][40] = 9'b111111111;
assign micromatr[2][41] = 9'b111111111;
assign micromatr[2][42] = 9'b111111111;
assign micromatr[2][43] = 9'b111111111;
assign micromatr[2][44] = 9'b111111111;
assign micromatr[2][45] = 9'b111111111;
assign micromatr[2][46] = 9'b111111111;
assign micromatr[2][47] = 9'b111111111;
assign micromatr[2][48] = 9'b111111111;
assign micromatr[2][49] = 9'b111111111;
assign micromatr[2][50] = 9'b111111111;
assign micromatr[2][51] = 9'b111111111;
assign micromatr[2][52] = 9'b111111111;
assign micromatr[2][53] = 9'b111111111;
assign micromatr[2][54] = 9'b111111111;
assign micromatr[2][55] = 9'b111111111;
assign micromatr[2][56] = 9'b111111111;
assign micromatr[2][57] = 9'b111111111;
assign micromatr[2][58] = 9'b111111111;
assign micromatr[2][59] = 9'b111111111;
assign micromatr[2][60] = 9'b111111111;
assign micromatr[2][61] = 9'b111111111;
assign micromatr[2][62] = 9'b111111111;
assign micromatr[2][63] = 9'b111111111;
assign micromatr[2][64] = 9'b111111111;
assign micromatr[2][65] = 9'b111111111;
assign micromatr[2][66] = 9'b111111111;
assign micromatr[2][67] = 9'b111111111;
assign micromatr[2][68] = 9'b111111111;
assign micromatr[2][69] = 9'b111111111;
assign micromatr[2][70] = 9'b111111111;
assign micromatr[2][71] = 9'b111111111;
assign micromatr[2][72] = 9'b111111111;
assign micromatr[2][73] = 9'b111111111;
assign micromatr[2][74] = 9'b111111111;
assign micromatr[2][75] = 9'b111111111;
assign micromatr[2][76] = 9'b111111111;
assign micromatr[2][77] = 9'b111111111;
assign micromatr[2][78] = 9'b111111111;
assign micromatr[2][79] = 9'b111111111;
assign micromatr[2][80] = 9'b111111111;
assign micromatr[2][81] = 9'b111111111;
assign micromatr[2][82] = 9'b111111111;
assign micromatr[2][83] = 9'b111111111;
assign micromatr[2][84] = 9'b111111111;
assign micromatr[2][85] = 9'b111111111;
assign micromatr[2][86] = 9'b111111111;
assign micromatr[2][87] = 9'b111111111;
assign micromatr[2][88] = 9'b111111111;
assign micromatr[2][89] = 9'b111111111;
assign micromatr[2][90] = 9'b111111111;
assign micromatr[2][91] = 9'b111111111;
assign micromatr[2][92] = 9'b111111111;
assign micromatr[2][93] = 9'b111111111;
assign micromatr[2][94] = 9'b111111111;
assign micromatr[2][95] = 9'b111111111;
assign micromatr[2][96] = 9'b111111111;
assign micromatr[2][97] = 9'b111111111;
assign micromatr[2][98] = 9'b111111111;
assign micromatr[2][99] = 9'b111111111;
assign micromatr[3][0] = 9'b111111111;
assign micromatr[3][1] = 9'b111111111;
assign micromatr[3][2] = 9'b111111111;
assign micromatr[3][3] = 9'b111111111;
assign micromatr[3][4] = 9'b111111111;
assign micromatr[3][5] = 9'b111111111;
assign micromatr[3][6] = 9'b111111111;
assign micromatr[3][7] = 9'b111111111;
assign micromatr[3][8] = 9'b111111111;
assign micromatr[3][9] = 9'b111111111;
assign micromatr[3][10] = 9'b111111111;
assign micromatr[3][11] = 9'b111111111;
assign micromatr[3][12] = 9'b111111111;
assign micromatr[3][13] = 9'b111111111;
assign micromatr[3][14] = 9'b111111111;
assign micromatr[3][15] = 9'b111111111;
assign micromatr[3][16] = 9'b111111111;
assign micromatr[3][17] = 9'b111111111;
assign micromatr[3][18] = 9'b111111111;
assign micromatr[3][19] = 9'b111111111;
assign micromatr[3][20] = 9'b111111111;
assign micromatr[3][21] = 9'b111111111;
assign micromatr[3][22] = 9'b111111111;
assign micromatr[3][23] = 9'b111111111;
assign micromatr[3][24] = 9'b111111111;
assign micromatr[3][25] = 9'b111111111;
assign micromatr[3][26] = 9'b111111111;
assign micromatr[3][27] = 9'b111111111;
assign micromatr[3][28] = 9'b111111111;
assign micromatr[3][29] = 9'b111111111;
assign micromatr[3][30] = 9'b111111111;
assign micromatr[3][31] = 9'b111111111;
assign micromatr[3][32] = 9'b111111111;
assign micromatr[3][33] = 9'b111111111;
assign micromatr[3][34] = 9'b111111111;
assign micromatr[3][35] = 9'b111111111;
assign micromatr[3][36] = 9'b111111111;
assign micromatr[3][37] = 9'b111111111;
assign micromatr[3][38] = 9'b111111111;
assign micromatr[3][39] = 9'b111111111;
assign micromatr[3][40] = 9'b111111111;
assign micromatr[3][41] = 9'b111111111;
assign micromatr[3][42] = 9'b111111111;
assign micromatr[3][43] = 9'b111111111;
assign micromatr[3][44] = 9'b111111111;
assign micromatr[3][45] = 9'b111111111;
assign micromatr[3][46] = 9'b111111111;
assign micromatr[3][47] = 9'b111111111;
assign micromatr[3][48] = 9'b111111111;
assign micromatr[3][49] = 9'b111111111;
assign micromatr[3][50] = 9'b111111111;
assign micromatr[3][51] = 9'b111111111;
assign micromatr[3][52] = 9'b111111111;
assign micromatr[3][53] = 9'b111111111;
assign micromatr[3][54] = 9'b111111111;
assign micromatr[3][55] = 9'b111111111;
assign micromatr[3][56] = 9'b111111111;
assign micromatr[3][57] = 9'b111111111;
assign micromatr[3][58] = 9'b111111111;
assign micromatr[3][59] = 9'b111111111;
assign micromatr[3][60] = 9'b111111111;
assign micromatr[3][61] = 9'b111111111;
assign micromatr[3][62] = 9'b111111111;
assign micromatr[3][63] = 9'b111111111;
assign micromatr[3][64] = 9'b111111111;
assign micromatr[3][65] = 9'b111111111;
assign micromatr[3][66] = 9'b111111111;
assign micromatr[3][67] = 9'b111111111;
assign micromatr[3][68] = 9'b111111111;
assign micromatr[3][69] = 9'b111111111;
assign micromatr[3][70] = 9'b111111111;
assign micromatr[3][71] = 9'b111111111;
assign micromatr[3][72] = 9'b111111111;
assign micromatr[3][73] = 9'b111111111;
assign micromatr[3][74] = 9'b111111111;
assign micromatr[3][75] = 9'b111111111;
assign micromatr[3][76] = 9'b111111111;
assign micromatr[3][77] = 9'b111111111;
assign micromatr[3][78] = 9'b111111111;
assign micromatr[3][79] = 9'b111111111;
assign micromatr[3][80] = 9'b111111111;
assign micromatr[3][81] = 9'b111111111;
assign micromatr[3][82] = 9'b111111111;
assign micromatr[3][83] = 9'b111111111;
assign micromatr[3][84] = 9'b111111111;
assign micromatr[3][85] = 9'b111111111;
assign micromatr[3][86] = 9'b111111111;
assign micromatr[3][87] = 9'b111111111;
assign micromatr[3][88] = 9'b111111111;
assign micromatr[3][89] = 9'b111111111;
assign micromatr[3][90] = 9'b111111111;
assign micromatr[3][91] = 9'b111111111;
assign micromatr[3][92] = 9'b111111111;
assign micromatr[3][93] = 9'b111111111;
assign micromatr[3][94] = 9'b111111111;
assign micromatr[3][95] = 9'b111111111;
assign micromatr[3][96] = 9'b111111111;
assign micromatr[3][97] = 9'b111111111;
assign micromatr[3][98] = 9'b111111111;
assign micromatr[3][99] = 9'b111111111;
assign micromatr[4][0] = 9'b111111111;
assign micromatr[4][1] = 9'b111111111;
assign micromatr[4][2] = 9'b111111111;
assign micromatr[4][3] = 9'b111111111;
assign micromatr[4][4] = 9'b111111111;
assign micromatr[4][5] = 9'b111111111;
assign micromatr[4][6] = 9'b111111111;
assign micromatr[4][7] = 9'b111111111;
assign micromatr[4][8] = 9'b111111111;
assign micromatr[4][9] = 9'b111111111;
assign micromatr[4][10] = 9'b111111111;
assign micromatr[4][11] = 9'b111111111;
assign micromatr[4][12] = 9'b111111111;
assign micromatr[4][13] = 9'b111111111;
assign micromatr[4][14] = 9'b111111111;
assign micromatr[4][15] = 9'b111111111;
assign micromatr[4][16] = 9'b111111111;
assign micromatr[4][17] = 9'b111111111;
assign micromatr[4][18] = 9'b111111111;
assign micromatr[4][19] = 9'b111111111;
assign micromatr[4][20] = 9'b111111111;
assign micromatr[4][21] = 9'b111111111;
assign micromatr[4][22] = 9'b111111111;
assign micromatr[4][23] = 9'b111111111;
assign micromatr[4][24] = 9'b111111111;
assign micromatr[4][25] = 9'b111111111;
assign micromatr[4][26] = 9'b111111111;
assign micromatr[4][27] = 9'b111111111;
assign micromatr[4][28] = 9'b111111111;
assign micromatr[4][29] = 9'b111111111;
assign micromatr[4][30] = 9'b111111111;
assign micromatr[4][31] = 9'b111111111;
assign micromatr[4][32] = 9'b111111111;
assign micromatr[4][33] = 9'b111111111;
assign micromatr[4][34] = 9'b111111111;
assign micromatr[4][35] = 9'b111111111;
assign micromatr[4][36] = 9'b111111111;
assign micromatr[4][37] = 9'b111111111;
assign micromatr[4][38] = 9'b111111111;
assign micromatr[4][39] = 9'b111111111;
assign micromatr[4][40] = 9'b111111111;
assign micromatr[4][41] = 9'b111111111;
assign micromatr[4][42] = 9'b111111111;
assign micromatr[4][43] = 9'b111111111;
assign micromatr[4][44] = 9'b111111111;
assign micromatr[4][45] = 9'b111111111;
assign micromatr[4][46] = 9'b111111111;
assign micromatr[4][47] = 9'b111111111;
assign micromatr[4][48] = 9'b111111111;
assign micromatr[4][49] = 9'b111111111;
assign micromatr[4][50] = 9'b111111111;
assign micromatr[4][51] = 9'b111111111;
assign micromatr[4][52] = 9'b111111111;
assign micromatr[4][53] = 9'b111111111;
assign micromatr[4][54] = 9'b111111111;
assign micromatr[4][55] = 9'b111111111;
assign micromatr[4][56] = 9'b111111111;
assign micromatr[4][57] = 9'b111111111;
assign micromatr[4][58] = 9'b111111111;
assign micromatr[4][59] = 9'b111111111;
assign micromatr[4][60] = 9'b111111111;
assign micromatr[4][61] = 9'b111111111;
assign micromatr[4][62] = 9'b111111111;
assign micromatr[4][63] = 9'b111111111;
assign micromatr[4][64] = 9'b111111111;
assign micromatr[4][65] = 9'b111111111;
assign micromatr[4][66] = 9'b111111111;
assign micromatr[4][67] = 9'b111111111;
assign micromatr[4][68] = 9'b111111111;
assign micromatr[4][69] = 9'b111111111;
assign micromatr[4][70] = 9'b111111111;
assign micromatr[4][71] = 9'b111111111;
assign micromatr[4][72] = 9'b111111111;
assign micromatr[4][73] = 9'b111111111;
assign micromatr[4][74] = 9'b111111111;
assign micromatr[4][75] = 9'b111111111;
assign micromatr[4][76] = 9'b111111111;
assign micromatr[4][77] = 9'b111111111;
assign micromatr[4][78] = 9'b111111111;
assign micromatr[4][79] = 9'b111111111;
assign micromatr[4][80] = 9'b111111111;
assign micromatr[4][81] = 9'b111111111;
assign micromatr[4][82] = 9'b111111111;
assign micromatr[4][83] = 9'b111111111;
assign micromatr[4][84] = 9'b111111111;
assign micromatr[4][85] = 9'b111111111;
assign micromatr[4][86] = 9'b111111111;
assign micromatr[4][87] = 9'b111111111;
assign micromatr[4][88] = 9'b111111111;
assign micromatr[4][89] = 9'b111111111;
assign micromatr[4][90] = 9'b111111111;
assign micromatr[4][91] = 9'b111111111;
assign micromatr[4][92] = 9'b111111111;
assign micromatr[4][93] = 9'b111111111;
assign micromatr[4][94] = 9'b111111111;
assign micromatr[4][95] = 9'b111111111;
assign micromatr[4][96] = 9'b111111111;
assign micromatr[4][97] = 9'b111111111;
assign micromatr[4][98] = 9'b111111111;
assign micromatr[4][99] = 9'b111111111;
assign micromatr[5][0] = 9'b111111111;
assign micromatr[5][1] = 9'b111111111;
assign micromatr[5][2] = 9'b111111111;
assign micromatr[5][3] = 9'b111111111;
assign micromatr[5][4] = 9'b111111111;
assign micromatr[5][5] = 9'b111111111;
assign micromatr[5][6] = 9'b111111111;
assign micromatr[5][7] = 9'b111111111;
assign micromatr[5][8] = 9'b111111111;
assign micromatr[5][9] = 9'b111111111;
assign micromatr[5][10] = 9'b111111111;
assign micromatr[5][11] = 9'b111111111;
assign micromatr[5][12] = 9'b111111111;
assign micromatr[5][13] = 9'b111111111;
assign micromatr[5][14] = 9'b111111111;
assign micromatr[5][15] = 9'b111111111;
assign micromatr[5][16] = 9'b111111111;
assign micromatr[5][17] = 9'b111111111;
assign micromatr[5][18] = 9'b111111111;
assign micromatr[5][19] = 9'b111111111;
assign micromatr[5][20] = 9'b111111111;
assign micromatr[5][21] = 9'b111111111;
assign micromatr[5][22] = 9'b111111111;
assign micromatr[5][23] = 9'b111111111;
assign micromatr[5][24] = 9'b111111111;
assign micromatr[5][25] = 9'b111111111;
assign micromatr[5][26] = 9'b111111111;
assign micromatr[5][27] = 9'b111111111;
assign micromatr[5][28] = 9'b111111111;
assign micromatr[5][29] = 9'b111111111;
assign micromatr[5][30] = 9'b111111111;
assign micromatr[5][31] = 9'b111111111;
assign micromatr[5][32] = 9'b111111111;
assign micromatr[5][33] = 9'b111111111;
assign micromatr[5][34] = 9'b111111111;
assign micromatr[5][35] = 9'b111111111;
assign micromatr[5][36] = 9'b111111111;
assign micromatr[5][37] = 9'b111111111;
assign micromatr[5][38] = 9'b111111111;
assign micromatr[5][39] = 9'b111111111;
assign micromatr[5][40] = 9'b111111111;
assign micromatr[5][41] = 9'b111111111;
assign micromatr[5][42] = 9'b111111111;
assign micromatr[5][43] = 9'b111111111;
assign micromatr[5][44] = 9'b111111111;
assign micromatr[5][45] = 9'b111111111;
assign micromatr[5][46] = 9'b111111111;
assign micromatr[5][47] = 9'b111111111;
assign micromatr[5][48] = 9'b111111111;
assign micromatr[5][49] = 9'b111111111;
assign micromatr[5][50] = 9'b111111111;
assign micromatr[5][51] = 9'b111111111;
assign micromatr[5][52] = 9'b111111111;
assign micromatr[5][53] = 9'b111111111;
assign micromatr[5][54] = 9'b111111111;
assign micromatr[5][55] = 9'b111111111;
assign micromatr[5][56] = 9'b111111111;
assign micromatr[5][57] = 9'b111111111;
assign micromatr[5][58] = 9'b111111111;
assign micromatr[5][59] = 9'b111111111;
assign micromatr[5][60] = 9'b111111111;
assign micromatr[5][61] = 9'b111111111;
assign micromatr[5][62] = 9'b111111111;
assign micromatr[5][63] = 9'b111111111;
assign micromatr[5][64] = 9'b111111111;
assign micromatr[5][65] = 9'b111111111;
assign micromatr[5][66] = 9'b111111111;
assign micromatr[5][67] = 9'b111111111;
assign micromatr[5][68] = 9'b111111111;
assign micromatr[5][69] = 9'b111111111;
assign micromatr[5][70] = 9'b111111111;
assign micromatr[5][71] = 9'b111111111;
assign micromatr[5][72] = 9'b111111111;
assign micromatr[5][73] = 9'b111111111;
assign micromatr[5][74] = 9'b111111111;
assign micromatr[5][75] = 9'b111111111;
assign micromatr[5][76] = 9'b111111111;
assign micromatr[5][77] = 9'b111111111;
assign micromatr[5][78] = 9'b111111111;
assign micromatr[5][79] = 9'b111111111;
assign micromatr[5][80] = 9'b111111111;
assign micromatr[5][81] = 9'b111111111;
assign micromatr[5][82] = 9'b111111111;
assign micromatr[5][83] = 9'b111111111;
assign micromatr[5][84] = 9'b111111111;
assign micromatr[5][85] = 9'b111111111;
assign micromatr[5][86] = 9'b111111111;
assign micromatr[5][87] = 9'b111111111;
assign micromatr[5][88] = 9'b111111111;
assign micromatr[5][89] = 9'b111111111;
assign micromatr[5][90] = 9'b111111111;
assign micromatr[5][91] = 9'b111111111;
assign micromatr[5][92] = 9'b111111111;
assign micromatr[5][93] = 9'b111111111;
assign micromatr[5][94] = 9'b111111111;
assign micromatr[5][95] = 9'b111111111;
assign micromatr[5][96] = 9'b111111111;
assign micromatr[5][97] = 9'b111111111;
assign micromatr[5][98] = 9'b111111111;
assign micromatr[5][99] = 9'b111111111;
assign micromatr[6][0] = 9'b111111111;
assign micromatr[6][1] = 9'b111111111;
assign micromatr[6][2] = 9'b111111111;
assign micromatr[6][3] = 9'b111111111;
assign micromatr[6][4] = 9'b111111111;
assign micromatr[6][5] = 9'b111111111;
assign micromatr[6][6] = 9'b111111111;
assign micromatr[6][7] = 9'b111111111;
assign micromatr[6][8] = 9'b111111111;
assign micromatr[6][9] = 9'b111111111;
assign micromatr[6][10] = 9'b111111111;
assign micromatr[6][11] = 9'b111111111;
assign micromatr[6][12] = 9'b111111111;
assign micromatr[6][13] = 9'b111111111;
assign micromatr[6][14] = 9'b111111111;
assign micromatr[6][15] = 9'b111111111;
assign micromatr[6][16] = 9'b111111111;
assign micromatr[6][17] = 9'b111111111;
assign micromatr[6][18] = 9'b111111111;
assign micromatr[6][19] = 9'b111111111;
assign micromatr[6][20] = 9'b111111111;
assign micromatr[6][21] = 9'b111111111;
assign micromatr[6][22] = 9'b111111111;
assign micromatr[6][23] = 9'b111111111;
assign micromatr[6][24] = 9'b111111111;
assign micromatr[6][25] = 9'b111111111;
assign micromatr[6][26] = 9'b111111111;
assign micromatr[6][27] = 9'b111111111;
assign micromatr[6][28] = 9'b111111111;
assign micromatr[6][29] = 9'b111111111;
assign micromatr[6][30] = 9'b111111111;
assign micromatr[6][31] = 9'b111111111;
assign micromatr[6][32] = 9'b111111111;
assign micromatr[6][33] = 9'b111111111;
assign micromatr[6][34] = 9'b111111111;
assign micromatr[6][35] = 9'b111111111;
assign micromatr[6][36] = 9'b111111111;
assign micromatr[6][37] = 9'b111111111;
assign micromatr[6][38] = 9'b111111111;
assign micromatr[6][39] = 9'b111111111;
assign micromatr[6][40] = 9'b111111111;
assign micromatr[6][41] = 9'b111111111;
assign micromatr[6][42] = 9'b111111111;
assign micromatr[6][43] = 9'b111111111;
assign micromatr[6][44] = 9'b111111111;
assign micromatr[6][45] = 9'b111111111;
assign micromatr[6][46] = 9'b111111111;
assign micromatr[6][47] = 9'b111111111;
assign micromatr[6][48] = 9'b111111111;
assign micromatr[6][49] = 9'b111111111;
assign micromatr[6][50] = 9'b111111111;
assign micromatr[6][51] = 9'b111111111;
assign micromatr[6][52] = 9'b111111111;
assign micromatr[6][53] = 9'b111111111;
assign micromatr[6][54] = 9'b111111111;
assign micromatr[6][55] = 9'b111111111;
assign micromatr[6][56] = 9'b111111111;
assign micromatr[6][57] = 9'b111111111;
assign micromatr[6][58] = 9'b111111111;
assign micromatr[6][59] = 9'b111111111;
assign micromatr[6][60] = 9'b111111111;
assign micromatr[6][61] = 9'b111111111;
assign micromatr[6][62] = 9'b111111111;
assign micromatr[6][63] = 9'b111111111;
assign micromatr[6][64] = 9'b111111111;
assign micromatr[6][65] = 9'b111111111;
assign micromatr[6][66] = 9'b111111111;
assign micromatr[6][67] = 9'b111111111;
assign micromatr[6][68] = 9'b111111111;
assign micromatr[6][69] = 9'b111111111;
assign micromatr[6][70] = 9'b111111111;
assign micromatr[6][71] = 9'b111111111;
assign micromatr[6][72] = 9'b111111111;
assign micromatr[6][73] = 9'b111111111;
assign micromatr[6][74] = 9'b111111111;
assign micromatr[6][75] = 9'b111111111;
assign micromatr[6][76] = 9'b111111111;
assign micromatr[6][77] = 9'b111111111;
assign micromatr[6][78] = 9'b111111111;
assign micromatr[6][79] = 9'b111111111;
assign micromatr[6][80] = 9'b111111111;
assign micromatr[6][81] = 9'b111111111;
assign micromatr[6][82] = 9'b111111111;
assign micromatr[6][83] = 9'b111111111;
assign micromatr[6][84] = 9'b111111111;
assign micromatr[6][85] = 9'b111111111;
assign micromatr[6][86] = 9'b111111111;
assign micromatr[6][87] = 9'b111111111;
assign micromatr[6][88] = 9'b111111111;
assign micromatr[6][89] = 9'b111111111;
assign micromatr[6][90] = 9'b111111111;
assign micromatr[6][91] = 9'b111111111;
assign micromatr[6][92] = 9'b111111111;
assign micromatr[6][93] = 9'b111111111;
assign micromatr[6][94] = 9'b111111111;
assign micromatr[6][95] = 9'b111111111;
assign micromatr[6][96] = 9'b111111111;
assign micromatr[6][97] = 9'b111111111;
assign micromatr[6][98] = 9'b111111111;
assign micromatr[6][99] = 9'b111111111;
assign micromatr[7][0] = 9'b111111111;
assign micromatr[7][1] = 9'b111111111;
assign micromatr[7][2] = 9'b111111111;
assign micromatr[7][3] = 9'b111111111;
assign micromatr[7][4] = 9'b111111111;
assign micromatr[7][5] = 9'b111111111;
assign micromatr[7][6] = 9'b111111111;
assign micromatr[7][7] = 9'b111111111;
assign micromatr[7][8] = 9'b111111111;
assign micromatr[7][9] = 9'b111111111;
assign micromatr[7][10] = 9'b111111111;
assign micromatr[7][11] = 9'b111111111;
assign micromatr[7][12] = 9'b111111111;
assign micromatr[7][13] = 9'b111111111;
assign micromatr[7][14] = 9'b111111111;
assign micromatr[7][15] = 9'b111111111;
assign micromatr[7][16] = 9'b111111111;
assign micromatr[7][17] = 9'b111111111;
assign micromatr[7][18] = 9'b111111111;
assign micromatr[7][19] = 9'b111111111;
assign micromatr[7][20] = 9'b111111111;
assign micromatr[7][21] = 9'b111111111;
assign micromatr[7][22] = 9'b111111111;
assign micromatr[7][23] = 9'b111111111;
assign micromatr[7][24] = 9'b111111111;
assign micromatr[7][25] = 9'b111111111;
assign micromatr[7][26] = 9'b111111111;
assign micromatr[7][27] = 9'b111111111;
assign micromatr[7][28] = 9'b111111111;
assign micromatr[7][29] = 9'b111111111;
assign micromatr[7][30] = 9'b111111111;
assign micromatr[7][31] = 9'b111111111;
assign micromatr[7][32] = 9'b111111111;
assign micromatr[7][33] = 9'b111111111;
assign micromatr[7][34] = 9'b111111111;
assign micromatr[7][35] = 9'b111111111;
assign micromatr[7][36] = 9'b111111111;
assign micromatr[7][37] = 9'b111111111;
assign micromatr[7][38] = 9'b111111111;
assign micromatr[7][39] = 9'b111111111;
assign micromatr[7][40] = 9'b111111111;
assign micromatr[7][41] = 9'b111111111;
assign micromatr[7][42] = 9'b111111111;
assign micromatr[7][43] = 9'b111111111;
assign micromatr[7][44] = 9'b111111111;
assign micromatr[7][45] = 9'b111111111;
assign micromatr[7][46] = 9'b111111111;
assign micromatr[7][47] = 9'b111111111;
assign micromatr[7][48] = 9'b111111111;
assign micromatr[7][49] = 9'b111111111;
assign micromatr[7][50] = 9'b111111111;
assign micromatr[7][51] = 9'b111111111;
assign micromatr[7][52] = 9'b111111111;
assign micromatr[7][53] = 9'b111111111;
assign micromatr[7][54] = 9'b111111111;
assign micromatr[7][55] = 9'b111111111;
assign micromatr[7][56] = 9'b111111111;
assign micromatr[7][57] = 9'b111111111;
assign micromatr[7][58] = 9'b111111111;
assign micromatr[7][59] = 9'b111111111;
assign micromatr[7][60] = 9'b111111111;
assign micromatr[7][61] = 9'b111111111;
assign micromatr[7][62] = 9'b111111111;
assign micromatr[7][63] = 9'b111111111;
assign micromatr[7][64] = 9'b111111111;
assign micromatr[7][65] = 9'b111111111;
assign micromatr[7][66] = 9'b111111111;
assign micromatr[7][67] = 9'b111111111;
assign micromatr[7][68] = 9'b111111111;
assign micromatr[7][69] = 9'b111111111;
assign micromatr[7][70] = 9'b111111111;
assign micromatr[7][71] = 9'b111111111;
assign micromatr[7][72] = 9'b111111111;
assign micromatr[7][73] = 9'b111111111;
assign micromatr[7][74] = 9'b111111111;
assign micromatr[7][75] = 9'b111111111;
assign micromatr[7][76] = 9'b111111111;
assign micromatr[7][77] = 9'b111111111;
assign micromatr[7][78] = 9'b111111111;
assign micromatr[7][79] = 9'b111111111;
assign micromatr[7][80] = 9'b111111111;
assign micromatr[7][81] = 9'b111111111;
assign micromatr[7][82] = 9'b111111111;
assign micromatr[7][83] = 9'b111111111;
assign micromatr[7][84] = 9'b111111111;
assign micromatr[7][85] = 9'b111111111;
assign micromatr[7][86] = 9'b111111111;
assign micromatr[7][87] = 9'b111111111;
assign micromatr[7][88] = 9'b111111111;
assign micromatr[7][89] = 9'b111111111;
assign micromatr[7][90] = 9'b111111111;
assign micromatr[7][91] = 9'b111111111;
assign micromatr[7][92] = 9'b111111111;
assign micromatr[7][93] = 9'b111111111;
assign micromatr[7][94] = 9'b111111111;
assign micromatr[7][95] = 9'b111111111;
assign micromatr[7][96] = 9'b111111111;
assign micromatr[7][97] = 9'b111111111;
assign micromatr[7][98] = 9'b111111111;
assign micromatr[7][99] = 9'b111111111;
assign micromatr[8][0] = 9'b111111111;
assign micromatr[8][1] = 9'b111111111;
assign micromatr[8][2] = 9'b111111111;
assign micromatr[8][3] = 9'b111111111;
assign micromatr[8][4] = 9'b111111111;
assign micromatr[8][5] = 9'b111111111;
assign micromatr[8][6] = 9'b111111111;
assign micromatr[8][7] = 9'b111111111;
assign micromatr[8][8] = 9'b111111111;
assign micromatr[8][9] = 9'b111111111;
assign micromatr[8][10] = 9'b111111111;
assign micromatr[8][11] = 9'b111111111;
assign micromatr[8][12] = 9'b111111111;
assign micromatr[8][13] = 9'b111111111;
assign micromatr[8][14] = 9'b111111111;
assign micromatr[8][15] = 9'b111111111;
assign micromatr[8][16] = 9'b111111111;
assign micromatr[8][17] = 9'b111111111;
assign micromatr[8][18] = 9'b111111111;
assign micromatr[8][19] = 9'b111111111;
assign micromatr[8][20] = 9'b111111111;
assign micromatr[8][21] = 9'b111111111;
assign micromatr[8][22] = 9'b111111111;
assign micromatr[8][23] = 9'b111111111;
assign micromatr[8][24] = 9'b111111111;
assign micromatr[8][25] = 9'b111111111;
assign micromatr[8][26] = 9'b111111111;
assign micromatr[8][27] = 9'b111111111;
assign micromatr[8][28] = 9'b111111111;
assign micromatr[8][29] = 9'b111111111;
assign micromatr[8][30] = 9'b111111111;
assign micromatr[8][31] = 9'b111111111;
assign micromatr[8][32] = 9'b111111111;
assign micromatr[8][33] = 9'b111111111;
assign micromatr[8][34] = 9'b111111111;
assign micromatr[8][35] = 9'b111111111;
assign micromatr[8][36] = 9'b111111111;
assign micromatr[8][37] = 9'b111111111;
assign micromatr[8][38] = 9'b111111111;
assign micromatr[8][39] = 9'b111111111;
assign micromatr[8][40] = 9'b111111111;
assign micromatr[8][41] = 9'b111111111;
assign micromatr[8][42] = 9'b111111111;
assign micromatr[8][43] = 9'b111111111;
assign micromatr[8][44] = 9'b111111111;
assign micromatr[8][45] = 9'b111111111;
assign micromatr[8][46] = 9'b111111111;
assign micromatr[8][47] = 9'b111111111;
assign micromatr[8][48] = 9'b111111111;
assign micromatr[8][49] = 9'b111111111;
assign micromatr[8][50] = 9'b111111111;
assign micromatr[8][51] = 9'b111111111;
assign micromatr[8][52] = 9'b111111111;
assign micromatr[8][53] = 9'b111111111;
assign micromatr[8][54] = 9'b111111111;
assign micromatr[8][55] = 9'b111111111;
assign micromatr[8][56] = 9'b111111111;
assign micromatr[8][57] = 9'b111111111;
assign micromatr[8][58] = 9'b111111111;
assign micromatr[8][59] = 9'b111111111;
assign micromatr[8][60] = 9'b111111111;
assign micromatr[8][61] = 9'b111111111;
assign micromatr[8][62] = 9'b111111111;
assign micromatr[8][63] = 9'b111111111;
assign micromatr[8][64] = 9'b111111111;
assign micromatr[8][65] = 9'b111111111;
assign micromatr[8][66] = 9'b111111111;
assign micromatr[8][67] = 9'b111111111;
assign micromatr[8][68] = 9'b111111111;
assign micromatr[8][69] = 9'b111111111;
assign micromatr[8][70] = 9'b111111111;
assign micromatr[8][71] = 9'b111111111;
assign micromatr[8][72] = 9'b111111111;
assign micromatr[8][73] = 9'b111111111;
assign micromatr[8][74] = 9'b111111111;
assign micromatr[8][75] = 9'b111111111;
assign micromatr[8][76] = 9'b111111111;
assign micromatr[8][77] = 9'b111111111;
assign micromatr[8][78] = 9'b111111111;
assign micromatr[8][79] = 9'b111111111;
assign micromatr[8][80] = 9'b111111111;
assign micromatr[8][81] = 9'b111111111;
assign micromatr[8][82] = 9'b111111111;
assign micromatr[8][83] = 9'b111111111;
assign micromatr[8][84] = 9'b111111111;
assign micromatr[8][85] = 9'b111111111;
assign micromatr[8][86] = 9'b111111111;
assign micromatr[8][87] = 9'b111111111;
assign micromatr[8][88] = 9'b111111111;
assign micromatr[8][89] = 9'b111111111;
assign micromatr[8][90] = 9'b111111111;
assign micromatr[8][91] = 9'b111111111;
assign micromatr[8][92] = 9'b111111111;
assign micromatr[8][93] = 9'b111111111;
assign micromatr[8][94] = 9'b111111111;
assign micromatr[8][95] = 9'b111111111;
assign micromatr[8][96] = 9'b111111111;
assign micromatr[8][97] = 9'b111111111;
assign micromatr[8][98] = 9'b111111111;
assign micromatr[8][99] = 9'b111111111;
assign micromatr[9][0] = 9'b111111111;
assign micromatr[9][1] = 9'b111111111;
assign micromatr[9][2] = 9'b111111111;
assign micromatr[9][3] = 9'b111111111;
assign micromatr[9][4] = 9'b111111111;
assign micromatr[9][5] = 9'b111111111;
assign micromatr[9][6] = 9'b111111111;
assign micromatr[9][7] = 9'b111111111;
assign micromatr[9][8] = 9'b111111111;
assign micromatr[9][9] = 9'b111111111;
assign micromatr[9][10] = 9'b111111111;
assign micromatr[9][11] = 9'b111111111;
assign micromatr[9][12] = 9'b111111111;
assign micromatr[9][13] = 9'b111111111;
assign micromatr[9][14] = 9'b111111111;
assign micromatr[9][15] = 9'b111111111;
assign micromatr[9][16] = 9'b111111111;
assign micromatr[9][17] = 9'b111111111;
assign micromatr[9][18] = 9'b111111111;
assign micromatr[9][19] = 9'b111111111;
assign micromatr[9][20] = 9'b111111111;
assign micromatr[9][21] = 9'b111111111;
assign micromatr[9][22] = 9'b111111111;
assign micromatr[9][23] = 9'b111111111;
assign micromatr[9][24] = 9'b111111111;
assign micromatr[9][25] = 9'b111111111;
assign micromatr[9][26] = 9'b111111111;
assign micromatr[9][27] = 9'b111111111;
assign micromatr[9][28] = 9'b111111111;
assign micromatr[9][29] = 9'b111111111;
assign micromatr[9][30] = 9'b111111111;
assign micromatr[9][31] = 9'b111111111;
assign micromatr[9][32] = 9'b111111111;
assign micromatr[9][33] = 9'b111111111;
assign micromatr[9][34] = 9'b111111111;
assign micromatr[9][35] = 9'b111111111;
assign micromatr[9][36] = 9'b111111111;
assign micromatr[9][37] = 9'b111111111;
assign micromatr[9][38] = 9'b111111111;
assign micromatr[9][39] = 9'b111111111;
assign micromatr[9][40] = 9'b111111111;
assign micromatr[9][41] = 9'b111111111;
assign micromatr[9][42] = 9'b111111111;
assign micromatr[9][43] = 9'b111111111;
assign micromatr[9][44] = 9'b111111111;
assign micromatr[9][45] = 9'b111111111;
assign micromatr[9][46] = 9'b111111111;
assign micromatr[9][47] = 9'b111111111;
assign micromatr[9][48] = 9'b111111111;
assign micromatr[9][49] = 9'b111111111;
assign micromatr[9][50] = 9'b111111111;
assign micromatr[9][51] = 9'b111111111;
assign micromatr[9][52] = 9'b111111111;
assign micromatr[9][53] = 9'b111111111;
assign micromatr[9][54] = 9'b111111111;
assign micromatr[9][55] = 9'b111111111;
assign micromatr[9][56] = 9'b111111111;
assign micromatr[9][57] = 9'b111111111;
assign micromatr[9][58] = 9'b111111111;
assign micromatr[9][59] = 9'b111111111;
assign micromatr[9][60] = 9'b111111111;
assign micromatr[9][61] = 9'b111111111;
assign micromatr[9][62] = 9'b111111111;
assign micromatr[9][63] = 9'b111111111;
assign micromatr[9][64] = 9'b111111111;
assign micromatr[9][65] = 9'b111111111;
assign micromatr[9][66] = 9'b111111111;
assign micromatr[9][67] = 9'b111111111;
assign micromatr[9][68] = 9'b111111111;
assign micromatr[9][69] = 9'b111111111;
assign micromatr[9][70] = 9'b111111111;
assign micromatr[9][71] = 9'b111111111;
assign micromatr[9][72] = 9'b111111111;
assign micromatr[9][73] = 9'b111111111;
assign micromatr[9][74] = 9'b111111111;
assign micromatr[9][75] = 9'b111111111;
assign micromatr[9][76] = 9'b111111111;
assign micromatr[9][77] = 9'b111111111;
assign micromatr[9][78] = 9'b111111111;
assign micromatr[9][79] = 9'b111111111;
assign micromatr[9][80] = 9'b111111111;
assign micromatr[9][81] = 9'b111111111;
assign micromatr[9][82] = 9'b111111111;
assign micromatr[9][83] = 9'b111111111;
assign micromatr[9][84] = 9'b111111111;
assign micromatr[9][85] = 9'b111111111;
assign micromatr[9][86] = 9'b111111111;
assign micromatr[9][87] = 9'b111111111;
assign micromatr[9][88] = 9'b111111111;
assign micromatr[9][89] = 9'b111111111;
assign micromatr[9][90] = 9'b111111111;
assign micromatr[9][91] = 9'b111111111;
assign micromatr[9][92] = 9'b111111111;
assign micromatr[9][93] = 9'b111111111;
assign micromatr[9][94] = 9'b111111111;
assign micromatr[9][95] = 9'b111111111;
assign micromatr[9][96] = 9'b111111111;
assign micromatr[9][97] = 9'b111111111;
assign micromatr[9][98] = 9'b111111111;
assign micromatr[9][99] = 9'b111111111;
assign micromatr[10][0] = 9'b111111111;
assign micromatr[10][1] = 9'b111111111;
assign micromatr[10][2] = 9'b111111111;
assign micromatr[10][3] = 9'b111111111;
assign micromatr[10][4] = 9'b111111111;
assign micromatr[10][5] = 9'b111111111;
assign micromatr[10][6] = 9'b111111111;
assign micromatr[10][7] = 9'b111111111;
assign micromatr[10][8] = 9'b111111111;
assign micromatr[10][9] = 9'b111111111;
assign micromatr[10][10] = 9'b111111111;
assign micromatr[10][11] = 9'b111111111;
assign micromatr[10][12] = 9'b111111111;
assign micromatr[10][13] = 9'b111111111;
assign micromatr[10][14] = 9'b111111111;
assign micromatr[10][15] = 9'b111111111;
assign micromatr[10][16] = 9'b111111111;
assign micromatr[10][17] = 9'b111111111;
assign micromatr[10][18] = 9'b111111111;
assign micromatr[10][19] = 9'b111111111;
assign micromatr[10][20] = 9'b111111111;
assign micromatr[10][21] = 9'b111111111;
assign micromatr[10][22] = 9'b111111111;
assign micromatr[10][23] = 9'b111111111;
assign micromatr[10][24] = 9'b111111111;
assign micromatr[10][25] = 9'b111111111;
assign micromatr[10][26] = 9'b111111111;
assign micromatr[10][27] = 9'b111111111;
assign micromatr[10][28] = 9'b111111111;
assign micromatr[10][29] = 9'b111111111;
assign micromatr[10][30] = 9'b111111111;
assign micromatr[10][31] = 9'b111111111;
assign micromatr[10][32] = 9'b111111111;
assign micromatr[10][33] = 9'b111111111;
assign micromatr[10][34] = 9'b111111111;
assign micromatr[10][35] = 9'b111111111;
assign micromatr[10][36] = 9'b111111111;
assign micromatr[10][37] = 9'b111111111;
assign micromatr[10][38] = 9'b111111111;
assign micromatr[10][39] = 9'b111111111;
assign micromatr[10][40] = 9'b111111111;
assign micromatr[10][41] = 9'b111111111;
assign micromatr[10][42] = 9'b111111111;
assign micromatr[10][43] = 9'b111111111;
assign micromatr[10][44] = 9'b111111111;
assign micromatr[10][45] = 9'b111111111;
assign micromatr[10][46] = 9'b111111111;
assign micromatr[10][47] = 9'b111111111;
assign micromatr[10][48] = 9'b111111111;
assign micromatr[10][49] = 9'b111111111;
assign micromatr[10][50] = 9'b111111111;
assign micromatr[10][51] = 9'b111111111;
assign micromatr[10][52] = 9'b111111111;
assign micromatr[10][53] = 9'b111111111;
assign micromatr[10][54] = 9'b111111111;
assign micromatr[10][55] = 9'b111111111;
assign micromatr[10][56] = 9'b111111111;
assign micromatr[10][57] = 9'b111111111;
assign micromatr[10][58] = 9'b111111111;
assign micromatr[10][59] = 9'b111111111;
assign micromatr[10][60] = 9'b111111111;
assign micromatr[10][61] = 9'b111111111;
assign micromatr[10][62] = 9'b111111111;
assign micromatr[10][63] = 9'b111111111;
assign micromatr[10][64] = 9'b111111111;
assign micromatr[10][65] = 9'b111111111;
assign micromatr[10][66] = 9'b111111111;
assign micromatr[10][67] = 9'b111111111;
assign micromatr[10][68] = 9'b111111111;
assign micromatr[10][69] = 9'b111111111;
assign micromatr[10][70] = 9'b111111111;
assign micromatr[10][71] = 9'b111111111;
assign micromatr[10][72] = 9'b111111111;
assign micromatr[10][73] = 9'b111111111;
assign micromatr[10][74] = 9'b111111111;
assign micromatr[10][75] = 9'b111111111;
assign micromatr[10][76] = 9'b111111111;
assign micromatr[10][77] = 9'b111111111;
assign micromatr[10][78] = 9'b111111111;
assign micromatr[10][79] = 9'b111111111;
assign micromatr[10][80] = 9'b111111111;
assign micromatr[10][81] = 9'b111111111;
assign micromatr[10][82] = 9'b111111111;
assign micromatr[10][83] = 9'b111111111;
assign micromatr[10][84] = 9'b111111111;
assign micromatr[10][85] = 9'b111111111;
assign micromatr[10][86] = 9'b111111111;
assign micromatr[10][87] = 9'b111111111;
assign micromatr[10][88] = 9'b111111111;
assign micromatr[10][89] = 9'b111111111;
assign micromatr[10][90] = 9'b111111111;
assign micromatr[10][91] = 9'b111111111;
assign micromatr[10][92] = 9'b111111111;
assign micromatr[10][93] = 9'b111111111;
assign micromatr[10][94] = 9'b111111111;
assign micromatr[10][95] = 9'b111111111;
assign micromatr[10][96] = 9'b111111111;
assign micromatr[10][97] = 9'b111111111;
assign micromatr[10][98] = 9'b111111111;
assign micromatr[10][99] = 9'b111111111;
assign micromatr[11][0] = 9'b111111111;
assign micromatr[11][1] = 9'b111111111;
assign micromatr[11][2] = 9'b111111111;
assign micromatr[11][3] = 9'b111111111;
assign micromatr[11][4] = 9'b111111111;
assign micromatr[11][5] = 9'b111111111;
assign micromatr[11][6] = 9'b111111111;
assign micromatr[11][7] = 9'b111111111;
assign micromatr[11][8] = 9'b111111111;
assign micromatr[11][9] = 9'b111111111;
assign micromatr[11][10] = 9'b111111111;
assign micromatr[11][11] = 9'b111111111;
assign micromatr[11][12] = 9'b111111111;
assign micromatr[11][13] = 9'b111111111;
assign micromatr[11][14] = 9'b111111111;
assign micromatr[11][15] = 9'b111111111;
assign micromatr[11][16] = 9'b111111111;
assign micromatr[11][17] = 9'b111111111;
assign micromatr[11][18] = 9'b111111111;
assign micromatr[11][19] = 9'b111111111;
assign micromatr[11][20] = 9'b111111111;
assign micromatr[11][21] = 9'b111111111;
assign micromatr[11][22] = 9'b111111111;
assign micromatr[11][23] = 9'b111111111;
assign micromatr[11][24] = 9'b111111111;
assign micromatr[11][25] = 9'b111111111;
assign micromatr[11][26] = 9'b111111111;
assign micromatr[11][27] = 9'b111111111;
assign micromatr[11][28] = 9'b111111111;
assign micromatr[11][29] = 9'b111111111;
assign micromatr[11][30] = 9'b111111111;
assign micromatr[11][31] = 9'b111111111;
assign micromatr[11][32] = 9'b111111111;
assign micromatr[11][33] = 9'b111111111;
assign micromatr[11][34] = 9'b111111111;
assign micromatr[11][35] = 9'b111111111;
assign micromatr[11][36] = 9'b111111111;
assign micromatr[11][37] = 9'b111111111;
assign micromatr[11][38] = 9'b111111111;
assign micromatr[11][39] = 9'b111111111;
assign micromatr[11][40] = 9'b111111111;
assign micromatr[11][41] = 9'b111111111;
assign micromatr[11][42] = 9'b111111111;
assign micromatr[11][43] = 9'b111111111;
assign micromatr[11][44] = 9'b111111111;
assign micromatr[11][45] = 9'b111111111;
assign micromatr[11][46] = 9'b111111111;
assign micromatr[11][47] = 9'b111111111;
assign micromatr[11][48] = 9'b111111111;
assign micromatr[11][49] = 9'b111111111;
assign micromatr[11][50] = 9'b111111111;
assign micromatr[11][51] = 9'b111111111;
assign micromatr[11][52] = 9'b111111111;
assign micromatr[11][53] = 9'b111111111;
assign micromatr[11][54] = 9'b111111111;
assign micromatr[11][55] = 9'b111111111;
assign micromatr[11][56] = 9'b111111111;
assign micromatr[11][57] = 9'b111111111;
assign micromatr[11][58] = 9'b111111111;
assign micromatr[11][59] = 9'b111111111;
assign micromatr[11][60] = 9'b111111111;
assign micromatr[11][61] = 9'b111111111;
assign micromatr[11][62] = 9'b111111111;
assign micromatr[11][63] = 9'b111111111;
assign micromatr[11][64] = 9'b111111111;
assign micromatr[11][65] = 9'b111111111;
assign micromatr[11][66] = 9'b111111111;
assign micromatr[11][67] = 9'b111111111;
assign micromatr[11][68] = 9'b111111111;
assign micromatr[11][69] = 9'b111111111;
assign micromatr[11][70] = 9'b111111111;
assign micromatr[11][71] = 9'b111111111;
assign micromatr[11][72] = 9'b111111111;
assign micromatr[11][73] = 9'b111111111;
assign micromatr[11][74] = 9'b111111111;
assign micromatr[11][75] = 9'b111111111;
assign micromatr[11][76] = 9'b111111111;
assign micromatr[11][77] = 9'b111111111;
assign micromatr[11][78] = 9'b111111111;
assign micromatr[11][79] = 9'b111111111;
assign micromatr[11][80] = 9'b111111111;
assign micromatr[11][81] = 9'b111111111;
assign micromatr[11][82] = 9'b111111111;
assign micromatr[11][83] = 9'b111111111;
assign micromatr[11][84] = 9'b111111111;
assign micromatr[11][85] = 9'b111111111;
assign micromatr[11][86] = 9'b111111111;
assign micromatr[11][87] = 9'b111111111;
assign micromatr[11][88] = 9'b111111111;
assign micromatr[11][89] = 9'b111111111;
assign micromatr[11][90] = 9'b111111111;
assign micromatr[11][91] = 9'b111111111;
assign micromatr[11][92] = 9'b111111111;
assign micromatr[11][93] = 9'b111111111;
assign micromatr[11][94] = 9'b111111111;
assign micromatr[11][95] = 9'b111111111;
assign micromatr[11][96] = 9'b111111111;
assign micromatr[11][97] = 9'b111111111;
assign micromatr[11][98] = 9'b111111111;
assign micromatr[11][99] = 9'b111111111;
assign micromatr[12][0] = 9'b111111111;
assign micromatr[12][1] = 9'b111111111;
assign micromatr[12][2] = 9'b111111111;
assign micromatr[12][3] = 9'b111111111;
assign micromatr[12][4] = 9'b111111111;
assign micromatr[12][5] = 9'b111111111;
assign micromatr[12][6] = 9'b111111111;
assign micromatr[12][7] = 9'b111111111;
assign micromatr[12][8] = 9'b111111111;
assign micromatr[12][9] = 9'b111111111;
assign micromatr[12][10] = 9'b111111111;
assign micromatr[12][11] = 9'b111111111;
assign micromatr[12][12] = 9'b111111111;
assign micromatr[12][13] = 9'b111111111;
assign micromatr[12][14] = 9'b111111111;
assign micromatr[12][15] = 9'b111111111;
assign micromatr[12][16] = 9'b111111111;
assign micromatr[12][17] = 9'b111111111;
assign micromatr[12][18] = 9'b111111111;
assign micromatr[12][19] = 9'b111111111;
assign micromatr[12][20] = 9'b111111111;
assign micromatr[12][21] = 9'b111111111;
assign micromatr[12][22] = 9'b111111111;
assign micromatr[12][23] = 9'b111111111;
assign micromatr[12][24] = 9'b111111111;
assign micromatr[12][25] = 9'b111111111;
assign micromatr[12][26] = 9'b111111111;
assign micromatr[12][27] = 9'b111111111;
assign micromatr[12][28] = 9'b111111111;
assign micromatr[12][29] = 9'b111111111;
assign micromatr[12][30] = 9'b111111111;
assign micromatr[12][31] = 9'b111111111;
assign micromatr[12][32] = 9'b111111111;
assign micromatr[12][33] = 9'b111111111;
assign micromatr[12][34] = 9'b111111111;
assign micromatr[12][35] = 9'b111111111;
assign micromatr[12][36] = 9'b111111111;
assign micromatr[12][37] = 9'b111111111;
assign micromatr[12][38] = 9'b111111111;
assign micromatr[12][39] = 9'b111111111;
assign micromatr[12][40] = 9'b111111111;
assign micromatr[12][41] = 9'b111111111;
assign micromatr[12][42] = 9'b111111111;
assign micromatr[12][43] = 9'b111111111;
assign micromatr[12][44] = 9'b111111111;
assign micromatr[12][45] = 9'b111111111;
assign micromatr[12][46] = 9'b111111111;
assign micromatr[12][47] = 9'b111111111;
assign micromatr[12][48] = 9'b111111111;
assign micromatr[12][49] = 9'b111111111;
assign micromatr[12][50] = 9'b111111111;
assign micromatr[12][51] = 9'b111111111;
assign micromatr[12][52] = 9'b111111111;
assign micromatr[12][53] = 9'b111111111;
assign micromatr[12][54] = 9'b111111111;
assign micromatr[12][55] = 9'b111111111;
assign micromatr[12][56] = 9'b111111111;
assign micromatr[12][57] = 9'b111111111;
assign micromatr[12][58] = 9'b111111111;
assign micromatr[12][59] = 9'b111111111;
assign micromatr[12][60] = 9'b111111111;
assign micromatr[12][61] = 9'b111111111;
assign micromatr[12][62] = 9'b111111111;
assign micromatr[12][63] = 9'b111111111;
assign micromatr[12][64] = 9'b111111111;
assign micromatr[12][65] = 9'b111111111;
assign micromatr[12][66] = 9'b111111111;
assign micromatr[12][67] = 9'b111111111;
assign micromatr[12][68] = 9'b111111111;
assign micromatr[12][69] = 9'b111111111;
assign micromatr[12][70] = 9'b111111111;
assign micromatr[12][71] = 9'b111111111;
assign micromatr[12][72] = 9'b111111111;
assign micromatr[12][73] = 9'b111111111;
assign micromatr[12][74] = 9'b111111111;
assign micromatr[12][75] = 9'b111111111;
assign micromatr[12][76] = 9'b111111111;
assign micromatr[12][77] = 9'b111111111;
assign micromatr[12][78] = 9'b111111111;
assign micromatr[12][79] = 9'b111111111;
assign micromatr[12][80] = 9'b111111111;
assign micromatr[12][81] = 9'b111111111;
assign micromatr[12][82] = 9'b111111111;
assign micromatr[12][83] = 9'b111111111;
assign micromatr[12][84] = 9'b111111111;
assign micromatr[12][85] = 9'b111111111;
assign micromatr[12][86] = 9'b111111111;
assign micromatr[12][87] = 9'b111111111;
assign micromatr[12][88] = 9'b111111111;
assign micromatr[12][89] = 9'b111111111;
assign micromatr[12][90] = 9'b111111111;
assign micromatr[12][91] = 9'b111111111;
assign micromatr[12][92] = 9'b111111111;
assign micromatr[12][93] = 9'b111111111;
assign micromatr[12][94] = 9'b111111111;
assign micromatr[12][95] = 9'b111111111;
assign micromatr[12][96] = 9'b111111111;
assign micromatr[12][97] = 9'b111111111;
assign micromatr[12][98] = 9'b111111111;
assign micromatr[12][99] = 9'b111111111;
assign micromatr[13][0] = 9'b111111111;
assign micromatr[13][1] = 9'b111111111;
assign micromatr[13][2] = 9'b111111111;
assign micromatr[13][3] = 9'b111111111;
assign micromatr[13][4] = 9'b111111111;
assign micromatr[13][5] = 9'b111111111;
assign micromatr[13][6] = 9'b111111111;
assign micromatr[13][7] = 9'b111111111;
assign micromatr[13][8] = 9'b111111111;
assign micromatr[13][9] = 9'b111111111;
assign micromatr[13][10] = 9'b111111111;
assign micromatr[13][11] = 9'b111111111;
assign micromatr[13][12] = 9'b111111111;
assign micromatr[13][13] = 9'b111111111;
assign micromatr[13][14] = 9'b111111111;
assign micromatr[13][15] = 9'b111111111;
assign micromatr[13][16] = 9'b111111111;
assign micromatr[13][17] = 9'b111111111;
assign micromatr[13][18] = 9'b111111111;
assign micromatr[13][19] = 9'b111111111;
assign micromatr[13][20] = 9'b111111111;
assign micromatr[13][21] = 9'b111111111;
assign micromatr[13][22] = 9'b111111111;
assign micromatr[13][23] = 9'b111111111;
assign micromatr[13][24] = 9'b111111111;
assign micromatr[13][25] = 9'b111111111;
assign micromatr[13][26] = 9'b111111111;
assign micromatr[13][27] = 9'b111111111;
assign micromatr[13][28] = 9'b111111111;
assign micromatr[13][29] = 9'b111111111;
assign micromatr[13][30] = 9'b111111111;
assign micromatr[13][31] = 9'b111111111;
assign micromatr[13][32] = 9'b111111111;
assign micromatr[13][33] = 9'b111111111;
assign micromatr[13][34] = 9'b111111111;
assign micromatr[13][35] = 9'b111111111;
assign micromatr[13][36] = 9'b111111111;
assign micromatr[13][37] = 9'b111111111;
assign micromatr[13][38] = 9'b111111111;
assign micromatr[13][39] = 9'b111111111;
assign micromatr[13][40] = 9'b111111111;
assign micromatr[13][41] = 9'b111111111;
assign micromatr[13][42] = 9'b111111111;
assign micromatr[13][43] = 9'b111111111;
assign micromatr[13][44] = 9'b111111111;
assign micromatr[13][45] = 9'b111111111;
assign micromatr[13][46] = 9'b111111111;
assign micromatr[13][47] = 9'b111111111;
assign micromatr[13][48] = 9'b111111111;
assign micromatr[13][49] = 9'b111111111;
assign micromatr[13][50] = 9'b111111111;
assign micromatr[13][51] = 9'b111111111;
assign micromatr[13][52] = 9'b111111111;
assign micromatr[13][53] = 9'b111111111;
assign micromatr[13][54] = 9'b111111111;
assign micromatr[13][55] = 9'b111111111;
assign micromatr[13][56] = 9'b111111111;
assign micromatr[13][57] = 9'b111111111;
assign micromatr[13][58] = 9'b111111111;
assign micromatr[13][59] = 9'b111111111;
assign micromatr[13][60] = 9'b111111111;
assign micromatr[13][61] = 9'b111111111;
assign micromatr[13][62] = 9'b111111111;
assign micromatr[13][63] = 9'b111111111;
assign micromatr[13][64] = 9'b111111111;
assign micromatr[13][65] = 9'b111111111;
assign micromatr[13][66] = 9'b111111111;
assign micromatr[13][67] = 9'b111111111;
assign micromatr[13][68] = 9'b111111111;
assign micromatr[13][69] = 9'b111111111;
assign micromatr[13][70] = 9'b111111111;
assign micromatr[13][71] = 9'b111111111;
assign micromatr[13][72] = 9'b111111111;
assign micromatr[13][73] = 9'b111111111;
assign micromatr[13][74] = 9'b111111111;
assign micromatr[13][75] = 9'b111111111;
assign micromatr[13][76] = 9'b111111111;
assign micromatr[13][77] = 9'b111111111;
assign micromatr[13][78] = 9'b111111111;
assign micromatr[13][79] = 9'b111111111;
assign micromatr[13][80] = 9'b111111111;
assign micromatr[13][81] = 9'b111111111;
assign micromatr[13][82] = 9'b111111111;
assign micromatr[13][83] = 9'b111111111;
assign micromatr[13][84] = 9'b111111111;
assign micromatr[13][85] = 9'b111111111;
assign micromatr[13][86] = 9'b111111111;
assign micromatr[13][87] = 9'b111111111;
assign micromatr[13][88] = 9'b111111111;
assign micromatr[13][89] = 9'b111111111;
assign micromatr[13][90] = 9'b111111111;
assign micromatr[13][91] = 9'b111111111;
assign micromatr[13][92] = 9'b111111111;
assign micromatr[13][93] = 9'b111111111;
assign micromatr[13][94] = 9'b111111111;
assign micromatr[13][95] = 9'b111111111;
assign micromatr[13][96] = 9'b111111111;
assign micromatr[13][97] = 9'b111111111;
assign micromatr[13][98] = 9'b111111111;
assign micromatr[13][99] = 9'b111111111;
assign micromatr[14][0] = 9'b111111111;
assign micromatr[14][1] = 9'b111111111;
assign micromatr[14][2] = 9'b111111111;
assign micromatr[14][3] = 9'b111111111;
assign micromatr[14][4] = 9'b111111111;
assign micromatr[14][5] = 9'b111111111;
assign micromatr[14][6] = 9'b111111111;
assign micromatr[14][7] = 9'b111111111;
assign micromatr[14][8] = 9'b111111111;
assign micromatr[14][9] = 9'b111111111;
assign micromatr[14][10] = 9'b111111111;
assign micromatr[14][11] = 9'b111111111;
assign micromatr[14][12] = 9'b111111111;
assign micromatr[14][13] = 9'b111111111;
assign micromatr[14][14] = 9'b111111111;
assign micromatr[14][15] = 9'b111111111;
assign micromatr[14][16] = 9'b111111111;
assign micromatr[14][17] = 9'b111111111;
assign micromatr[14][18] = 9'b111111111;
assign micromatr[14][19] = 9'b111111111;
assign micromatr[14][20] = 9'b111111111;
assign micromatr[14][21] = 9'b111111111;
assign micromatr[14][22] = 9'b111111111;
assign micromatr[14][23] = 9'b111111111;
assign micromatr[14][24] = 9'b111111111;
assign micromatr[14][25] = 9'b111111111;
assign micromatr[14][26] = 9'b111111111;
assign micromatr[14][27] = 9'b111111111;
assign micromatr[14][28] = 9'b111111111;
assign micromatr[14][29] = 9'b111111111;
assign micromatr[14][30] = 9'b111111111;
assign micromatr[14][31] = 9'b111111111;
assign micromatr[14][32] = 9'b111111111;
assign micromatr[14][33] = 9'b111111111;
assign micromatr[14][34] = 9'b111111111;
assign micromatr[14][35] = 9'b111111111;
assign micromatr[14][36] = 9'b111111111;
assign micromatr[14][37] = 9'b111111111;
assign micromatr[14][38] = 9'b111111111;
assign micromatr[14][39] = 9'b111111111;
assign micromatr[14][40] = 9'b111111111;
assign micromatr[14][41] = 9'b111111111;
assign micromatr[14][42] = 9'b111111111;
assign micromatr[14][43] = 9'b111111111;
assign micromatr[14][44] = 9'b111111111;
assign micromatr[14][45] = 9'b111111111;
assign micromatr[14][46] = 9'b111111111;
assign micromatr[14][47] = 9'b111111111;
assign micromatr[14][48] = 9'b111111111;
assign micromatr[14][49] = 9'b111111111;
assign micromatr[14][50] = 9'b111111111;
assign micromatr[14][51] = 9'b111111111;
assign micromatr[14][52] = 9'b111111111;
assign micromatr[14][53] = 9'b111111111;
assign micromatr[14][54] = 9'b111111111;
assign micromatr[14][55] = 9'b111111111;
assign micromatr[14][56] = 9'b111111111;
assign micromatr[14][57] = 9'b111111111;
assign micromatr[14][58] = 9'b111111111;
assign micromatr[14][59] = 9'b111111111;
assign micromatr[14][60] = 9'b111111111;
assign micromatr[14][61] = 9'b111111111;
assign micromatr[14][62] = 9'b111111111;
assign micromatr[14][63] = 9'b111111111;
assign micromatr[14][64] = 9'b111111111;
assign micromatr[14][65] = 9'b111111111;
assign micromatr[14][66] = 9'b111111111;
assign micromatr[14][67] = 9'b111111111;
assign micromatr[14][68] = 9'b111111111;
assign micromatr[14][69] = 9'b111111111;
assign micromatr[14][70] = 9'b111111111;
assign micromatr[14][71] = 9'b111111111;
assign micromatr[14][72] = 9'b111111111;
assign micromatr[14][73] = 9'b111111111;
assign micromatr[14][74] = 9'b111111111;
assign micromatr[14][75] = 9'b111111111;
assign micromatr[14][76] = 9'b111111111;
assign micromatr[14][77] = 9'b111111111;
assign micromatr[14][78] = 9'b111111111;
assign micromatr[14][79] = 9'b111111111;
assign micromatr[14][80] = 9'b111111111;
assign micromatr[14][81] = 9'b111111111;
assign micromatr[14][82] = 9'b111111111;
assign micromatr[14][83] = 9'b111111111;
assign micromatr[14][84] = 9'b111111111;
assign micromatr[14][85] = 9'b111111111;
assign micromatr[14][86] = 9'b111111111;
assign micromatr[14][87] = 9'b111111111;
assign micromatr[14][88] = 9'b111111111;
assign micromatr[14][89] = 9'b111111111;
assign micromatr[14][90] = 9'b111111111;
assign micromatr[14][91] = 9'b111111111;
assign micromatr[14][92] = 9'b111111111;
assign micromatr[14][93] = 9'b111111111;
assign micromatr[14][94] = 9'b111111111;
assign micromatr[14][95] = 9'b111111111;
assign micromatr[14][96] = 9'b111111111;
assign micromatr[14][97] = 9'b111111111;
assign micromatr[14][98] = 9'b111111111;
assign micromatr[14][99] = 9'b111111111;
assign micromatr[15][0] = 9'b111111111;
assign micromatr[15][1] = 9'b111111111;
assign micromatr[15][2] = 9'b111111111;
assign micromatr[15][3] = 9'b111111111;
assign micromatr[15][4] = 9'b111111111;
assign micromatr[15][5] = 9'b111111111;
assign micromatr[15][6] = 9'b111111111;
assign micromatr[15][7] = 9'b111111111;
assign micromatr[15][8] = 9'b111111111;
assign micromatr[15][9] = 9'b111111111;
assign micromatr[15][10] = 9'b111111111;
assign micromatr[15][11] = 9'b111111111;
assign micromatr[15][12] = 9'b111111111;
assign micromatr[15][13] = 9'b111111111;
assign micromatr[15][14] = 9'b111111111;
assign micromatr[15][15] = 9'b111111111;
assign micromatr[15][16] = 9'b111111111;
assign micromatr[15][17] = 9'b111111111;
assign micromatr[15][18] = 9'b110110110;
assign micromatr[15][19] = 9'b110110110;
assign micromatr[15][20] = 9'b110110010;
assign micromatr[15][21] = 9'b110110110;
assign micromatr[15][22] = 9'b111111111;
assign micromatr[15][23] = 9'b111111111;
assign micromatr[15][24] = 9'b111111111;
assign micromatr[15][25] = 9'b111111111;
assign micromatr[15][26] = 9'b111111111;
assign micromatr[15][27] = 9'b111111111;
assign micromatr[15][28] = 9'b111111111;
assign micromatr[15][29] = 9'b111111111;
assign micromatr[15][30] = 9'b111111111;
assign micromatr[15][31] = 9'b111111111;
assign micromatr[15][32] = 9'b111111111;
assign micromatr[15][33] = 9'b110010001;
assign micromatr[15][34] = 9'b110001110;
assign micromatr[15][35] = 9'b110010001;
assign micromatr[15][36] = 9'b110010010;
assign micromatr[15][37] = 9'b111111111;
assign micromatr[15][38] = 9'b111111111;
assign micromatr[15][39] = 9'b111111111;
assign micromatr[15][40] = 9'b111111111;
assign micromatr[15][41] = 9'b111111111;
assign micromatr[15][42] = 9'b111111111;
assign micromatr[15][43] = 9'b111111111;
assign micromatr[15][44] = 9'b111111111;
assign micromatr[15][45] = 9'b110110110;
assign micromatr[15][46] = 9'b110010010;
assign micromatr[15][47] = 9'b110111111;
assign micromatr[15][48] = 9'b110011111;
assign micromatr[15][49] = 9'b110010001;
assign micromatr[15][50] = 9'b111111111;
assign micromatr[15][51] = 9'b111111111;
assign micromatr[15][52] = 9'b111111111;
assign micromatr[15][53] = 9'b111111111;
assign micromatr[15][54] = 9'b111111111;
assign micromatr[15][55] = 9'b111111111;
assign micromatr[15][56] = 9'b111111111;
assign micromatr[15][57] = 9'b111111111;
assign micromatr[15][58] = 9'b111111111;
assign micromatr[15][59] = 9'b111111111;
assign micromatr[15][60] = 9'b111111111;
assign micromatr[15][61] = 9'b111111111;
assign micromatr[15][62] = 9'b111111111;
assign micromatr[15][63] = 9'b111111111;
assign micromatr[15][64] = 9'b111111111;
assign micromatr[15][65] = 9'b111111111;
assign micromatr[15][66] = 9'b110001101;
assign micromatr[15][67] = 9'b110010010;
assign micromatr[15][68] = 9'b110110011;
assign micromatr[15][69] = 9'b110001110;
assign micromatr[15][70] = 9'b110110110;
assign micromatr[15][71] = 9'b111111111;
assign micromatr[15][72] = 9'b111111111;
assign micromatr[15][73] = 9'b111111111;
assign micromatr[15][74] = 9'b111111111;
assign micromatr[15][75] = 9'b111111111;
assign micromatr[15][76] = 9'b111111111;
assign micromatr[15][77] = 9'b111111111;
assign micromatr[15][78] = 9'b111111111;
assign micromatr[15][79] = 9'b111111111;
assign micromatr[15][80] = 9'b111111111;
assign micromatr[15][81] = 9'b111111111;
assign micromatr[15][82] = 9'b111111111;
assign micromatr[15][83] = 9'b111111111;
assign micromatr[15][84] = 9'b111111111;
assign micromatr[15][85] = 9'b111111111;
assign micromatr[15][86] = 9'b111111111;
assign micromatr[15][87] = 9'b111111111;
assign micromatr[15][88] = 9'b111111111;
assign micromatr[15][89] = 9'b111111111;
assign micromatr[15][90] = 9'b111111111;
assign micromatr[15][91] = 9'b111111111;
assign micromatr[15][92] = 9'b111111111;
assign micromatr[15][93] = 9'b111111111;
assign micromatr[15][94] = 9'b111111111;
assign micromatr[15][95] = 9'b111111111;
assign micromatr[15][96] = 9'b111111111;
assign micromatr[15][97] = 9'b111111111;
assign micromatr[15][98] = 9'b111111111;
assign micromatr[15][99] = 9'b111111111;
assign micromatr[16][0] = 9'b111111111;
assign micromatr[16][1] = 9'b111111111;
assign micromatr[16][2] = 9'b111111111;
assign micromatr[16][3] = 9'b111111111;
assign micromatr[16][4] = 9'b111111111;
assign micromatr[16][5] = 9'b111111111;
assign micromatr[16][6] = 9'b111111111;
assign micromatr[16][7] = 9'b111111111;
assign micromatr[16][8] = 9'b111111111;
assign micromatr[16][9] = 9'b111111111;
assign micromatr[16][10] = 9'b111111111;
assign micromatr[16][11] = 9'b111111111;
assign micromatr[16][12] = 9'b111111111;
assign micromatr[16][13] = 9'b111111111;
assign micromatr[16][14] = 9'b111111111;
assign micromatr[16][15] = 9'b110110010;
assign micromatr[16][16] = 9'b110110010;
assign micromatr[16][17] = 9'b111110010;
assign micromatr[16][18] = 9'b111110010;
assign micromatr[16][19] = 9'b111110011;
assign micromatr[16][20] = 9'b111110011;
assign micromatr[16][21] = 9'b110001101;
assign micromatr[16][22] = 9'b111111111;
assign micromatr[16][23] = 9'b111111111;
assign micromatr[16][24] = 9'b111111111;
assign micromatr[16][25] = 9'b111111111;
assign micromatr[16][26] = 9'b111111111;
assign micromatr[16][27] = 9'b111111111;
assign micromatr[16][28] = 9'b111111111;
assign micromatr[16][29] = 9'b111111111;
assign micromatr[16][30] = 9'b111111111;
assign micromatr[16][31] = 9'b111111111;
assign micromatr[16][32] = 9'b111111111;
assign micromatr[16][33] = 9'b110001110;
assign micromatr[16][34] = 9'b111111111;
assign micromatr[16][35] = 9'b111110111;
assign micromatr[16][36] = 9'b111110011;
assign micromatr[16][37] = 9'b110001110;
assign micromatr[16][38] = 9'b110010010;
assign micromatr[16][39] = 9'b111111111;
assign micromatr[16][40] = 9'b111111111;
assign micromatr[16][41] = 9'b111111111;
assign micromatr[16][42] = 9'b111111111;
assign micromatr[16][43] = 9'b111111111;
assign micromatr[16][44] = 9'b111111111;
assign micromatr[16][45] = 9'b110010010;
assign micromatr[16][46] = 9'b111111111;
assign micromatr[16][47] = 9'b111111111;
assign micromatr[16][48] = 9'b111111111;
assign micromatr[16][49] = 9'b111111111;
assign micromatr[16][50] = 9'b110010001;
assign micromatr[16][51] = 9'b111111111;
assign micromatr[16][52] = 9'b110110110;
assign micromatr[16][53] = 9'b110001101;
assign micromatr[16][54] = 9'b111110010;
assign micromatr[16][55] = 9'b111110010;
assign micromatr[16][56] = 9'b111110010;
assign micromatr[16][57] = 9'b111110010;
assign micromatr[16][58] = 9'b110001101;
assign micromatr[16][59] = 9'b111111111;
assign micromatr[16][60] = 9'b111111111;
assign micromatr[16][61] = 9'b111111111;
assign micromatr[16][62] = 9'b111111111;
assign micromatr[16][63] = 9'b111111111;
assign micromatr[16][64] = 9'b111111111;
assign micromatr[16][65] = 9'b110001101;
assign micromatr[16][66] = 9'b111110011;
assign micromatr[16][67] = 9'b111110111;
assign micromatr[16][68] = 9'b111110111;
assign micromatr[16][69] = 9'b111110111;
assign micromatr[16][70] = 9'b110001110;
assign micromatr[16][71] = 9'b110110110;
assign micromatr[16][72] = 9'b111111111;
assign micromatr[16][73] = 9'b110110110;
assign micromatr[16][74] = 9'b110010110;
assign micromatr[16][75] = 9'b110010010;
assign micromatr[16][76] = 9'b110010110;
assign micromatr[16][77] = 9'b110010010;
assign micromatr[16][78] = 9'b110010110;
assign micromatr[16][79] = 9'b110010110;
assign micromatr[16][80] = 9'b110010110;
assign micromatr[16][81] = 9'b110011111;
assign micromatr[16][82] = 9'b110010111;
assign micromatr[16][83] = 9'b110010010;
assign micromatr[16][84] = 9'b111111111;
assign micromatr[16][85] = 9'b111111111;
assign micromatr[16][86] = 9'b111111111;
assign micromatr[16][87] = 9'b111111111;
assign micromatr[16][88] = 9'b111111111;
assign micromatr[16][89] = 9'b111111111;
assign micromatr[16][90] = 9'b111111111;
assign micromatr[16][91] = 9'b111111111;
assign micromatr[16][92] = 9'b111111111;
assign micromatr[16][93] = 9'b111111111;
assign micromatr[16][94] = 9'b111111111;
assign micromatr[16][95] = 9'b111111111;
assign micromatr[16][96] = 9'b111111111;
assign micromatr[16][97] = 9'b111111111;
assign micromatr[16][98] = 9'b111111111;
assign micromatr[16][99] = 9'b111111111;
assign micromatr[17][0] = 9'b111111111;
assign micromatr[17][1] = 9'b111111111;
assign micromatr[17][2] = 9'b111111111;
assign micromatr[17][3] = 9'b111111111;
assign micromatr[17][4] = 9'b111111111;
assign micromatr[17][5] = 9'b111111111;
assign micromatr[17][6] = 9'b111111111;
assign micromatr[17][7] = 9'b111111111;
assign micromatr[17][8] = 9'b111111111;
assign micromatr[17][9] = 9'b111111111;
assign micromatr[17][10] = 9'b111111111;
assign micromatr[17][11] = 9'b111111111;
assign micromatr[17][12] = 9'b111111111;
assign micromatr[17][13] = 9'b111111111;
assign micromatr[17][14] = 9'b111111111;
assign micromatr[17][15] = 9'b110110010;
assign micromatr[17][16] = 9'b111110111;
assign micromatr[17][17] = 9'b111111111;
assign micromatr[17][18] = 9'b111110111;
assign micromatr[17][19] = 9'b111110111;
assign micromatr[17][20] = 9'b111111111;
assign micromatr[17][21] = 9'b110010001;
assign micromatr[17][22] = 9'b110001101;
assign micromatr[17][23] = 9'b110010001;
assign micromatr[17][24] = 9'b110110010;
assign micromatr[17][25] = 9'b110110010;
assign micromatr[17][26] = 9'b110001101;
assign micromatr[17][27] = 9'b111111111;
assign micromatr[17][28] = 9'b111111111;
assign micromatr[17][29] = 9'b111111111;
assign micromatr[17][30] = 9'b111111111;
assign micromatr[17][31] = 9'b111111111;
assign micromatr[17][32] = 9'b110010010;
assign micromatr[17][33] = 9'b111110011;
assign micromatr[17][34] = 9'b111110111;
assign micromatr[17][35] = 9'b111110111;
assign micromatr[17][36] = 9'b111110111;
assign micromatr[17][37] = 9'b111111111;
assign micromatr[17][38] = 9'b110001101;
assign micromatr[17][39] = 9'b110110110;
assign micromatr[17][40] = 9'b111111111;
assign micromatr[17][41] = 9'b111111111;
assign micromatr[17][42] = 9'b111111111;
assign micromatr[17][43] = 9'b111111111;
assign micromatr[17][44] = 9'b110010110;
assign micromatr[17][45] = 9'b111111111;
assign micromatr[17][46] = 9'b111111111;
assign micromatr[17][47] = 9'b111111111;
assign micromatr[17][48] = 9'b111111111;
assign micromatr[17][49] = 9'b111111111;
assign micromatr[17][50] = 9'b110010110;
assign micromatr[17][51] = 9'b110010110;
assign micromatr[17][52] = 9'b110110010;
assign micromatr[17][53] = 9'b111110111;
assign micromatr[17][54] = 9'b111111111;
assign micromatr[17][55] = 9'b111111111;
assign micromatr[17][56] = 9'b111111111;
assign micromatr[17][57] = 9'b111111111;
assign micromatr[17][58] = 9'b110001101;
assign micromatr[17][59] = 9'b111110110;
assign micromatr[17][60] = 9'b111111111;
assign micromatr[17][61] = 9'b111111111;
assign micromatr[17][62] = 9'b111111111;
assign micromatr[17][63] = 9'b111111111;
assign micromatr[17][64] = 9'b111111111;
assign micromatr[17][65] = 9'b110010010;
assign micromatr[17][66] = 9'b111110111;
assign micromatr[17][67] = 9'b111110111;
assign micromatr[17][68] = 9'b111110111;
assign micromatr[17][69] = 9'b111110111;
assign micromatr[17][70] = 9'b111110011;
assign micromatr[17][71] = 9'b110001101;
assign micromatr[17][72] = 9'b111111111;
assign micromatr[17][73] = 9'b110010010;
assign micromatr[17][74] = 9'b111111111;
assign micromatr[17][75] = 9'b111111111;
assign micromatr[17][76] = 9'b111111111;
assign micromatr[17][77] = 9'b111111111;
assign micromatr[17][78] = 9'b111111111;
assign micromatr[17][79] = 9'b111111111;
assign micromatr[17][80] = 9'b111111111;
assign micromatr[17][81] = 9'b111111111;
assign micromatr[17][82] = 9'b111111111;
assign micromatr[17][83] = 9'b110010001;
assign micromatr[17][84] = 9'b111111111;
assign micromatr[17][85] = 9'b111111111;
assign micromatr[17][86] = 9'b111111111;
assign micromatr[17][87] = 9'b111111111;
assign micromatr[17][88] = 9'b111111111;
assign micromatr[17][89] = 9'b111111111;
assign micromatr[17][90] = 9'b111111111;
assign micromatr[17][91] = 9'b111111111;
assign micromatr[17][92] = 9'b111111111;
assign micromatr[17][93] = 9'b111111111;
assign micromatr[17][94] = 9'b111111111;
assign micromatr[17][95] = 9'b111111111;
assign micromatr[17][96] = 9'b111111111;
assign micromatr[17][97] = 9'b111111111;
assign micromatr[17][98] = 9'b111111111;
assign micromatr[17][99] = 9'b111111111;
assign micromatr[18][0] = 9'b111111111;
assign micromatr[18][1] = 9'b111111111;
assign micromatr[18][2] = 9'b111111111;
assign micromatr[18][3] = 9'b111111111;
assign micromatr[18][4] = 9'b111111111;
assign micromatr[18][5] = 9'b111111111;
assign micromatr[18][6] = 9'b111111111;
assign micromatr[18][7] = 9'b111111111;
assign micromatr[18][8] = 9'b111111111;
assign micromatr[18][9] = 9'b111111111;
assign micromatr[18][10] = 9'b111111111;
assign micromatr[18][11] = 9'b111111111;
assign micromatr[18][12] = 9'b111111111;
assign micromatr[18][13] = 9'b111111111;
assign micromatr[18][14] = 9'b111111111;
assign micromatr[18][15] = 9'b110010010;
assign micromatr[18][16] = 9'b111110111;
assign micromatr[18][17] = 9'b111110111;
assign micromatr[18][18] = 9'b111110111;
assign micromatr[18][19] = 9'b111110111;
assign micromatr[18][20] = 9'b111110111;
assign micromatr[18][21] = 9'b110001101;
assign micromatr[18][22] = 9'b110001101;
assign micromatr[18][23] = 9'b111110111;
assign micromatr[18][24] = 9'b111110111;
assign micromatr[18][25] = 9'b111110111;
assign micromatr[18][26] = 9'b111110011;
assign micromatr[18][27] = 9'b110010001;
assign micromatr[18][28] = 9'b111111111;
assign micromatr[18][29] = 9'b111111111;
assign micromatr[18][30] = 9'b111111111;
assign micromatr[18][31] = 9'b111111111;
assign micromatr[18][32] = 9'b110001110;
assign micromatr[18][33] = 9'b111110111;
assign micromatr[18][34] = 9'b111110111;
assign micromatr[18][35] = 9'b111110111;
assign micromatr[18][36] = 9'b111110111;
assign micromatr[18][37] = 9'b111110111;
assign micromatr[18][38] = 9'b111110011;
assign micromatr[18][39] = 9'b101101101;
assign micromatr[18][40] = 9'b111111111;
assign micromatr[18][41] = 9'b111111111;
assign micromatr[18][42] = 9'b111111111;
assign micromatr[18][43] = 9'b111111111;
assign micromatr[18][44] = 9'b110010110;
assign micromatr[18][45] = 9'b111111111;
assign micromatr[18][46] = 9'b111111111;
assign micromatr[18][47] = 9'b111111111;
assign micromatr[18][48] = 9'b111111111;
assign micromatr[18][49] = 9'b111111111;
assign micromatr[18][50] = 9'b110111111;
assign micromatr[18][51] = 9'b110111111;
assign micromatr[18][52] = 9'b110010001;
assign micromatr[18][53] = 9'b111110011;
assign micromatr[18][54] = 9'b111110111;
assign micromatr[18][55] = 9'b111110111;
assign micromatr[18][56] = 9'b111110111;
assign micromatr[18][57] = 9'b111110111;
assign micromatr[18][58] = 9'b110010001;
assign micromatr[18][59] = 9'b111111111;
assign micromatr[18][60] = 9'b111111111;
assign micromatr[18][61] = 9'b111111111;
assign micromatr[18][62] = 9'b111111111;
assign micromatr[18][63] = 9'b111111111;
assign micromatr[18][64] = 9'b111111111;
assign micromatr[18][65] = 9'b110010010;
assign micromatr[18][66] = 9'b111110111;
assign micromatr[18][67] = 9'b111110111;
assign micromatr[18][68] = 9'b111110111;
assign micromatr[18][69] = 9'b111110111;
assign micromatr[18][70] = 9'b111110011;
assign micromatr[18][71] = 9'b110010010;
assign micromatr[18][72] = 9'b110110111;
assign micromatr[18][73] = 9'b110010110;
assign micromatr[18][74] = 9'b111111111;
assign micromatr[18][75] = 9'b111111111;
assign micromatr[18][76] = 9'b111111111;
assign micromatr[18][77] = 9'b111111111;
assign micromatr[18][78] = 9'b111111111;
assign micromatr[18][79] = 9'b111111111;
assign micromatr[18][80] = 9'b111111111;
assign micromatr[18][81] = 9'b111111111;
assign micromatr[18][82] = 9'b111111111;
assign micromatr[18][83] = 9'b110010110;
assign micromatr[18][84] = 9'b111111111;
assign micromatr[18][85] = 9'b111111111;
assign micromatr[18][86] = 9'b111111111;
assign micromatr[18][87] = 9'b111111111;
assign micromatr[18][88] = 9'b111111111;
assign micromatr[18][89] = 9'b111111111;
assign micromatr[18][90] = 9'b111111111;
assign micromatr[18][91] = 9'b111111111;
assign micromatr[18][92] = 9'b111111111;
assign micromatr[18][93] = 9'b111111111;
assign micromatr[18][94] = 9'b111111111;
assign micromatr[18][95] = 9'b111111111;
assign micromatr[18][96] = 9'b111111111;
assign micromatr[18][97] = 9'b111111111;
assign micromatr[18][98] = 9'b111111111;
assign micromatr[18][99] = 9'b111111111;
assign micromatr[19][0] = 9'b111111111;
assign micromatr[19][1] = 9'b111111111;
assign micromatr[19][2] = 9'b111111111;
assign micromatr[19][3] = 9'b111111111;
assign micromatr[19][4] = 9'b111111111;
assign micromatr[19][5] = 9'b111111111;
assign micromatr[19][6] = 9'b111111111;
assign micromatr[19][7] = 9'b111111111;
assign micromatr[19][8] = 9'b111111111;
assign micromatr[19][9] = 9'b111111111;
assign micromatr[19][10] = 9'b111111111;
assign micromatr[19][11] = 9'b111111111;
assign micromatr[19][12] = 9'b111111111;
assign micromatr[19][13] = 9'b111111111;
assign micromatr[19][14] = 9'b111111111;
assign micromatr[19][15] = 9'b110010010;
assign micromatr[19][16] = 9'b111110111;
assign micromatr[19][17] = 9'b111110111;
assign micromatr[19][18] = 9'b111110111;
assign micromatr[19][19] = 9'b111110111;
assign micromatr[19][20] = 9'b111110111;
assign micromatr[19][21] = 9'b110001101;
assign micromatr[19][22] = 9'b110010001;
assign micromatr[19][23] = 9'b111111111;
assign micromatr[19][24] = 9'b111110111;
assign micromatr[19][25] = 9'b111110111;
assign micromatr[19][26] = 9'b111110011;
assign micromatr[19][27] = 9'b110010010;
assign micromatr[19][28] = 9'b111111111;
assign micromatr[19][29] = 9'b111111111;
assign micromatr[19][30] = 9'b111111111;
assign micromatr[19][31] = 9'b111111111;
assign micromatr[19][32] = 9'b110010010;
assign micromatr[19][33] = 9'b111110111;
assign micromatr[19][34] = 9'b111110111;
assign micromatr[19][35] = 9'b111110111;
assign micromatr[19][36] = 9'b111110111;
assign micromatr[19][37] = 9'b111110111;
assign micromatr[19][38] = 9'b111110111;
assign micromatr[19][39] = 9'b110001101;
assign micromatr[19][40] = 9'b110110110;
assign micromatr[19][41] = 9'b111111111;
assign micromatr[19][42] = 9'b111111111;
assign micromatr[19][43] = 9'b111111111;
assign micromatr[19][44] = 9'b111111111;
assign micromatr[19][45] = 9'b110011111;
assign micromatr[19][46] = 9'b111111111;
assign micromatr[19][47] = 9'b111111111;
assign micromatr[19][48] = 9'b111111111;
assign micromatr[19][49] = 9'b111111111;
assign micromatr[19][50] = 9'b110010010;
assign micromatr[19][51] = 9'b111111111;
assign micromatr[19][52] = 9'b110010001;
assign micromatr[19][53] = 9'b111110011;
assign micromatr[19][54] = 9'b111110111;
assign micromatr[19][55] = 9'b111110111;
assign micromatr[19][56] = 9'b111110111;
assign micromatr[19][57] = 9'b111110111;
assign micromatr[19][58] = 9'b110010001;
assign micromatr[19][59] = 9'b111111111;
assign micromatr[19][60] = 9'b111111111;
assign micromatr[19][61] = 9'b111111111;
assign micromatr[19][62] = 9'b111111111;
assign micromatr[19][63] = 9'b111111111;
assign micromatr[19][64] = 9'b111111111;
assign micromatr[19][65] = 9'b110010010;
assign micromatr[19][66] = 9'b111110111;
assign micromatr[19][67] = 9'b111110111;
assign micromatr[19][68] = 9'b111110111;
assign micromatr[19][69] = 9'b111110111;
assign micromatr[19][70] = 9'b110010010;
assign micromatr[19][71] = 9'b111110111;
assign micromatr[19][72] = 9'b111110111;
assign micromatr[19][73] = 9'b110010010;
assign micromatr[19][74] = 9'b111111111;
assign micromatr[19][75] = 9'b111111111;
assign micromatr[19][76] = 9'b111111111;
assign micromatr[19][77] = 9'b111111111;
assign micromatr[19][78] = 9'b111111111;
assign micromatr[19][79] = 9'b111111111;
assign micromatr[19][80] = 9'b111111111;
assign micromatr[19][81] = 9'b111111111;
assign micromatr[19][82] = 9'b111111111;
assign micromatr[19][83] = 9'b110010110;
assign micromatr[19][84] = 9'b111111111;
assign micromatr[19][85] = 9'b111111111;
assign micromatr[19][86] = 9'b111111111;
assign micromatr[19][87] = 9'b111111111;
assign micromatr[19][88] = 9'b111111111;
assign micromatr[19][89] = 9'b111111111;
assign micromatr[19][90] = 9'b111111111;
assign micromatr[19][91] = 9'b111111111;
assign micromatr[19][92] = 9'b111111111;
assign micromatr[19][93] = 9'b111111111;
assign micromatr[19][94] = 9'b111111111;
assign micromatr[19][95] = 9'b111111111;
assign micromatr[19][96] = 9'b111111111;
assign micromatr[19][97] = 9'b111111111;
assign micromatr[19][98] = 9'b111111111;
assign micromatr[19][99] = 9'b111111111;
assign micromatr[20][0] = 9'b111111111;
assign micromatr[20][1] = 9'b111111111;
assign micromatr[20][2] = 9'b111111111;
assign micromatr[20][3] = 9'b111111111;
assign micromatr[20][4] = 9'b111111111;
assign micromatr[20][5] = 9'b111111111;
assign micromatr[20][6] = 9'b111111111;
assign micromatr[20][7] = 9'b111111111;
assign micromatr[20][8] = 9'b111111111;
assign micromatr[20][9] = 9'b111111111;
assign micromatr[20][10] = 9'b111111111;
assign micromatr[20][11] = 9'b111111111;
assign micromatr[20][12] = 9'b111111111;
assign micromatr[20][13] = 9'b111111111;
assign micromatr[20][14] = 9'b111111111;
assign micromatr[20][15] = 9'b110110010;
assign micromatr[20][16] = 9'b111110111;
assign micromatr[20][17] = 9'b111110111;
assign micromatr[20][18] = 9'b111110111;
assign micromatr[20][19] = 9'b111110111;
assign micromatr[20][20] = 9'b111110111;
assign micromatr[20][21] = 9'b110001101;
assign micromatr[20][22] = 9'b110110010;
assign micromatr[20][23] = 9'b111111111;
assign micromatr[20][24] = 9'b111110111;
assign micromatr[20][25] = 9'b111110111;
assign micromatr[20][26] = 9'b111110011;
assign micromatr[20][27] = 9'b110110010;
assign micromatr[20][28] = 9'b111111111;
assign micromatr[20][29] = 9'b111111111;
assign micromatr[20][30] = 9'b111111111;
assign micromatr[20][31] = 9'b110010010;
assign micromatr[20][32] = 9'b111110011;
assign micromatr[20][33] = 9'b111110111;
assign micromatr[20][34] = 9'b111110111;
assign micromatr[20][35] = 9'b111110111;
assign micromatr[20][36] = 9'b111110111;
assign micromatr[20][37] = 9'b111110111;
assign micromatr[20][38] = 9'b111110111;
assign micromatr[20][39] = 9'b110110011;
assign micromatr[20][40] = 9'b110001101;
assign micromatr[20][41] = 9'b111111111;
assign micromatr[20][42] = 9'b111111111;
assign micromatr[20][43] = 9'b111111111;
assign micromatr[20][44] = 9'b111111111;
assign micromatr[20][45] = 9'b101101101;
assign micromatr[20][46] = 9'b110011111;
assign micromatr[20][47] = 9'b111111111;
assign micromatr[20][48] = 9'b111111111;
assign micromatr[20][49] = 9'b110010111;
assign micromatr[20][50] = 9'b101101101;
assign micromatr[20][51] = 9'b111111111;
assign micromatr[20][52] = 9'b110010001;
assign micromatr[20][53] = 9'b111110011;
assign micromatr[20][54] = 9'b111110111;
assign micromatr[20][55] = 9'b111110111;
assign micromatr[20][56] = 9'b111110111;
assign micromatr[20][57] = 9'b111110111;
assign micromatr[20][58] = 9'b110010001;
assign micromatr[20][59] = 9'b111111111;
assign micromatr[20][60] = 9'b111111111;
assign micromatr[20][61] = 9'b111111111;
assign micromatr[20][62] = 9'b111111111;
assign micromatr[20][63] = 9'b111111111;
assign micromatr[20][64] = 9'b111111111;
assign micromatr[20][65] = 9'b110010001;
assign micromatr[20][66] = 9'b101101101;
assign micromatr[20][67] = 9'b111110111;
assign micromatr[20][68] = 9'b111110111;
assign micromatr[20][69] = 9'b111110011;
assign micromatr[20][70] = 9'b101101001;
assign micromatr[20][71] = 9'b110110011;
assign micromatr[20][72] = 9'b111110111;
assign micromatr[20][73] = 9'b110010110;
assign micromatr[20][74] = 9'b111111111;
assign micromatr[20][75] = 9'b111111111;
assign micromatr[20][76] = 9'b111111111;
assign micromatr[20][77] = 9'b111111111;
assign micromatr[20][78] = 9'b111111111;
assign micromatr[20][79] = 9'b111111111;
assign micromatr[20][80] = 9'b111111111;
assign micromatr[20][81] = 9'b111111111;
assign micromatr[20][82] = 9'b111111111;
assign micromatr[20][83] = 9'b110010110;
assign micromatr[20][84] = 9'b111111111;
assign micromatr[20][85] = 9'b111111111;
assign micromatr[20][86] = 9'b111111111;
assign micromatr[20][87] = 9'b111111111;
assign micromatr[20][88] = 9'b111111111;
assign micromatr[20][89] = 9'b111111111;
assign micromatr[20][90] = 9'b111111111;
assign micromatr[20][91] = 9'b111111111;
assign micromatr[20][92] = 9'b111111111;
assign micromatr[20][93] = 9'b111111111;
assign micromatr[20][94] = 9'b111111111;
assign micromatr[20][95] = 9'b111111111;
assign micromatr[20][96] = 9'b111111111;
assign micromatr[20][97] = 9'b111111111;
assign micromatr[20][98] = 9'b111111111;
assign micromatr[20][99] = 9'b111111111;
assign micromatr[21][0] = 9'b111111111;
assign micromatr[21][1] = 9'b111111111;
assign micromatr[21][2] = 9'b111111111;
assign micromatr[21][3] = 9'b111111111;
assign micromatr[21][4] = 9'b111111111;
assign micromatr[21][5] = 9'b111111111;
assign micromatr[21][6] = 9'b111111111;
assign micromatr[21][7] = 9'b111111111;
assign micromatr[21][8] = 9'b111111111;
assign micromatr[21][9] = 9'b111111111;
assign micromatr[21][10] = 9'b111111111;
assign micromatr[21][11] = 9'b111111111;
assign micromatr[21][12] = 9'b111111111;
assign micromatr[21][13] = 9'b111111111;
assign micromatr[21][14] = 9'b111111111;
assign micromatr[21][15] = 9'b110110010;
assign micromatr[21][16] = 9'b111110111;
assign micromatr[21][17] = 9'b111110111;
assign micromatr[21][18] = 9'b111110111;
assign micromatr[21][19] = 9'b111110111;
assign micromatr[21][20] = 9'b111110111;
assign micromatr[21][21] = 9'b110001101;
assign micromatr[21][22] = 9'b110110010;
assign micromatr[21][23] = 9'b111111111;
assign micromatr[21][24] = 9'b111110111;
assign micromatr[21][25] = 9'b111110111;
assign micromatr[21][26] = 9'b111110011;
assign micromatr[21][27] = 9'b110110010;
assign micromatr[21][28] = 9'b111111111;
assign micromatr[21][29] = 9'b111111111;
assign micromatr[21][30] = 9'b111111111;
assign micromatr[21][31] = 9'b110001110;
assign micromatr[21][32] = 9'b111110111;
assign micromatr[21][33] = 9'b111110111;
assign micromatr[21][34] = 9'b111110111;
assign micromatr[21][35] = 9'b111110111;
assign micromatr[21][36] = 9'b111110111;
assign micromatr[21][37] = 9'b111110111;
assign micromatr[21][38] = 9'b111110111;
assign micromatr[21][39] = 9'b111110111;
assign micromatr[21][40] = 9'b110001101;
assign micromatr[21][41] = 9'b110110110;
assign micromatr[21][42] = 9'b111111111;
assign micromatr[21][43] = 9'b111111111;
assign micromatr[21][44] = 9'b110010110;
assign micromatr[21][45] = 9'b110010110;
assign micromatr[21][46] = 9'b110111111;
assign micromatr[21][47] = 9'b111111111;
assign micromatr[21][48] = 9'b111111111;
assign micromatr[21][49] = 9'b111111111;
assign micromatr[21][50] = 9'b110011111;
assign micromatr[21][51] = 9'b110010010;
assign micromatr[21][52] = 9'b110010010;
assign micromatr[21][53] = 9'b111110010;
assign micromatr[21][54] = 9'b111111111;
assign micromatr[21][55] = 9'b111110111;
assign micromatr[21][56] = 9'b111110111;
assign micromatr[21][57] = 9'b111110111;
assign micromatr[21][58] = 9'b110010001;
assign micromatr[21][59] = 9'b111111111;
assign micromatr[21][60] = 9'b111111111;
assign micromatr[21][61] = 9'b111111111;
assign micromatr[21][62] = 9'b111111111;
assign micromatr[21][63] = 9'b111111111;
assign micromatr[21][64] = 9'b111111111;
assign micromatr[21][65] = 9'b110001101;
assign micromatr[21][66] = 9'b110110011;
assign micromatr[21][67] = 9'b111110111;
assign micromatr[21][68] = 9'b111110111;
assign micromatr[21][69] = 9'b111110111;
assign micromatr[21][70] = 9'b111110011;
assign micromatr[21][71] = 9'b110001101;
assign micromatr[21][72] = 9'b111110111;
assign micromatr[21][73] = 9'b110010110;
assign micromatr[21][74] = 9'b111111111;
assign micromatr[21][75] = 9'b111111111;
assign micromatr[21][76] = 9'b111111111;
assign micromatr[21][77] = 9'b111111111;
assign micromatr[21][78] = 9'b111111111;
assign micromatr[21][79] = 9'b111111111;
assign micromatr[21][80] = 9'b111111111;
assign micromatr[21][81] = 9'b111111111;
assign micromatr[21][82] = 9'b111111111;
assign micromatr[21][83] = 9'b110010110;
assign micromatr[21][84] = 9'b111111111;
assign micromatr[21][85] = 9'b111111111;
assign micromatr[21][86] = 9'b111111111;
assign micromatr[21][87] = 9'b111111111;
assign micromatr[21][88] = 9'b111111111;
assign micromatr[21][89] = 9'b111111111;
assign micromatr[21][90] = 9'b111111111;
assign micromatr[21][91] = 9'b111111111;
assign micromatr[21][92] = 9'b111111111;
assign micromatr[21][93] = 9'b111111111;
assign micromatr[21][94] = 9'b111111111;
assign micromatr[21][95] = 9'b111111111;
assign micromatr[21][96] = 9'b111111111;
assign micromatr[21][97] = 9'b111111111;
assign micromatr[21][98] = 9'b111111111;
assign micromatr[21][99] = 9'b111111111;
assign micromatr[22][0] = 9'b111111111;
assign micromatr[22][1] = 9'b111111111;
assign micromatr[22][2] = 9'b111111111;
assign micromatr[22][3] = 9'b111111111;
assign micromatr[22][4] = 9'b111111111;
assign micromatr[22][5] = 9'b111111111;
assign micromatr[22][6] = 9'b111111111;
assign micromatr[22][7] = 9'b111111111;
assign micromatr[22][8] = 9'b111111111;
assign micromatr[22][9] = 9'b111111111;
assign micromatr[22][10] = 9'b111111111;
assign micromatr[22][11] = 9'b111111111;
assign micromatr[22][12] = 9'b111111111;
assign micromatr[22][13] = 9'b111111111;
assign micromatr[22][14] = 9'b111111111;
assign micromatr[22][15] = 9'b110010010;
assign micromatr[22][16] = 9'b111110111;
assign micromatr[22][17] = 9'b111110111;
assign micromatr[22][18] = 9'b111110111;
assign micromatr[22][19] = 9'b111110111;
assign micromatr[22][20] = 9'b111110111;
assign micromatr[22][21] = 9'b101101101;
assign micromatr[22][22] = 9'b110110010;
assign micromatr[22][23] = 9'b111111111;
assign micromatr[22][24] = 9'b111110111;
assign micromatr[22][25] = 9'b111110111;
assign micromatr[22][26] = 9'b111110011;
assign micromatr[22][27] = 9'b110110010;
assign micromatr[22][28] = 9'b111111111;
assign micromatr[22][29] = 9'b111111111;
assign micromatr[22][30] = 9'b110110110;
assign micromatr[22][31] = 9'b110110011;
assign micromatr[22][32] = 9'b111110111;
assign micromatr[22][33] = 9'b111110111;
assign micromatr[22][34] = 9'b111110111;
assign micromatr[22][35] = 9'b111110011;
assign micromatr[22][36] = 9'b111110111;
assign micromatr[22][37] = 9'b111110111;
assign micromatr[22][38] = 9'b111110111;
assign micromatr[22][39] = 9'b111110111;
assign micromatr[22][40] = 9'b110110011;
assign micromatr[22][41] = 9'b110001101;
assign micromatr[22][42] = 9'b111111111;
assign micromatr[22][43] = 9'b111111111;
assign micromatr[22][44] = 9'b110010110;
assign micromatr[22][45] = 9'b111111111;
assign micromatr[22][46] = 9'b111111111;
assign micromatr[22][47] = 9'b111111111;
assign micromatr[22][48] = 9'b111111111;
assign micromatr[22][49] = 9'b111111111;
assign micromatr[22][50] = 9'b110011111;
assign micromatr[22][51] = 9'b110010110;
assign micromatr[22][52] = 9'b110010001;
assign micromatr[22][53] = 9'b111110010;
assign micromatr[22][54] = 9'b111111111;
assign micromatr[22][55] = 9'b111110111;
assign micromatr[22][56] = 9'b111110111;
assign micromatr[22][57] = 9'b111110111;
assign micromatr[22][58] = 9'b110010001;
assign micromatr[22][59] = 9'b111111111;
assign micromatr[22][60] = 9'b111111111;
assign micromatr[22][61] = 9'b111111111;
assign micromatr[22][62] = 9'b111111111;
assign micromatr[22][63] = 9'b111111111;
assign micromatr[22][64] = 9'b111111111;
assign micromatr[22][65] = 9'b110110010;
assign micromatr[22][66] = 9'b111111111;
assign micromatr[22][67] = 9'b111110111;
assign micromatr[22][68] = 9'b111110111;
assign micromatr[22][69] = 9'b111110111;
assign micromatr[22][70] = 9'b111110011;
assign micromatr[22][71] = 9'b110001101;
assign micromatr[22][72] = 9'b111110111;
assign micromatr[22][73] = 9'b110010010;
assign micromatr[22][74] = 9'b111111111;
assign micromatr[22][75] = 9'b111111111;
assign micromatr[22][76] = 9'b111111111;
assign micromatr[22][77] = 9'b110111111;
assign micromatr[22][78] = 9'b110010001;
assign micromatr[22][79] = 9'b110010001;
assign micromatr[22][80] = 9'b110010010;
assign micromatr[22][81] = 9'b110010110;
assign micromatr[22][82] = 9'b110010010;
assign micromatr[22][83] = 9'b111111111;
assign micromatr[22][84] = 9'b111111111;
assign micromatr[22][85] = 9'b111111111;
assign micromatr[22][86] = 9'b111111111;
assign micromatr[22][87] = 9'b111111111;
assign micromatr[22][88] = 9'b111111111;
assign micromatr[22][89] = 9'b111111111;
assign micromatr[22][90] = 9'b111111111;
assign micromatr[22][91] = 9'b111111111;
assign micromatr[22][92] = 9'b111111111;
assign micromatr[22][93] = 9'b111111111;
assign micromatr[22][94] = 9'b111111111;
assign micromatr[22][95] = 9'b111111111;
assign micromatr[22][96] = 9'b111111111;
assign micromatr[22][97] = 9'b111111111;
assign micromatr[22][98] = 9'b111111111;
assign micromatr[22][99] = 9'b111111111;
assign micromatr[23][0] = 9'b111111111;
assign micromatr[23][1] = 9'b111111111;
assign micromatr[23][2] = 9'b111111111;
assign micromatr[23][3] = 9'b111111111;
assign micromatr[23][4] = 9'b111111111;
assign micromatr[23][5] = 9'b111111111;
assign micromatr[23][6] = 9'b111111111;
assign micromatr[23][7] = 9'b111111111;
assign micromatr[23][8] = 9'b111111111;
assign micromatr[23][9] = 9'b111111111;
assign micromatr[23][10] = 9'b111111111;
assign micromatr[23][11] = 9'b111111111;
assign micromatr[23][12] = 9'b111111111;
assign micromatr[23][13] = 9'b111111111;
assign micromatr[23][14] = 9'b111111111;
assign micromatr[23][15] = 9'b110010001;
assign micromatr[23][16] = 9'b111110111;
assign micromatr[23][17] = 9'b111110111;
assign micromatr[23][18] = 9'b111110111;
assign micromatr[23][19] = 9'b111110111;
assign micromatr[23][20] = 9'b111110111;
assign micromatr[23][21] = 9'b110110001;
assign micromatr[23][22] = 9'b111110010;
assign micromatr[23][23] = 9'b111111111;
assign micromatr[23][24] = 9'b111110111;
assign micromatr[23][25] = 9'b111110111;
assign micromatr[23][26] = 9'b111110011;
assign micromatr[23][27] = 9'b110110010;
assign micromatr[23][28] = 9'b111111111;
assign micromatr[23][29] = 9'b111111111;
assign micromatr[23][30] = 9'b110010001;
assign micromatr[23][31] = 9'b111110111;
assign micromatr[23][32] = 9'b111110111;
assign micromatr[23][33] = 9'b111110111;
assign micromatr[23][34] = 9'b111111111;
assign micromatr[23][35] = 9'b101101101;
assign micromatr[23][36] = 9'b110010010;
assign micromatr[23][37] = 9'b111110111;
assign micromatr[23][38] = 9'b111110111;
assign micromatr[23][39] = 9'b111110111;
assign micromatr[23][40] = 9'b111110111;
assign micromatr[23][41] = 9'b110001101;
assign micromatr[23][42] = 9'b111111111;
assign micromatr[23][43] = 9'b111111111;
assign micromatr[23][44] = 9'b110010110;
assign micromatr[23][45] = 9'b111111111;
assign micromatr[23][46] = 9'b111111111;
assign micromatr[23][47] = 9'b111111111;
assign micromatr[23][48] = 9'b111111111;
assign micromatr[23][49] = 9'b111111111;
assign micromatr[23][50] = 9'b110011111;
assign micromatr[23][51] = 9'b111111111;
assign micromatr[23][52] = 9'b110010010;
assign micromatr[23][53] = 9'b111110010;
assign micromatr[23][54] = 9'b111111111;
assign micromatr[23][55] = 9'b111110111;
assign micromatr[23][56] = 9'b111110111;
assign micromatr[23][57] = 9'b111110111;
assign micromatr[23][58] = 9'b110110010;
assign micromatr[23][59] = 9'b111111111;
assign micromatr[23][60] = 9'b111111111;
assign micromatr[23][61] = 9'b111111111;
assign micromatr[23][62] = 9'b111111111;
assign micromatr[23][63] = 9'b111111111;
assign micromatr[23][64] = 9'b111111111;
assign micromatr[23][65] = 9'b110010010;
assign micromatr[23][66] = 9'b111110111;
assign micromatr[23][67] = 9'b111110111;
assign micromatr[23][68] = 9'b111110111;
assign micromatr[23][69] = 9'b111110111;
assign micromatr[23][70] = 9'b111110011;
assign micromatr[23][71] = 9'b110010010;
assign micromatr[23][72] = 9'b111111111;
assign micromatr[23][73] = 9'b110010010;
assign micromatr[23][74] = 9'b111111111;
assign micromatr[23][75] = 9'b111111111;
assign micromatr[23][76] = 9'b111111111;
assign micromatr[23][77] = 9'b110010111;
assign micromatr[23][78] = 9'b110010010;
assign micromatr[23][79] = 9'b110010110;
assign micromatr[23][80] = 9'b101110001;
assign micromatr[23][81] = 9'b111111111;
assign micromatr[23][82] = 9'b111111111;
assign micromatr[23][83] = 9'b111111111;
assign micromatr[23][84] = 9'b111111111;
assign micromatr[23][85] = 9'b111111111;
assign micromatr[23][86] = 9'b111111111;
assign micromatr[23][87] = 9'b111111111;
assign micromatr[23][88] = 9'b111111111;
assign micromatr[23][89] = 9'b111111111;
assign micromatr[23][90] = 9'b111111111;
assign micromatr[23][91] = 9'b111111111;
assign micromatr[23][92] = 9'b111111111;
assign micromatr[23][93] = 9'b111111111;
assign micromatr[23][94] = 9'b111111111;
assign micromatr[23][95] = 9'b111111111;
assign micromatr[23][96] = 9'b111111111;
assign micromatr[23][97] = 9'b111111111;
assign micromatr[23][98] = 9'b111111111;
assign micromatr[23][99] = 9'b111111111;
assign micromatr[24][0] = 9'b111111111;
assign micromatr[24][1] = 9'b111111111;
assign micromatr[24][2] = 9'b111111111;
assign micromatr[24][3] = 9'b111111111;
assign micromatr[24][4] = 9'b111111111;
assign micromatr[24][5] = 9'b111111111;
assign micromatr[24][6] = 9'b111111111;
assign micromatr[24][7] = 9'b111111111;
assign micromatr[24][8] = 9'b111111111;
assign micromatr[24][9] = 9'b111111111;
assign micromatr[24][10] = 9'b111111111;
assign micromatr[24][11] = 9'b111111111;
assign micromatr[24][12] = 9'b111111111;
assign micromatr[24][13] = 9'b111111111;
assign micromatr[24][14] = 9'b111111111;
assign micromatr[24][15] = 9'b110110010;
assign micromatr[24][16] = 9'b111110111;
assign micromatr[24][17] = 9'b111110111;
assign micromatr[24][18] = 9'b111110111;
assign micromatr[24][19] = 9'b111110111;
assign micromatr[24][20] = 9'b111110111;
assign micromatr[24][21] = 9'b111111111;
assign micromatr[24][22] = 9'b111110111;
assign micromatr[24][23] = 9'b111110111;
assign micromatr[24][24] = 9'b111110111;
assign micromatr[24][25] = 9'b111110111;
assign micromatr[24][26] = 9'b111110011;
assign micromatr[24][27] = 9'b110110010;
assign micromatr[24][28] = 9'b111111111;
assign micromatr[24][29] = 9'b111111111;
assign micromatr[24][30] = 9'b110010010;
assign micromatr[24][31] = 9'b111110111;
assign micromatr[24][32] = 9'b111110111;
assign micromatr[24][33] = 9'b111110111;
assign micromatr[24][34] = 9'b111110111;
assign micromatr[24][35] = 9'b110001101;
assign micromatr[24][36] = 9'b110001110;
assign micromatr[24][37] = 9'b111110111;
assign micromatr[24][38] = 9'b111110111;
assign micromatr[24][39] = 9'b111110111;
assign micromatr[24][40] = 9'b111110111;
assign micromatr[24][41] = 9'b110110010;
assign micromatr[24][42] = 9'b110010001;
assign micromatr[24][43] = 9'b111111111;
assign micromatr[24][44] = 9'b110110110;
assign micromatr[24][45] = 9'b111111111;
assign micromatr[24][46] = 9'b111111111;
assign micromatr[24][47] = 9'b111111111;
assign micromatr[24][48] = 9'b111111111;
assign micromatr[24][49] = 9'b111111111;
assign micromatr[24][50] = 9'b110011111;
assign micromatr[24][51] = 9'b111111111;
assign micromatr[24][52] = 9'b110010010;
assign micromatr[24][53] = 9'b111110010;
assign micromatr[24][54] = 9'b111111111;
assign micromatr[24][55] = 9'b111110111;
assign micromatr[24][56] = 9'b111110111;
assign micromatr[24][57] = 9'b111110111;
assign micromatr[24][58] = 9'b110001101;
assign micromatr[24][59] = 9'b110110010;
assign micromatr[24][60] = 9'b110010010;
assign micromatr[24][61] = 9'b110110110;
assign micromatr[24][62] = 9'b110110010;
assign micromatr[24][63] = 9'b110110110;
assign micromatr[24][64] = 9'b111111111;
assign micromatr[24][65] = 9'b110010010;
assign micromatr[24][66] = 9'b111110111;
assign micromatr[24][67] = 9'b111110111;
assign micromatr[24][68] = 9'b111110111;
assign micromatr[24][69] = 9'b111110111;
assign micromatr[24][70] = 9'b111110011;
assign micromatr[24][71] = 9'b110010010;
assign micromatr[24][72] = 9'b111111111;
assign micromatr[24][73] = 9'b110010010;
assign micromatr[24][74] = 9'b111111111;
assign micromatr[24][75] = 9'b111111111;
assign micromatr[24][76] = 9'b111111111;
assign micromatr[24][77] = 9'b111111111;
assign micromatr[24][78] = 9'b111111111;
assign micromatr[24][79] = 9'b111111111;
assign micromatr[24][80] = 9'b110010110;
assign micromatr[24][81] = 9'b110010001;
assign micromatr[24][82] = 9'b111111111;
assign micromatr[24][83] = 9'b111111111;
assign micromatr[24][84] = 9'b111111111;
assign micromatr[24][85] = 9'b111111111;
assign micromatr[24][86] = 9'b111111111;
assign micromatr[24][87] = 9'b111111111;
assign micromatr[24][88] = 9'b111111111;
assign micromatr[24][89] = 9'b111111111;
assign micromatr[24][90] = 9'b111111111;
assign micromatr[24][91] = 9'b111111111;
assign micromatr[24][92] = 9'b111111111;
assign micromatr[24][93] = 9'b111111111;
assign micromatr[24][94] = 9'b111111111;
assign micromatr[24][95] = 9'b111111111;
assign micromatr[24][96] = 9'b111111111;
assign micromatr[24][97] = 9'b111111111;
assign micromatr[24][98] = 9'b111111111;
assign micromatr[24][99] = 9'b111111111;
assign micromatr[25][0] = 9'b111111111;
assign micromatr[25][1] = 9'b111111111;
assign micromatr[25][2] = 9'b111111111;
assign micromatr[25][3] = 9'b111111111;
assign micromatr[25][4] = 9'b111111111;
assign micromatr[25][5] = 9'b111111111;
assign micromatr[25][6] = 9'b111111111;
assign micromatr[25][7] = 9'b111111111;
assign micromatr[25][8] = 9'b111111111;
assign micromatr[25][9] = 9'b111111111;
assign micromatr[25][10] = 9'b111111111;
assign micromatr[25][11] = 9'b111111111;
assign micromatr[25][12] = 9'b111111111;
assign micromatr[25][13] = 9'b111111111;
assign micromatr[25][14] = 9'b111111111;
assign micromatr[25][15] = 9'b110110010;
assign micromatr[25][16] = 9'b111110111;
assign micromatr[25][17] = 9'b111110111;
assign micromatr[25][18] = 9'b111110111;
assign micromatr[25][19] = 9'b111110111;
assign micromatr[25][20] = 9'b111110111;
assign micromatr[25][21] = 9'b111110111;
assign micromatr[25][22] = 9'b111110111;
assign micromatr[25][23] = 9'b111110111;
assign micromatr[25][24] = 9'b111110111;
assign micromatr[25][25] = 9'b111110111;
assign micromatr[25][26] = 9'b111110011;
assign micromatr[25][27] = 9'b110110010;
assign micromatr[25][28] = 9'b111111111;
assign micromatr[25][29] = 9'b110010010;
assign micromatr[25][30] = 9'b111110011;
assign micromatr[25][31] = 9'b111110111;
assign micromatr[25][32] = 9'b111110111;
assign micromatr[25][33] = 9'b111110111;
assign micromatr[25][34] = 9'b111110011;
assign micromatr[25][35] = 9'b101101101;
assign micromatr[25][36] = 9'b110001101;
assign micromatr[25][37] = 9'b111110111;
assign micromatr[25][38] = 9'b111110111;
assign micromatr[25][39] = 9'b111110111;
assign micromatr[25][40] = 9'b111110111;
assign micromatr[25][41] = 9'b111110111;
assign micromatr[25][42] = 9'b101101101;
assign micromatr[25][43] = 9'b111111111;
assign micromatr[25][44] = 9'b110110110;
assign micromatr[25][45] = 9'b111111111;
assign micromatr[25][46] = 9'b111111111;
assign micromatr[25][47] = 9'b111111111;
assign micromatr[25][48] = 9'b111111111;
assign micromatr[25][49] = 9'b111111111;
assign micromatr[25][50] = 9'b110011111;
assign micromatr[25][51] = 9'b111111111;
assign micromatr[25][52] = 9'b110010010;
assign micromatr[25][53] = 9'b111110010;
assign micromatr[25][54] = 9'b111111111;
assign micromatr[25][55] = 9'b111110111;
assign micromatr[25][56] = 9'b111110111;
assign micromatr[25][57] = 9'b111110111;
assign micromatr[25][58] = 9'b111110011;
assign micromatr[25][59] = 9'b111110010;
assign micromatr[25][60] = 9'b111110010;
assign micromatr[25][61] = 9'b111110011;
assign micromatr[25][62] = 9'b111110011;
assign micromatr[25][63] = 9'b110110010;
assign micromatr[25][64] = 9'b110110110;
assign micromatr[25][65] = 9'b110010010;
assign micromatr[25][66] = 9'b111110111;
assign micromatr[25][67] = 9'b111110111;
assign micromatr[25][68] = 9'b111110111;
assign micromatr[25][69] = 9'b111110111;
assign micromatr[25][70] = 9'b111110011;
assign micromatr[25][71] = 9'b110010010;
assign micromatr[25][72] = 9'b111111111;
assign micromatr[25][73] = 9'b110010010;
assign micromatr[25][74] = 9'b111111111;
assign micromatr[25][75] = 9'b111111111;
assign micromatr[25][76] = 9'b111111111;
assign micromatr[25][77] = 9'b111111111;
assign micromatr[25][78] = 9'b111111111;
assign micromatr[25][79] = 9'b111111111;
assign micromatr[25][80] = 9'b110010010;
assign micromatr[25][81] = 9'b111111111;
assign micromatr[25][82] = 9'b111111111;
assign micromatr[25][83] = 9'b111111111;
assign micromatr[25][84] = 9'b111111111;
assign micromatr[25][85] = 9'b111111111;
assign micromatr[25][86] = 9'b111111111;
assign micromatr[25][87] = 9'b111111111;
assign micromatr[25][88] = 9'b111111111;
assign micromatr[25][89] = 9'b111111111;
assign micromatr[25][90] = 9'b111111111;
assign micromatr[25][91] = 9'b111111111;
assign micromatr[25][92] = 9'b111111111;
assign micromatr[25][93] = 9'b111111111;
assign micromatr[25][94] = 9'b111111111;
assign micromatr[25][95] = 9'b111111111;
assign micromatr[25][96] = 9'b111111111;
assign micromatr[25][97] = 9'b111111111;
assign micromatr[25][98] = 9'b111111111;
assign micromatr[25][99] = 9'b111111111;
assign micromatr[26][0] = 9'b111111111;
assign micromatr[26][1] = 9'b111111111;
assign micromatr[26][2] = 9'b111111111;
assign micromatr[26][3] = 9'b111111111;
assign micromatr[26][4] = 9'b111111111;
assign micromatr[26][5] = 9'b111111111;
assign micromatr[26][6] = 9'b111111111;
assign micromatr[26][7] = 9'b111111111;
assign micromatr[26][8] = 9'b111111111;
assign micromatr[26][9] = 9'b111111111;
assign micromatr[26][10] = 9'b111111111;
assign micromatr[26][11] = 9'b111111111;
assign micromatr[26][12] = 9'b111111111;
assign micromatr[26][13] = 9'b111111111;
assign micromatr[26][14] = 9'b111111111;
assign micromatr[26][15] = 9'b110110010;
assign micromatr[26][16] = 9'b111110111;
assign micromatr[26][17] = 9'b111110111;
assign micromatr[26][18] = 9'b111110111;
assign micromatr[26][19] = 9'b111110111;
assign micromatr[26][20] = 9'b111110111;
assign micromatr[26][21] = 9'b111110111;
assign micromatr[26][22] = 9'b111110111;
assign micromatr[26][23] = 9'b111110111;
assign micromatr[26][24] = 9'b111110111;
assign micromatr[26][25] = 9'b111110111;
assign micromatr[26][26] = 9'b111110011;
assign micromatr[26][27] = 9'b110110010;
assign micromatr[26][28] = 9'b111111111;
assign micromatr[26][29] = 9'b110001101;
assign micromatr[26][30] = 9'b111110111;
assign micromatr[26][31] = 9'b111110111;
assign micromatr[26][32] = 9'b111110111;
assign micromatr[26][33] = 9'b111110111;
assign micromatr[26][34] = 9'b111110111;
assign micromatr[26][35] = 9'b110110011;
assign micromatr[26][36] = 9'b111110011;
assign micromatr[26][37] = 9'b111110111;
assign micromatr[26][38] = 9'b111110111;
assign micromatr[26][39] = 9'b111110111;
assign micromatr[26][40] = 9'b111110111;
assign micromatr[26][41] = 9'b111110111;
assign micromatr[26][42] = 9'b110010010;
assign micromatr[26][43] = 9'b110010010;
assign micromatr[26][44] = 9'b110010110;
assign micromatr[26][45] = 9'b111111111;
assign micromatr[26][46] = 9'b111111111;
assign micromatr[26][47] = 9'b111111111;
assign micromatr[26][48] = 9'b111111111;
assign micromatr[26][49] = 9'b111111111;
assign micromatr[26][50] = 9'b110011111;
assign micromatr[26][51] = 9'b111111111;
assign micromatr[26][52] = 9'b110010110;
assign micromatr[26][53] = 9'b111110010;
assign micromatr[26][54] = 9'b111111111;
assign micromatr[26][55] = 9'b111110111;
assign micromatr[26][56] = 9'b111110111;
assign micromatr[26][57] = 9'b111110111;
assign micromatr[26][58] = 9'b111110111;
assign micromatr[26][59] = 9'b111111111;
assign micromatr[26][60] = 9'b111110111;
assign micromatr[26][61] = 9'b111110111;
assign micromatr[26][62] = 9'b111111111;
assign micromatr[26][63] = 9'b110110010;
assign micromatr[26][64] = 9'b110010001;
assign micromatr[26][65] = 9'b110010010;
assign micromatr[26][66] = 9'b111110111;
assign micromatr[26][67] = 9'b111110111;
assign micromatr[26][68] = 9'b111110111;
assign micromatr[26][69] = 9'b111110111;
assign micromatr[26][70] = 9'b111110011;
assign micromatr[26][71] = 9'b110010010;
assign micromatr[26][72] = 9'b111111111;
assign micromatr[26][73] = 9'b110010001;
assign micromatr[26][74] = 9'b111111111;
assign micromatr[26][75] = 9'b111111111;
assign micromatr[26][76] = 9'b111111111;
assign micromatr[26][77] = 9'b111111111;
assign micromatr[26][78] = 9'b101101101;
assign micromatr[26][79] = 9'b101101101;
assign micromatr[26][80] = 9'b101101101;
assign micromatr[26][81] = 9'b110010110;
assign micromatr[26][82] = 9'b110010010;
assign micromatr[26][83] = 9'b111111111;
assign micromatr[26][84] = 9'b111111111;
assign micromatr[26][85] = 9'b111111111;
assign micromatr[26][86] = 9'b111111111;
assign micromatr[26][87] = 9'b111111111;
assign micromatr[26][88] = 9'b111111111;
assign micromatr[26][89] = 9'b111111111;
assign micromatr[26][90] = 9'b111111111;
assign micromatr[26][91] = 9'b111111111;
assign micromatr[26][92] = 9'b111111111;
assign micromatr[26][93] = 9'b111111111;
assign micromatr[26][94] = 9'b111111111;
assign micromatr[26][95] = 9'b111111111;
assign micromatr[26][96] = 9'b111111111;
assign micromatr[26][97] = 9'b111111111;
assign micromatr[26][98] = 9'b111111111;
assign micromatr[26][99] = 9'b111111111;
assign micromatr[27][0] = 9'b111111111;
assign micromatr[27][1] = 9'b111111111;
assign micromatr[27][2] = 9'b111111111;
assign micromatr[27][3] = 9'b111111111;
assign micromatr[27][4] = 9'b111111111;
assign micromatr[27][5] = 9'b111111111;
assign micromatr[27][6] = 9'b111111111;
assign micromatr[27][7] = 9'b111111111;
assign micromatr[27][8] = 9'b111111111;
assign micromatr[27][9] = 9'b111111111;
assign micromatr[27][10] = 9'b111111111;
assign micromatr[27][11] = 9'b111111111;
assign micromatr[27][12] = 9'b111111111;
assign micromatr[27][13] = 9'b111111111;
assign micromatr[27][14] = 9'b111111111;
assign micromatr[27][15] = 9'b110010010;
assign micromatr[27][16] = 9'b111110111;
assign micromatr[27][17] = 9'b111110111;
assign micromatr[27][18] = 9'b111110111;
assign micromatr[27][19] = 9'b111110111;
assign micromatr[27][20] = 9'b110001101;
assign micromatr[27][21] = 9'b110110010;
assign micromatr[27][22] = 9'b111110111;
assign micromatr[27][23] = 9'b111110111;
assign micromatr[27][24] = 9'b111110111;
assign micromatr[27][25] = 9'b111110111;
assign micromatr[27][26] = 9'b111110011;
assign micromatr[27][27] = 9'b111110010;
assign micromatr[27][28] = 9'b110010010;
assign micromatr[27][29] = 9'b110010010;
assign micromatr[27][30] = 9'b111110111;
assign micromatr[27][31] = 9'b111110111;
assign micromatr[27][32] = 9'b111110111;
assign micromatr[27][33] = 9'b111110111;
assign micromatr[27][34] = 9'b111110111;
assign micromatr[27][35] = 9'b111110111;
assign micromatr[27][36] = 9'b111110111;
assign micromatr[27][37] = 9'b111110111;
assign micromatr[27][38] = 9'b111110111;
assign micromatr[27][39] = 9'b111110111;
assign micromatr[27][40] = 9'b111110111;
assign micromatr[27][41] = 9'b111110111;
assign micromatr[27][42] = 9'b111110111;
assign micromatr[27][43] = 9'b110001101;
assign micromatr[27][44] = 9'b110010001;
assign micromatr[27][45] = 9'b111111111;
assign micromatr[27][46] = 9'b111111111;
assign micromatr[27][47] = 9'b111111111;
assign micromatr[27][48] = 9'b111111111;
assign micromatr[27][49] = 9'b111111111;
assign micromatr[27][50] = 9'b110011111;
assign micromatr[27][51] = 9'b111111111;
assign micromatr[27][52] = 9'b110010110;
assign micromatr[27][53] = 9'b111110010;
assign micromatr[27][54] = 9'b111111111;
assign micromatr[27][55] = 9'b111110111;
assign micromatr[27][56] = 9'b111110111;
assign micromatr[27][57] = 9'b111110111;
assign micromatr[27][58] = 9'b111110111;
assign micromatr[27][59] = 9'b111110111;
assign micromatr[27][60] = 9'b111110111;
assign micromatr[27][61] = 9'b111110111;
assign micromatr[27][62] = 9'b111110111;
assign micromatr[27][63] = 9'b110110010;
assign micromatr[27][64] = 9'b111110110;
assign micromatr[27][65] = 9'b110010010;
assign micromatr[27][66] = 9'b111110111;
assign micromatr[27][67] = 9'b111110111;
assign micromatr[27][68] = 9'b111110111;
assign micromatr[27][69] = 9'b111110111;
assign micromatr[27][70] = 9'b111110011;
assign micromatr[27][71] = 9'b110010010;
assign micromatr[27][72] = 9'b111111111;
assign micromatr[27][73] = 9'b110010001;
assign micromatr[27][74] = 9'b111111111;
assign micromatr[27][75] = 9'b111111111;
assign micromatr[27][76] = 9'b111111111;
assign micromatr[27][77] = 9'b111111111;
assign micromatr[27][78] = 9'b111111111;
assign micromatr[27][79] = 9'b111111111;
assign micromatr[27][80] = 9'b111111111;
assign micromatr[27][81] = 9'b110111111;
assign micromatr[27][82] = 9'b110010010;
assign micromatr[27][83] = 9'b111111111;
assign micromatr[27][84] = 9'b111111111;
assign micromatr[27][85] = 9'b111111111;
assign micromatr[27][86] = 9'b111111111;
assign micromatr[27][87] = 9'b111111111;
assign micromatr[27][88] = 9'b111111111;
assign micromatr[27][89] = 9'b111111111;
assign micromatr[27][90] = 9'b111111111;
assign micromatr[27][91] = 9'b111111111;
assign micromatr[27][92] = 9'b111111111;
assign micromatr[27][93] = 9'b111111111;
assign micromatr[27][94] = 9'b111111111;
assign micromatr[27][95] = 9'b111111111;
assign micromatr[27][96] = 9'b111111111;
assign micromatr[27][97] = 9'b111111111;
assign micromatr[27][98] = 9'b111111111;
assign micromatr[27][99] = 9'b111111111;
assign micromatr[28][0] = 9'b111111111;
assign micromatr[28][1] = 9'b111111111;
assign micromatr[28][2] = 9'b111111111;
assign micromatr[28][3] = 9'b111111111;
assign micromatr[28][4] = 9'b111111111;
assign micromatr[28][5] = 9'b111111111;
assign micromatr[28][6] = 9'b111111111;
assign micromatr[28][7] = 9'b111111111;
assign micromatr[28][8] = 9'b111111111;
assign micromatr[28][9] = 9'b111111111;
assign micromatr[28][10] = 9'b111111111;
assign micromatr[28][11] = 9'b111111111;
assign micromatr[28][12] = 9'b111111111;
assign micromatr[28][13] = 9'b111111111;
assign micromatr[28][14] = 9'b111111111;
assign micromatr[28][15] = 9'b110110010;
assign micromatr[28][16] = 9'b111110111;
assign micromatr[28][17] = 9'b111110111;
assign micromatr[28][18] = 9'b111110111;
assign micromatr[28][19] = 9'b111110011;
assign micromatr[28][20] = 9'b110010001;
assign micromatr[28][21] = 9'b110110010;
assign micromatr[28][22] = 9'b111110111;
assign micromatr[28][23] = 9'b111110111;
assign micromatr[28][24] = 9'b111110111;
assign micromatr[28][25] = 9'b111110111;
assign micromatr[28][26] = 9'b111110011;
assign micromatr[28][27] = 9'b110110010;
assign micromatr[28][28] = 9'b110010010;
assign micromatr[28][29] = 9'b111110011;
assign micromatr[28][30] = 9'b111110111;
assign micromatr[28][31] = 9'b111110111;
assign micromatr[28][32] = 9'b111110111;
assign micromatr[28][33] = 9'b111110111;
assign micromatr[28][34] = 9'b111110111;
assign micromatr[28][35] = 9'b111110111;
assign micromatr[28][36] = 9'b111110111;
assign micromatr[28][37] = 9'b111110111;
assign micromatr[28][38] = 9'b111110111;
assign micromatr[28][39] = 9'b111110111;
assign micromatr[28][40] = 9'b111110111;
assign micromatr[28][41] = 9'b111110111;
assign micromatr[28][42] = 9'b111110111;
assign micromatr[28][43] = 9'b110010010;
assign micromatr[28][44] = 9'b101101101;
assign micromatr[28][45] = 9'b111111111;
assign micromatr[28][46] = 9'b111111111;
assign micromatr[28][47] = 9'b111111111;
assign micromatr[28][48] = 9'b111111111;
assign micromatr[28][49] = 9'b111111111;
assign micromatr[28][50] = 9'b110011111;
assign micromatr[28][51] = 9'b111111111;
assign micromatr[28][52] = 9'b110110110;
assign micromatr[28][53] = 9'b111110010;
assign micromatr[28][54] = 9'b111111111;
assign micromatr[28][55] = 9'b111110111;
assign micromatr[28][56] = 9'b111110111;
assign micromatr[28][57] = 9'b111110111;
assign micromatr[28][58] = 9'b111110111;
assign micromatr[28][59] = 9'b111110111;
assign micromatr[28][60] = 9'b111110111;
assign micromatr[28][61] = 9'b111110111;
assign micromatr[28][62] = 9'b111110111;
assign micromatr[28][63] = 9'b110110010;
assign micromatr[28][64] = 9'b111110010;
assign micromatr[28][65] = 9'b110010010;
assign micromatr[28][66] = 9'b111110111;
assign micromatr[28][67] = 9'b111110111;
assign micromatr[28][68] = 9'b111110111;
assign micromatr[28][69] = 9'b111110111;
assign micromatr[28][70] = 9'b111110011;
assign micromatr[28][71] = 9'b110010010;
assign micromatr[28][72] = 9'b111111111;
assign micromatr[28][73] = 9'b110010010;
assign micromatr[28][74] = 9'b111111111;
assign micromatr[28][75] = 9'b111111111;
assign micromatr[28][76] = 9'b111111111;
assign micromatr[28][77] = 9'b111111111;
assign micromatr[28][78] = 9'b111111111;
assign micromatr[28][79] = 9'b111111111;
assign micromatr[28][80] = 9'b111111111;
assign micromatr[28][81] = 9'b111111111;
assign micromatr[28][82] = 9'b110111111;
assign micromatr[28][83] = 9'b110010001;
assign micromatr[28][84] = 9'b111111111;
assign micromatr[28][85] = 9'b111111111;
assign micromatr[28][86] = 9'b111111111;
assign micromatr[28][87] = 9'b111111111;
assign micromatr[28][88] = 9'b111111111;
assign micromatr[28][89] = 9'b111111111;
assign micromatr[28][90] = 9'b111111111;
assign micromatr[28][91] = 9'b111111111;
assign micromatr[28][92] = 9'b111111111;
assign micromatr[28][93] = 9'b111111111;
assign micromatr[28][94] = 9'b111111111;
assign micromatr[28][95] = 9'b111111111;
assign micromatr[28][96] = 9'b111111111;
assign micromatr[28][97] = 9'b111111111;
assign micromatr[28][98] = 9'b111111111;
assign micromatr[28][99] = 9'b111111111;
assign micromatr[29][0] = 9'b111111111;
assign micromatr[29][1] = 9'b111111111;
assign micromatr[29][2] = 9'b111111111;
assign micromatr[29][3] = 9'b111111111;
assign micromatr[29][4] = 9'b111111111;
assign micromatr[29][5] = 9'b111111111;
assign micromatr[29][6] = 9'b111111111;
assign micromatr[29][7] = 9'b111111111;
assign micromatr[29][8] = 9'b111111111;
assign micromatr[29][9] = 9'b111111111;
assign micromatr[29][10] = 9'b111111111;
assign micromatr[29][11] = 9'b111111111;
assign micromatr[29][12] = 9'b111111111;
assign micromatr[29][13] = 9'b111111111;
assign micromatr[29][14] = 9'b111111111;
assign micromatr[29][15] = 9'b110110010;
assign micromatr[29][16] = 9'b111111111;
assign micromatr[29][17] = 9'b111110111;
assign micromatr[29][18] = 9'b111110111;
assign micromatr[29][19] = 9'b111110011;
assign micromatr[29][20] = 9'b110010010;
assign micromatr[29][21] = 9'b110110010;
assign micromatr[29][22] = 9'b111110111;
assign micromatr[29][23] = 9'b111110111;
assign micromatr[29][24] = 9'b111110111;
assign micromatr[29][25] = 9'b111110111;
assign micromatr[29][26] = 9'b111110011;
assign micromatr[29][27] = 9'b110001101;
assign micromatr[29][28] = 9'b110010010;
assign micromatr[29][29] = 9'b111110111;
assign micromatr[29][30] = 9'b111110111;
assign micromatr[29][31] = 9'b111110111;
assign micromatr[29][32] = 9'b111110111;
assign micromatr[29][33] = 9'b111110111;
assign micromatr[29][34] = 9'b111110111;
assign micromatr[29][35] = 9'b111110011;
assign micromatr[29][36] = 9'b110001110;
assign micromatr[29][37] = 9'b110110011;
assign micromatr[29][38] = 9'b111110111;
assign micromatr[29][39] = 9'b111110111;
assign micromatr[29][40] = 9'b111110111;
assign micromatr[29][41] = 9'b111110111;
assign micromatr[29][42] = 9'b111110111;
assign micromatr[29][43] = 9'b111110111;
assign micromatr[29][44] = 9'b101001001;
assign micromatr[29][45] = 9'b111111111;
assign micromatr[29][46] = 9'b111111111;
assign micromatr[29][47] = 9'b111111111;
assign micromatr[29][48] = 9'b111111111;
assign micromatr[29][49] = 9'b111111111;
assign micromatr[29][50] = 9'b110011111;
assign micromatr[29][51] = 9'b111111111;
assign micromatr[29][52] = 9'b110110110;
assign micromatr[29][53] = 9'b111110010;
assign micromatr[29][54] = 9'b111111111;
assign micromatr[29][55] = 9'b111110111;
assign micromatr[29][56] = 9'b111110111;
assign micromatr[29][57] = 9'b111110111;
assign micromatr[29][58] = 9'b111110111;
assign micromatr[29][59] = 9'b111110111;
assign micromatr[29][60] = 9'b111110111;
assign micromatr[29][61] = 9'b111110111;
assign micromatr[29][62] = 9'b111110111;
assign micromatr[29][63] = 9'b110110010;
assign micromatr[29][64] = 9'b111110010;
assign micromatr[29][65] = 9'b110010010;
assign micromatr[29][66] = 9'b111110111;
assign micromatr[29][67] = 9'b111110111;
assign micromatr[29][68] = 9'b111110111;
assign micromatr[29][69] = 9'b111110111;
assign micromatr[29][70] = 9'b111110011;
assign micromatr[29][71] = 9'b110010010;
assign micromatr[29][72] = 9'b111111111;
assign micromatr[29][73] = 9'b110010010;
assign micromatr[29][74] = 9'b111111111;
assign micromatr[29][75] = 9'b111111111;
assign micromatr[29][76] = 9'b111111111;
assign micromatr[29][77] = 9'b111111111;
assign micromatr[29][78] = 9'b111111111;
assign micromatr[29][79] = 9'b111111111;
assign micromatr[29][80] = 9'b111111111;
assign micromatr[29][81] = 9'b111111111;
assign micromatr[29][82] = 9'b111111111;
assign micromatr[29][83] = 9'b110010110;
assign micromatr[29][84] = 9'b111111111;
assign micromatr[29][85] = 9'b111111111;
assign micromatr[29][86] = 9'b111111111;
assign micromatr[29][87] = 9'b111111111;
assign micromatr[29][88] = 9'b111111111;
assign micromatr[29][89] = 9'b111111111;
assign micromatr[29][90] = 9'b111111111;
assign micromatr[29][91] = 9'b111111111;
assign micromatr[29][92] = 9'b111111111;
assign micromatr[29][93] = 9'b111111111;
assign micromatr[29][94] = 9'b111111111;
assign micromatr[29][95] = 9'b111111111;
assign micromatr[29][96] = 9'b111111111;
assign micromatr[29][97] = 9'b111111111;
assign micromatr[29][98] = 9'b111111111;
assign micromatr[29][99] = 9'b111111111;
assign micromatr[30][0] = 9'b111111111;
assign micromatr[30][1] = 9'b111111111;
assign micromatr[30][2] = 9'b111111111;
assign micromatr[30][3] = 9'b111111111;
assign micromatr[30][4] = 9'b111111111;
assign micromatr[30][5] = 9'b111111111;
assign micromatr[30][6] = 9'b111111111;
assign micromatr[30][7] = 9'b111111111;
assign micromatr[30][8] = 9'b111111111;
assign micromatr[30][9] = 9'b111111111;
assign micromatr[30][10] = 9'b111111111;
assign micromatr[30][11] = 9'b111111111;
assign micromatr[30][12] = 9'b111111111;
assign micromatr[30][13] = 9'b111111111;
assign micromatr[30][14] = 9'b111111111;
assign micromatr[30][15] = 9'b110110010;
assign micromatr[30][16] = 9'b111111111;
assign micromatr[30][17] = 9'b111110111;
assign micromatr[30][18] = 9'b111110111;
assign micromatr[30][19] = 9'b111110011;
assign micromatr[30][20] = 9'b110010010;
assign micromatr[30][21] = 9'b110110010;
assign micromatr[30][22] = 9'b111111111;
assign micromatr[30][23] = 9'b111111111;
assign micromatr[30][24] = 9'b111111111;
assign micromatr[30][25] = 9'b111111111;
assign micromatr[30][26] = 9'b111110111;
assign micromatr[30][27] = 9'b101101101;
assign micromatr[30][28] = 9'b110010010;
assign micromatr[30][29] = 9'b111111111;
assign micromatr[30][30] = 9'b111110111;
assign micromatr[30][31] = 9'b111110111;
assign micromatr[30][32] = 9'b111110111;
assign micromatr[30][33] = 9'b111110111;
assign micromatr[30][34] = 9'b110110011;
assign micromatr[30][35] = 9'b110001101;
assign micromatr[30][36] = 9'b111110111;
assign micromatr[30][37] = 9'b110001101;
assign micromatr[30][38] = 9'b111110111;
assign micromatr[30][39] = 9'b111110111;
assign micromatr[30][40] = 9'b111110111;
assign micromatr[30][41] = 9'b111110111;
assign micromatr[30][42] = 9'b111110011;
assign micromatr[30][43] = 9'b110001110;
assign micromatr[30][44] = 9'b101101101;
assign micromatr[30][45] = 9'b111111111;
assign micromatr[30][46] = 9'b111111111;
assign micromatr[30][47] = 9'b111111111;
assign micromatr[30][48] = 9'b111111111;
assign micromatr[30][49] = 9'b111111111;
assign micromatr[30][50] = 9'b110011111;
assign micromatr[30][51] = 9'b111111111;
assign micromatr[30][52] = 9'b110110110;
assign micromatr[30][53] = 9'b110110010;
assign micromatr[30][54] = 9'b111111111;
assign micromatr[30][55] = 9'b111110111;
assign micromatr[30][56] = 9'b111110111;
assign micromatr[30][57] = 9'b111110111;
assign micromatr[30][58] = 9'b111110111;
assign micromatr[30][59] = 9'b111110111;
assign micromatr[30][60] = 9'b111110111;
assign micromatr[30][61] = 9'b111111111;
assign micromatr[30][62] = 9'b111111111;
assign micromatr[30][63] = 9'b110110010;
assign micromatr[30][64] = 9'b111110010;
assign micromatr[30][65] = 9'b110010010;
assign micromatr[30][66] = 9'b111110111;
assign micromatr[30][67] = 9'b111110111;
assign micromatr[30][68] = 9'b111110111;
assign micromatr[30][69] = 9'b111110111;
assign micromatr[30][70] = 9'b111110011;
assign micromatr[30][71] = 9'b110010010;
assign micromatr[30][72] = 9'b111111111;
assign micromatr[30][73] = 9'b110010010;
assign micromatr[30][74] = 9'b111111111;
assign micromatr[30][75] = 9'b111111111;
assign micromatr[30][76] = 9'b111111111;
assign micromatr[30][77] = 9'b111111111;
assign micromatr[30][78] = 9'b111111111;
assign micromatr[30][79] = 9'b111111111;
assign micromatr[30][80] = 9'b110111111;
assign micromatr[30][81] = 9'b110011111;
assign micromatr[30][82] = 9'b110010010;
assign micromatr[30][83] = 9'b110110110;
assign micromatr[30][84] = 9'b111111111;
assign micromatr[30][85] = 9'b111111111;
assign micromatr[30][86] = 9'b111111111;
assign micromatr[30][87] = 9'b111111111;
assign micromatr[30][88] = 9'b111111111;
assign micromatr[30][89] = 9'b111111111;
assign micromatr[30][90] = 9'b111111111;
assign micromatr[30][91] = 9'b111111111;
assign micromatr[30][92] = 9'b111111111;
assign micromatr[30][93] = 9'b111111111;
assign micromatr[30][94] = 9'b111111111;
assign micromatr[30][95] = 9'b111111111;
assign micromatr[30][96] = 9'b111111111;
assign micromatr[30][97] = 9'b111111111;
assign micromatr[30][98] = 9'b111111111;
assign micromatr[30][99] = 9'b111111111;
assign micromatr[31][0] = 9'b111111111;
assign micromatr[31][1] = 9'b111111111;
assign micromatr[31][2] = 9'b111111111;
assign micromatr[31][3] = 9'b111111111;
assign micromatr[31][4] = 9'b111111111;
assign micromatr[31][5] = 9'b111111111;
assign micromatr[31][6] = 9'b111111111;
assign micromatr[31][7] = 9'b111111111;
assign micromatr[31][8] = 9'b111111111;
assign micromatr[31][9] = 9'b111111111;
assign micromatr[31][10] = 9'b111111111;
assign micromatr[31][11] = 9'b111111111;
assign micromatr[31][12] = 9'b111111111;
assign micromatr[31][13] = 9'b111111111;
assign micromatr[31][14] = 9'b111111111;
assign micromatr[31][15] = 9'b110001101;
assign micromatr[31][16] = 9'b111110011;
assign micromatr[31][17] = 9'b111110111;
assign micromatr[31][18] = 9'b111111111;
assign micromatr[31][19] = 9'b111110011;
assign micromatr[31][20] = 9'b110110010;
assign micromatr[31][21] = 9'b110010001;
assign micromatr[31][22] = 9'b110110010;
assign micromatr[31][23] = 9'b110110010;
assign micromatr[31][24] = 9'b111110010;
assign micromatr[31][25] = 9'b111110010;
assign micromatr[31][26] = 9'b110101110;
assign micromatr[31][27] = 9'b110110010;
assign micromatr[31][28] = 9'b110010010;
assign micromatr[31][29] = 9'b101101101;
assign micromatr[31][30] = 9'b111110011;
assign micromatr[31][31] = 9'b111110111;
assign micromatr[31][32] = 9'b111110111;
assign micromatr[31][33] = 9'b111110111;
assign micromatr[31][34] = 9'b110001101;
assign micromatr[31][35] = 9'b111111111;
assign micromatr[31][36] = 9'b111111111;
assign micromatr[31][37] = 9'b110010001;
assign micromatr[31][38] = 9'b110010010;
assign micromatr[31][39] = 9'b111111111;
assign micromatr[31][40] = 9'b111110111;
assign micromatr[31][41] = 9'b110001110;
assign micromatr[31][42] = 9'b110001101;
assign micromatr[31][43] = 9'b111110111;
assign micromatr[31][44] = 9'b110010010;
assign micromatr[31][45] = 9'b111111111;
assign micromatr[31][46] = 9'b111111111;
assign micromatr[31][47] = 9'b111111111;
assign micromatr[31][48] = 9'b111111111;
assign micromatr[31][49] = 9'b111111111;
assign micromatr[31][50] = 9'b110010010;
assign micromatr[31][51] = 9'b110111111;
assign micromatr[31][52] = 9'b110110110;
assign micromatr[31][53] = 9'b110001101;
assign micromatr[31][54] = 9'b111110111;
assign micromatr[31][55] = 9'b111110111;
assign micromatr[31][56] = 9'b111110011;
assign micromatr[31][57] = 9'b111110011;
assign micromatr[31][58] = 9'b111110011;
assign micromatr[31][59] = 9'b111110011;
assign micromatr[31][60] = 9'b111110010;
assign micromatr[31][61] = 9'b111110010;
assign micromatr[31][62] = 9'b111110010;
assign micromatr[31][63] = 9'b110010001;
assign micromatr[31][64] = 9'b111110110;
assign micromatr[31][65] = 9'b110110010;
assign micromatr[31][66] = 9'b111111111;
assign micromatr[31][67] = 9'b111110111;
assign micromatr[31][68] = 9'b111110111;
assign micromatr[31][69] = 9'b111110011;
assign micromatr[31][70] = 9'b110110011;
assign micromatr[31][71] = 9'b110010010;
assign micromatr[31][72] = 9'b111111111;
assign micromatr[31][73] = 9'b110010001;
assign micromatr[31][74] = 9'b110111111;
assign micromatr[31][75] = 9'b110111111;
assign micromatr[31][76] = 9'b110011111;
assign micromatr[31][77] = 9'b110010110;
assign micromatr[31][78] = 9'b110010010;
assign micromatr[31][79] = 9'b110010010;
assign micromatr[31][80] = 9'b110010110;
assign micromatr[31][81] = 9'b110111111;
assign micromatr[31][82] = 9'b111111111;
assign micromatr[31][83] = 9'b111111111;
assign micromatr[31][84] = 9'b111111111;
assign micromatr[31][85] = 9'b111111111;
assign micromatr[31][86] = 9'b111111111;
assign micromatr[31][87] = 9'b111111111;
assign micromatr[31][88] = 9'b111111111;
assign micromatr[31][89] = 9'b111111111;
assign micromatr[31][90] = 9'b111111111;
assign micromatr[31][91] = 9'b111111111;
assign micromatr[31][92] = 9'b111111111;
assign micromatr[31][93] = 9'b111111111;
assign micromatr[31][94] = 9'b111111111;
assign micromatr[31][95] = 9'b111111111;
assign micromatr[31][96] = 9'b111111111;
assign micromatr[31][97] = 9'b111111111;
assign micromatr[31][98] = 9'b111111111;
assign micromatr[31][99] = 9'b111111111;
assign micromatr[32][0] = 9'b111111111;
assign micromatr[32][1] = 9'b111111111;
assign micromatr[32][2] = 9'b111111111;
assign micromatr[32][3] = 9'b111111111;
assign micromatr[32][4] = 9'b111111111;
assign micromatr[32][5] = 9'b111111111;
assign micromatr[32][6] = 9'b111111111;
assign micromatr[32][7] = 9'b111111111;
assign micromatr[32][8] = 9'b111111111;
assign micromatr[32][9] = 9'b111111111;
assign micromatr[32][10] = 9'b111111111;
assign micromatr[32][11] = 9'b111111111;
assign micromatr[32][12] = 9'b111111111;
assign micromatr[32][13] = 9'b111111111;
assign micromatr[32][14] = 9'b111111111;
assign micromatr[32][15] = 9'b111111111;
assign micromatr[32][16] = 9'b110010001;
assign micromatr[32][17] = 9'b110001101;
assign micromatr[32][18] = 9'b110110010;
assign micromatr[32][19] = 9'b110001101;
assign micromatr[32][20] = 9'b110110010;
assign micromatr[32][21] = 9'b111111111;
assign micromatr[32][22] = 9'b110111110;
assign micromatr[32][23] = 9'b110110010;
assign micromatr[32][24] = 9'b111110110;
assign micromatr[32][25] = 9'b111110010;
assign micromatr[32][26] = 9'b110110010;
assign micromatr[32][27] = 9'b111111111;
assign micromatr[32][28] = 9'b111111111;
assign micromatr[32][29] = 9'b110110110;
assign micromatr[32][30] = 9'b101101101;
assign micromatr[32][31] = 9'b110001110;
assign micromatr[32][32] = 9'b111110111;
assign micromatr[32][33] = 9'b110001110;
assign micromatr[32][34] = 9'b110110010;
assign micromatr[32][35] = 9'b111111111;
assign micromatr[32][36] = 9'b111111111;
assign micromatr[32][37] = 9'b111111111;
assign micromatr[32][38] = 9'b110001101;
assign micromatr[32][39] = 9'b110001110;
assign micromatr[32][40] = 9'b110001101;
assign micromatr[32][41] = 9'b110110010;
assign micromatr[32][42] = 9'b111111111;
assign micromatr[32][43] = 9'b111111111;
assign micromatr[32][44] = 9'b110010001;
assign micromatr[32][45] = 9'b110010010;
assign micromatr[32][46] = 9'b110010110;
assign micromatr[32][47] = 9'b110010110;
assign micromatr[32][48] = 9'b110010110;
assign micromatr[32][49] = 9'b110010110;
assign micromatr[32][50] = 9'b110010110;
assign micromatr[32][51] = 9'b111111111;
assign micromatr[32][52] = 9'b111111111;
assign micromatr[32][53] = 9'b110010010;
assign micromatr[32][54] = 9'b110010001;
assign micromatr[32][55] = 9'b110110010;
assign micromatr[32][56] = 9'b110110010;
assign micromatr[32][57] = 9'b110110010;
assign micromatr[32][58] = 9'b110110010;
assign micromatr[32][59] = 9'b111110010;
assign micromatr[32][60] = 9'b110110010;
assign micromatr[32][61] = 9'b110110010;
assign micromatr[32][62] = 9'b111110010;
assign micromatr[32][63] = 9'b111111111;
assign micromatr[32][64] = 9'b111110111;
assign micromatr[32][65] = 9'b101101101;
assign micromatr[32][66] = 9'b110010010;
assign micromatr[32][67] = 9'b110010010;
assign micromatr[32][68] = 9'b110010010;
assign micromatr[32][69] = 9'b110010010;
assign micromatr[32][70] = 9'b110010010;
assign micromatr[32][71] = 9'b111111111;
assign micromatr[32][72] = 9'b111111111;
assign micromatr[32][73] = 9'b110110110;
assign micromatr[32][74] = 9'b110010001;
assign micromatr[32][75] = 9'b110010010;
assign micromatr[32][76] = 9'b111111111;
assign micromatr[32][77] = 9'b111111111;
assign micromatr[32][78] = 9'b111111111;
assign micromatr[32][79] = 9'b111111111;
assign micromatr[32][80] = 9'b111111111;
assign micromatr[32][81] = 9'b111111111;
assign micromatr[32][82] = 9'b111111111;
assign micromatr[32][83] = 9'b111111111;
assign micromatr[32][84] = 9'b111111111;
assign micromatr[32][85] = 9'b111111111;
assign micromatr[32][86] = 9'b111111111;
assign micromatr[32][87] = 9'b111111111;
assign micromatr[32][88] = 9'b111111111;
assign micromatr[32][89] = 9'b111111111;
assign micromatr[32][90] = 9'b111111111;
assign micromatr[32][91] = 9'b111111111;
assign micromatr[32][92] = 9'b111111111;
assign micromatr[32][93] = 9'b111111111;
assign micromatr[32][94] = 9'b111111111;
assign micromatr[32][95] = 9'b111111111;
assign micromatr[32][96] = 9'b111111111;
assign micromatr[32][97] = 9'b111111111;
assign micromatr[32][98] = 9'b111111111;
assign micromatr[32][99] = 9'b111111111;
assign micromatr[33][0] = 9'b111111111;
assign micromatr[33][1] = 9'b111111111;
assign micromatr[33][2] = 9'b111111111;
assign micromatr[33][3] = 9'b111111111;
assign micromatr[33][4] = 9'b111111111;
assign micromatr[33][5] = 9'b111111111;
assign micromatr[33][6] = 9'b111111111;
assign micromatr[33][7] = 9'b111111111;
assign micromatr[33][8] = 9'b111111111;
assign micromatr[33][9] = 9'b111111111;
assign micromatr[33][10] = 9'b111111111;
assign micromatr[33][11] = 9'b111111111;
assign micromatr[33][12] = 9'b111111111;
assign micromatr[33][13] = 9'b111111111;
assign micromatr[33][14] = 9'b111111111;
assign micromatr[33][15] = 9'b111111111;
assign micromatr[33][16] = 9'b111111111;
assign micromatr[33][17] = 9'b111111111;
assign micromatr[33][18] = 9'b110110110;
assign micromatr[33][19] = 9'b110010010;
assign micromatr[33][20] = 9'b111111111;
assign micromatr[33][21] = 9'b111111111;
assign micromatr[33][22] = 9'b111111111;
assign micromatr[33][23] = 9'b111111111;
assign micromatr[33][24] = 9'b111111111;
assign micromatr[33][25] = 9'b111111111;
assign micromatr[33][26] = 9'b111111111;
assign micromatr[33][27] = 9'b111111111;
assign micromatr[33][28] = 9'b111111111;
assign micromatr[33][29] = 9'b111111111;
assign micromatr[33][30] = 9'b111111111;
assign micromatr[33][31] = 9'b110010010;
assign micromatr[33][32] = 9'b101101101;
assign micromatr[33][33] = 9'b110001110;
assign micromatr[33][34] = 9'b111111111;
assign micromatr[33][35] = 9'b111110111;
assign micromatr[33][36] = 9'b111111111;
assign micromatr[33][37] = 9'b111111111;
assign micromatr[33][38] = 9'b111111111;
assign micromatr[33][39] = 9'b110010001;
assign micromatr[33][40] = 9'b111111111;
assign micromatr[33][41] = 9'b111111111;
assign micromatr[33][42] = 9'b111110111;
assign micromatr[33][43] = 9'b111111111;
assign micromatr[33][44] = 9'b111111111;
assign micromatr[33][45] = 9'b111111111;
assign micromatr[33][46] = 9'b110110110;
assign micromatr[33][47] = 9'b111111111;
assign micromatr[33][48] = 9'b111111111;
assign micromatr[33][49] = 9'b111111111;
assign micromatr[33][50] = 9'b111111111;
assign micromatr[33][51] = 9'b111111111;
assign micromatr[33][52] = 9'b111111111;
assign micromatr[33][53] = 9'b111111111;
assign micromatr[33][54] = 9'b111111111;
assign micromatr[33][55] = 9'b111111111;
assign micromatr[33][56] = 9'b111111111;
assign micromatr[33][57] = 9'b111111111;
assign micromatr[33][58] = 9'b111111111;
assign micromatr[33][59] = 9'b111111111;
assign micromatr[33][60] = 9'b111111111;
assign micromatr[33][61] = 9'b111111111;
assign micromatr[33][62] = 9'b111111111;
assign micromatr[33][63] = 9'b111111111;
assign micromatr[33][64] = 9'b111111111;
assign micromatr[33][65] = 9'b111111111;
assign micromatr[33][66] = 9'b110110110;
assign micromatr[33][67] = 9'b111111111;
assign micromatr[33][68] = 9'b111111111;
assign micromatr[33][69] = 9'b111111111;
assign micromatr[33][70] = 9'b111111111;
assign micromatr[33][71] = 9'b111111111;
assign micromatr[33][72] = 9'b111110111;
assign micromatr[33][73] = 9'b111111111;
assign micromatr[33][74] = 9'b111111111;
assign micromatr[33][75] = 9'b111111111;
assign micromatr[33][76] = 9'b111111111;
assign micromatr[33][77] = 9'b111111111;
assign micromatr[33][78] = 9'b111111111;
assign micromatr[33][79] = 9'b111111111;
assign micromatr[33][80] = 9'b111111111;
assign micromatr[33][81] = 9'b111111111;
assign micromatr[33][82] = 9'b111111111;
assign micromatr[33][83] = 9'b111111111;
assign micromatr[33][84] = 9'b111111111;
assign micromatr[33][85] = 9'b111111111;
assign micromatr[33][86] = 9'b111111111;
assign micromatr[33][87] = 9'b111111111;
assign micromatr[33][88] = 9'b111111111;
assign micromatr[33][89] = 9'b111111111;
assign micromatr[33][90] = 9'b111111111;
assign micromatr[33][91] = 9'b111111111;
assign micromatr[33][92] = 9'b111111111;
assign micromatr[33][93] = 9'b111111111;
assign micromatr[33][94] = 9'b111111111;
assign micromatr[33][95] = 9'b111111111;
assign micromatr[33][96] = 9'b111111111;
assign micromatr[33][97] = 9'b111111111;
assign micromatr[33][98] = 9'b111111111;
assign micromatr[33][99] = 9'b111111111;
assign micromatr[34][0] = 9'b111111111;
assign micromatr[34][1] = 9'b111111111;
assign micromatr[34][2] = 9'b111111111;
assign micromatr[34][3] = 9'b111111111;
assign micromatr[34][4] = 9'b111111111;
assign micromatr[34][5] = 9'b111111111;
assign micromatr[34][6] = 9'b111111111;
assign micromatr[34][7] = 9'b111111111;
assign micromatr[34][8] = 9'b111111111;
assign micromatr[34][9] = 9'b111111111;
assign micromatr[34][10] = 9'b111111111;
assign micromatr[34][11] = 9'b111111111;
assign micromatr[34][12] = 9'b111111111;
assign micromatr[34][13] = 9'b111111111;
assign micromatr[34][14] = 9'b111111111;
assign micromatr[34][15] = 9'b111111111;
assign micromatr[34][16] = 9'b111111111;
assign micromatr[34][17] = 9'b111111111;
assign micromatr[34][18] = 9'b111111111;
assign micromatr[34][19] = 9'b111111111;
assign micromatr[34][20] = 9'b111111111;
assign micromatr[34][21] = 9'b111111111;
assign micromatr[34][22] = 9'b111111111;
assign micromatr[34][23] = 9'b111111111;
assign micromatr[34][24] = 9'b111111111;
assign micromatr[34][25] = 9'b111111111;
assign micromatr[34][26] = 9'b111111111;
assign micromatr[34][27] = 9'b111111111;
assign micromatr[34][28] = 9'b111111111;
assign micromatr[34][29] = 9'b111111111;
assign micromatr[34][30] = 9'b111111111;
assign micromatr[34][31] = 9'b111111111;
assign micromatr[34][32] = 9'b111111111;
assign micromatr[34][33] = 9'b111111111;
assign micromatr[34][34] = 9'b111110111;
assign micromatr[34][35] = 9'b111111111;
assign micromatr[34][36] = 9'b111111111;
assign micromatr[34][37] = 9'b111111111;
assign micromatr[34][38] = 9'b111111111;
assign micromatr[34][39] = 9'b111111111;
assign micromatr[34][40] = 9'b110110111;
assign micromatr[34][41] = 9'b111111111;
assign micromatr[34][42] = 9'b111111111;
assign micromatr[34][43] = 9'b111111111;
assign micromatr[34][44] = 9'b111111111;
assign micromatr[34][45] = 9'b111111111;
assign micromatr[34][46] = 9'b111111111;
assign micromatr[34][47] = 9'b111111111;
assign micromatr[34][48] = 9'b111111111;
assign micromatr[34][49] = 9'b111111111;
assign micromatr[34][50] = 9'b111111111;
assign micromatr[34][51] = 9'b111111111;
assign micromatr[34][52] = 9'b111111111;
assign micromatr[34][53] = 9'b111111111;
assign micromatr[34][54] = 9'b111111111;
assign micromatr[34][55] = 9'b111111111;
assign micromatr[34][56] = 9'b111111111;
assign micromatr[34][57] = 9'b111111111;
assign micromatr[34][58] = 9'b111111111;
assign micromatr[34][59] = 9'b111111111;
assign micromatr[34][60] = 9'b111111111;
assign micromatr[34][61] = 9'b111111111;
assign micromatr[34][62] = 9'b111111111;
assign micromatr[34][63] = 9'b111111111;
assign micromatr[34][64] = 9'b111111111;
assign micromatr[34][65] = 9'b111111111;
assign micromatr[34][66] = 9'b111111111;
assign micromatr[34][67] = 9'b111111111;
assign micromatr[34][68] = 9'b111111111;
assign micromatr[34][69] = 9'b111111111;
assign micromatr[34][70] = 9'b111111111;
assign micromatr[34][71] = 9'b111111111;
assign micromatr[34][72] = 9'b111111111;
assign micromatr[34][73] = 9'b111111111;
assign micromatr[34][74] = 9'b111111111;
assign micromatr[34][75] = 9'b111111111;
assign micromatr[34][76] = 9'b111111111;
assign micromatr[34][77] = 9'b111111111;
assign micromatr[34][78] = 9'b111111111;
assign micromatr[34][79] = 9'b111111111;
assign micromatr[34][80] = 9'b111111111;
assign micromatr[34][81] = 9'b111111111;
assign micromatr[34][82] = 9'b111111111;
assign micromatr[34][83] = 9'b111111111;
assign micromatr[34][84] = 9'b111111111;
assign micromatr[34][85] = 9'b111111111;
assign micromatr[34][86] = 9'b111111111;
assign micromatr[34][87] = 9'b111111111;
assign micromatr[34][88] = 9'b111111111;
assign micromatr[34][89] = 9'b111111111;
assign micromatr[34][90] = 9'b111111111;
assign micromatr[34][91] = 9'b111111111;
assign micromatr[34][92] = 9'b111111111;
assign micromatr[34][93] = 9'b111111111;
assign micromatr[34][94] = 9'b111111111;
assign micromatr[34][95] = 9'b111111111;
assign micromatr[34][96] = 9'b111111111;
assign micromatr[34][97] = 9'b111111111;
assign micromatr[34][98] = 9'b111111111;
assign micromatr[34][99] = 9'b111111111;
assign micromatr[35][0] = 9'b111111111;
assign micromatr[35][1] = 9'b111111111;
assign micromatr[35][2] = 9'b111111111;
assign micromatr[35][3] = 9'b111111111;
assign micromatr[35][4] = 9'b111111111;
assign micromatr[35][5] = 9'b111111111;
assign micromatr[35][6] = 9'b111111111;
assign micromatr[35][7] = 9'b111111111;
assign micromatr[35][8] = 9'b111111111;
assign micromatr[35][9] = 9'b111111111;
assign micromatr[35][10] = 9'b111111111;
assign micromatr[35][11] = 9'b111111111;
assign micromatr[35][12] = 9'b111111111;
assign micromatr[35][13] = 9'b111111111;
assign micromatr[35][14] = 9'b111111111;
assign micromatr[35][15] = 9'b111111111;
assign micromatr[35][16] = 9'b111111111;
assign micromatr[35][17] = 9'b111111111;
assign micromatr[35][18] = 9'b111111111;
assign micromatr[35][19] = 9'b111111111;
assign micromatr[35][20] = 9'b111111111;
assign micromatr[35][21] = 9'b111111111;
assign micromatr[35][22] = 9'b111111111;
assign micromatr[35][23] = 9'b111111111;
assign micromatr[35][24] = 9'b111111111;
assign micromatr[35][25] = 9'b111111111;
assign micromatr[35][26] = 9'b111111111;
assign micromatr[35][27] = 9'b111111111;
assign micromatr[35][28] = 9'b111111111;
assign micromatr[35][29] = 9'b111111111;
assign micromatr[35][30] = 9'b111111111;
assign micromatr[35][31] = 9'b111111111;
assign micromatr[35][32] = 9'b111111111;
assign micromatr[35][33] = 9'b111111111;
assign micromatr[35][34] = 9'b111111111;
assign micromatr[35][35] = 9'b111111111;
assign micromatr[35][36] = 9'b111111111;
assign micromatr[35][37] = 9'b111111111;
assign micromatr[35][38] = 9'b111111111;
assign micromatr[35][39] = 9'b111111111;
assign micromatr[35][40] = 9'b111111111;
assign micromatr[35][41] = 9'b111111111;
assign micromatr[35][42] = 9'b111111111;
assign micromatr[35][43] = 9'b111111111;
assign micromatr[35][44] = 9'b111111111;
assign micromatr[35][45] = 9'b111111111;
assign micromatr[35][46] = 9'b111111111;
assign micromatr[35][47] = 9'b111111111;
assign micromatr[35][48] = 9'b111111111;
assign micromatr[35][49] = 9'b111111111;
assign micromatr[35][50] = 9'b111111111;
assign micromatr[35][51] = 9'b111111111;
assign micromatr[35][52] = 9'b111111111;
assign micromatr[35][53] = 9'b111111111;
assign micromatr[35][54] = 9'b111111111;
assign micromatr[35][55] = 9'b111111111;
assign micromatr[35][56] = 9'b111111111;
assign micromatr[35][57] = 9'b111111111;
assign micromatr[35][58] = 9'b111111111;
assign micromatr[35][59] = 9'b111111111;
assign micromatr[35][60] = 9'b111111111;
assign micromatr[35][61] = 9'b111111111;
assign micromatr[35][62] = 9'b111111111;
assign micromatr[35][63] = 9'b111111111;
assign micromatr[35][64] = 9'b111111111;
assign micromatr[35][65] = 9'b111111111;
assign micromatr[35][66] = 9'b111111111;
assign micromatr[35][67] = 9'b111111111;
assign micromatr[35][68] = 9'b111111111;
assign micromatr[35][69] = 9'b111111111;
assign micromatr[35][70] = 9'b111111111;
assign micromatr[35][71] = 9'b111111111;
assign micromatr[35][72] = 9'b111111111;
assign micromatr[35][73] = 9'b111111111;
assign micromatr[35][74] = 9'b111111111;
assign micromatr[35][75] = 9'b111111111;
assign micromatr[35][76] = 9'b111111111;
assign micromatr[35][77] = 9'b111111111;
assign micromatr[35][78] = 9'b111111111;
assign micromatr[35][79] = 9'b111111111;
assign micromatr[35][80] = 9'b111111111;
assign micromatr[35][81] = 9'b111111111;
assign micromatr[35][82] = 9'b111111111;
assign micromatr[35][83] = 9'b111111111;
assign micromatr[35][84] = 9'b111111111;
assign micromatr[35][85] = 9'b111111111;
assign micromatr[35][86] = 9'b111111111;
assign micromatr[35][87] = 9'b111111111;
assign micromatr[35][88] = 9'b111111111;
assign micromatr[35][89] = 9'b111111111;
assign micromatr[35][90] = 9'b111111111;
assign micromatr[35][91] = 9'b111111111;
assign micromatr[35][92] = 9'b111111111;
assign micromatr[35][93] = 9'b111111111;
assign micromatr[35][94] = 9'b111111111;
assign micromatr[35][95] = 9'b111111111;
assign micromatr[35][96] = 9'b111111111;
assign micromatr[35][97] = 9'b111111111;
assign micromatr[35][98] = 9'b111111111;
assign micromatr[35][99] = 9'b111111111;
assign micromatr[36][0] = 9'b111111111;
assign micromatr[36][1] = 9'b111111111;
assign micromatr[36][2] = 9'b111111111;
assign micromatr[36][3] = 9'b111111111;
assign micromatr[36][4] = 9'b111111111;
assign micromatr[36][5] = 9'b111111111;
assign micromatr[36][6] = 9'b111111111;
assign micromatr[36][7] = 9'b111111111;
assign micromatr[36][8] = 9'b111111111;
assign micromatr[36][9] = 9'b111111111;
assign micromatr[36][10] = 9'b111111111;
assign micromatr[36][11] = 9'b111111111;
assign micromatr[36][12] = 9'b111111111;
assign micromatr[36][13] = 9'b111111111;
assign micromatr[36][14] = 9'b111111111;
assign micromatr[36][15] = 9'b111111111;
assign micromatr[36][16] = 9'b111111111;
assign micromatr[36][17] = 9'b111111111;
assign micromatr[36][18] = 9'b111111111;
assign micromatr[36][19] = 9'b111111111;
assign micromatr[36][20] = 9'b111111111;
assign micromatr[36][21] = 9'b111111111;
assign micromatr[36][22] = 9'b111111111;
assign micromatr[36][23] = 9'b111111111;
assign micromatr[36][24] = 9'b111111111;
assign micromatr[36][25] = 9'b111111111;
assign micromatr[36][26] = 9'b111111111;
assign micromatr[36][27] = 9'b111111111;
assign micromatr[36][28] = 9'b111111111;
assign micromatr[36][29] = 9'b111111111;
assign micromatr[36][30] = 9'b111111111;
assign micromatr[36][31] = 9'b111111111;
assign micromatr[36][32] = 9'b111111111;
assign micromatr[36][33] = 9'b111111111;
assign micromatr[36][34] = 9'b111111111;
assign micromatr[36][35] = 9'b111111111;
assign micromatr[36][36] = 9'b111111111;
assign micromatr[36][37] = 9'b111111111;
assign micromatr[36][38] = 9'b111111111;
assign micromatr[36][39] = 9'b111111111;
assign micromatr[36][40] = 9'b111111111;
assign micromatr[36][41] = 9'b111111111;
assign micromatr[36][42] = 9'b111111111;
assign micromatr[36][43] = 9'b111111111;
assign micromatr[36][44] = 9'b111111111;
assign micromatr[36][45] = 9'b111111111;
assign micromatr[36][46] = 9'b111111111;
assign micromatr[36][47] = 9'b111111111;
assign micromatr[36][48] = 9'b111111111;
assign micromatr[36][49] = 9'b111111111;
assign micromatr[36][50] = 9'b111111111;
assign micromatr[36][51] = 9'b111111111;
assign micromatr[36][52] = 9'b111111111;
assign micromatr[36][53] = 9'b111111111;
assign micromatr[36][54] = 9'b111111111;
assign micromatr[36][55] = 9'b111111111;
assign micromatr[36][56] = 9'b111111111;
assign micromatr[36][57] = 9'b111111111;
assign micromatr[36][58] = 9'b111111111;
assign micromatr[36][59] = 9'b111111111;
assign micromatr[36][60] = 9'b111111111;
assign micromatr[36][61] = 9'b111111111;
assign micromatr[36][62] = 9'b111111111;
assign micromatr[36][63] = 9'b111111111;
assign micromatr[36][64] = 9'b111111111;
assign micromatr[36][65] = 9'b111111111;
assign micromatr[36][66] = 9'b111111111;
assign micromatr[36][67] = 9'b111111111;
assign micromatr[36][68] = 9'b111111111;
assign micromatr[36][69] = 9'b111111111;
assign micromatr[36][70] = 9'b111111111;
assign micromatr[36][71] = 9'b111111111;
assign micromatr[36][72] = 9'b111111111;
assign micromatr[36][73] = 9'b111111111;
assign micromatr[36][74] = 9'b111111111;
assign micromatr[36][75] = 9'b111111111;
assign micromatr[36][76] = 9'b111111111;
assign micromatr[36][77] = 9'b111111111;
assign micromatr[36][78] = 9'b111111111;
assign micromatr[36][79] = 9'b111111111;
assign micromatr[36][80] = 9'b111111111;
assign micromatr[36][81] = 9'b111111111;
assign micromatr[36][82] = 9'b111111111;
assign micromatr[36][83] = 9'b111111111;
assign micromatr[36][84] = 9'b111111111;
assign micromatr[36][85] = 9'b111111111;
assign micromatr[36][86] = 9'b111111111;
assign micromatr[36][87] = 9'b111111111;
assign micromatr[36][88] = 9'b111111111;
assign micromatr[36][89] = 9'b111111111;
assign micromatr[36][90] = 9'b111111111;
assign micromatr[36][91] = 9'b111111111;
assign micromatr[36][92] = 9'b111111111;
assign micromatr[36][93] = 9'b111111111;
assign micromatr[36][94] = 9'b111111111;
assign micromatr[36][95] = 9'b111111111;
assign micromatr[36][96] = 9'b111111111;
assign micromatr[36][97] = 9'b111111111;
assign micromatr[36][98] = 9'b111111111;
assign micromatr[36][99] = 9'b111111111;
assign micromatr[37][0] = 9'b111111111;
assign micromatr[37][1] = 9'b111111111;
assign micromatr[37][2] = 9'b111111111;
assign micromatr[37][3] = 9'b111111111;
assign micromatr[37][4] = 9'b111111111;
assign micromatr[37][5] = 9'b111111111;
assign micromatr[37][6] = 9'b111111111;
assign micromatr[37][7] = 9'b111111111;
assign micromatr[37][8] = 9'b111111111;
assign micromatr[37][9] = 9'b111111111;
assign micromatr[37][10] = 9'b111111111;
assign micromatr[37][11] = 9'b111111111;
assign micromatr[37][12] = 9'b111111111;
assign micromatr[37][13] = 9'b111111111;
assign micromatr[37][14] = 9'b111111111;
assign micromatr[37][15] = 9'b111111111;
assign micromatr[37][16] = 9'b111111111;
assign micromatr[37][17] = 9'b111111111;
assign micromatr[37][18] = 9'b111111111;
assign micromatr[37][19] = 9'b111111111;
assign micromatr[37][20] = 9'b111111111;
assign micromatr[37][21] = 9'b111111111;
assign micromatr[37][22] = 9'b111111111;
assign micromatr[37][23] = 9'b111111111;
assign micromatr[37][24] = 9'b111111111;
assign micromatr[37][25] = 9'b111111111;
assign micromatr[37][26] = 9'b111111111;
assign micromatr[37][27] = 9'b111111111;
assign micromatr[37][28] = 9'b111111111;
assign micromatr[37][29] = 9'b111111111;
assign micromatr[37][30] = 9'b111111111;
assign micromatr[37][31] = 9'b111111111;
assign micromatr[37][32] = 9'b111111111;
assign micromatr[37][33] = 9'b111111111;
assign micromatr[37][34] = 9'b111111111;
assign micromatr[37][35] = 9'b111111111;
assign micromatr[37][36] = 9'b111111111;
assign micromatr[37][37] = 9'b111111111;
assign micromatr[37][38] = 9'b111111111;
assign micromatr[37][39] = 9'b111111111;
assign micromatr[37][40] = 9'b111111111;
assign micromatr[37][41] = 9'b111111111;
assign micromatr[37][42] = 9'b111111111;
assign micromatr[37][43] = 9'b111111111;
assign micromatr[37][44] = 9'b111111111;
assign micromatr[37][45] = 9'b111111111;
assign micromatr[37][46] = 9'b111111111;
assign micromatr[37][47] = 9'b111111111;
assign micromatr[37][48] = 9'b111111111;
assign micromatr[37][49] = 9'b111111111;
assign micromatr[37][50] = 9'b111111111;
assign micromatr[37][51] = 9'b111111111;
assign micromatr[37][52] = 9'b111111111;
assign micromatr[37][53] = 9'b111111111;
assign micromatr[37][54] = 9'b111111111;
assign micromatr[37][55] = 9'b111111111;
assign micromatr[37][56] = 9'b111111111;
assign micromatr[37][57] = 9'b111111111;
assign micromatr[37][58] = 9'b111111111;
assign micromatr[37][59] = 9'b111111111;
assign micromatr[37][60] = 9'b111111111;
assign micromatr[37][61] = 9'b111111111;
assign micromatr[37][62] = 9'b111111111;
assign micromatr[37][63] = 9'b111111111;
assign micromatr[37][64] = 9'b111111111;
assign micromatr[37][65] = 9'b111111111;
assign micromatr[37][66] = 9'b111111111;
assign micromatr[37][67] = 9'b111111111;
assign micromatr[37][68] = 9'b111111111;
assign micromatr[37][69] = 9'b111111111;
assign micromatr[37][70] = 9'b111111111;
assign micromatr[37][71] = 9'b111111111;
assign micromatr[37][72] = 9'b111111111;
assign micromatr[37][73] = 9'b111111111;
assign micromatr[37][74] = 9'b111111111;
assign micromatr[37][75] = 9'b111111111;
assign micromatr[37][76] = 9'b111111111;
assign micromatr[37][77] = 9'b111111111;
assign micromatr[37][78] = 9'b111111111;
assign micromatr[37][79] = 9'b111111111;
assign micromatr[37][80] = 9'b111111111;
assign micromatr[37][81] = 9'b111111111;
assign micromatr[37][82] = 9'b111111111;
assign micromatr[37][83] = 9'b111111111;
assign micromatr[37][84] = 9'b111111111;
assign micromatr[37][85] = 9'b111111111;
assign micromatr[37][86] = 9'b111111111;
assign micromatr[37][87] = 9'b111111111;
assign micromatr[37][88] = 9'b111111111;
assign micromatr[37][89] = 9'b111111111;
assign micromatr[37][90] = 9'b111111111;
assign micromatr[37][91] = 9'b111111111;
assign micromatr[37][92] = 9'b111111111;
assign micromatr[37][93] = 9'b111111111;
assign micromatr[37][94] = 9'b111111111;
assign micromatr[37][95] = 9'b111111111;
assign micromatr[37][96] = 9'b111111111;
assign micromatr[37][97] = 9'b111111111;
assign micromatr[37][98] = 9'b111111111;
assign micromatr[37][99] = 9'b111111111;
assign micromatr[38][0] = 9'b111111111;
assign micromatr[38][1] = 9'b111111111;
assign micromatr[38][2] = 9'b111111111;
assign micromatr[38][3] = 9'b111111111;
assign micromatr[38][4] = 9'b111111111;
assign micromatr[38][5] = 9'b111111111;
assign micromatr[38][6] = 9'b111111111;
assign micromatr[38][7] = 9'b111111111;
assign micromatr[38][8] = 9'b111111111;
assign micromatr[38][9] = 9'b111111111;
assign micromatr[38][10] = 9'b111111111;
assign micromatr[38][11] = 9'b111111111;
assign micromatr[38][12] = 9'b111111111;
assign micromatr[38][13] = 9'b111111111;
assign micromatr[38][14] = 9'b111111111;
assign micromatr[38][15] = 9'b111111111;
assign micromatr[38][16] = 9'b111111111;
assign micromatr[38][17] = 9'b111111111;
assign micromatr[38][18] = 9'b111111111;
assign micromatr[38][19] = 9'b111111111;
assign micromatr[38][20] = 9'b111111111;
assign micromatr[38][21] = 9'b111111111;
assign micromatr[38][22] = 9'b111111111;
assign micromatr[38][23] = 9'b111111111;
assign micromatr[38][24] = 9'b111111111;
assign micromatr[38][25] = 9'b111111111;
assign micromatr[38][26] = 9'b111111111;
assign micromatr[38][27] = 9'b111111111;
assign micromatr[38][28] = 9'b111111111;
assign micromatr[38][29] = 9'b111111111;
assign micromatr[38][30] = 9'b111111111;
assign micromatr[38][31] = 9'b111111111;
assign micromatr[38][32] = 9'b111111111;
assign micromatr[38][33] = 9'b111111111;
assign micromatr[38][34] = 9'b111111111;
assign micromatr[38][35] = 9'b111111111;
assign micromatr[38][36] = 9'b111111111;
assign micromatr[38][37] = 9'b111111111;
assign micromatr[38][38] = 9'b111111111;
assign micromatr[38][39] = 9'b111111111;
assign micromatr[38][40] = 9'b111111111;
assign micromatr[38][41] = 9'b111111111;
assign micromatr[38][42] = 9'b111111111;
assign micromatr[38][43] = 9'b111111111;
assign micromatr[38][44] = 9'b111111111;
assign micromatr[38][45] = 9'b111111111;
assign micromatr[38][46] = 9'b111111111;
assign micromatr[38][47] = 9'b111111111;
assign micromatr[38][48] = 9'b111111111;
assign micromatr[38][49] = 9'b111111111;
assign micromatr[38][50] = 9'b111111111;
assign micromatr[38][51] = 9'b111111111;
assign micromatr[38][52] = 9'b111111111;
assign micromatr[38][53] = 9'b111111111;
assign micromatr[38][54] = 9'b111111111;
assign micromatr[38][55] = 9'b111111111;
assign micromatr[38][56] = 9'b111111111;
assign micromatr[38][57] = 9'b111111111;
assign micromatr[38][58] = 9'b111111111;
assign micromatr[38][59] = 9'b111111111;
assign micromatr[38][60] = 9'b111111111;
assign micromatr[38][61] = 9'b111111111;
assign micromatr[38][62] = 9'b111111111;
assign micromatr[38][63] = 9'b111111111;
assign micromatr[38][64] = 9'b111111111;
assign micromatr[38][65] = 9'b111111111;
assign micromatr[38][66] = 9'b111111111;
assign micromatr[38][67] = 9'b111111111;
assign micromatr[38][68] = 9'b111111111;
assign micromatr[38][69] = 9'b111111111;
assign micromatr[38][70] = 9'b111111111;
assign micromatr[38][71] = 9'b111111111;
assign micromatr[38][72] = 9'b111111111;
assign micromatr[38][73] = 9'b111111111;
assign micromatr[38][74] = 9'b111111111;
assign micromatr[38][75] = 9'b111111111;
assign micromatr[38][76] = 9'b111111111;
assign micromatr[38][77] = 9'b111111111;
assign micromatr[38][78] = 9'b111111111;
assign micromatr[38][79] = 9'b111111111;
assign micromatr[38][80] = 9'b111111111;
assign micromatr[38][81] = 9'b111111111;
assign micromatr[38][82] = 9'b111111111;
assign micromatr[38][83] = 9'b111111111;
assign micromatr[38][84] = 9'b111111111;
assign micromatr[38][85] = 9'b111111111;
assign micromatr[38][86] = 9'b111111111;
assign micromatr[38][87] = 9'b111111111;
assign micromatr[38][88] = 9'b111111111;
assign micromatr[38][89] = 9'b111111111;
assign micromatr[38][90] = 9'b111111111;
assign micromatr[38][91] = 9'b111111111;
assign micromatr[38][92] = 9'b111111111;
assign micromatr[38][93] = 9'b111111111;
assign micromatr[38][94] = 9'b111111111;
assign micromatr[38][95] = 9'b111111111;
assign micromatr[38][96] = 9'b111111111;
assign micromatr[38][97] = 9'b111111111;
assign micromatr[38][98] = 9'b111111111;
assign micromatr[38][99] = 9'b111111111;
assign micromatr[39][0] = 9'b111111111;
assign micromatr[39][1] = 9'b111111111;
assign micromatr[39][2] = 9'b111111111;
assign micromatr[39][3] = 9'b111111111;
assign micromatr[39][4] = 9'b111111111;
assign micromatr[39][5] = 9'b111111111;
assign micromatr[39][6] = 9'b111111111;
assign micromatr[39][7] = 9'b111111111;
assign micromatr[39][8] = 9'b111111111;
assign micromatr[39][9] = 9'b111111111;
assign micromatr[39][10] = 9'b111111111;
assign micromatr[39][11] = 9'b111111111;
assign micromatr[39][12] = 9'b111111111;
assign micromatr[39][13] = 9'b111111111;
assign micromatr[39][14] = 9'b111111111;
assign micromatr[39][15] = 9'b111111111;
assign micromatr[39][16] = 9'b111111111;
assign micromatr[39][17] = 9'b111111111;
assign micromatr[39][18] = 9'b111111111;
assign micromatr[39][19] = 9'b111111111;
assign micromatr[39][20] = 9'b111111111;
assign micromatr[39][21] = 9'b111111111;
assign micromatr[39][22] = 9'b111111111;
assign micromatr[39][23] = 9'b111111111;
assign micromatr[39][24] = 9'b111111111;
assign micromatr[39][25] = 9'b111111111;
assign micromatr[39][26] = 9'b111111111;
assign micromatr[39][27] = 9'b111111111;
assign micromatr[39][28] = 9'b111111111;
assign micromatr[39][29] = 9'b111111111;
assign micromatr[39][30] = 9'b111111111;
assign micromatr[39][31] = 9'b111111111;
assign micromatr[39][32] = 9'b111111111;
assign micromatr[39][33] = 9'b111111111;
assign micromatr[39][34] = 9'b111111111;
assign micromatr[39][35] = 9'b111111111;
assign micromatr[39][36] = 9'b111111111;
assign micromatr[39][37] = 9'b111111111;
assign micromatr[39][38] = 9'b111111111;
assign micromatr[39][39] = 9'b111111111;
assign micromatr[39][40] = 9'b111111111;
assign micromatr[39][41] = 9'b111111111;
assign micromatr[39][42] = 9'b111111111;
assign micromatr[39][43] = 9'b111111111;
assign micromatr[39][44] = 9'b111111111;
assign micromatr[39][45] = 9'b111111111;
assign micromatr[39][46] = 9'b111111111;
assign micromatr[39][47] = 9'b111111111;
assign micromatr[39][48] = 9'b111111111;
assign micromatr[39][49] = 9'b111111111;
assign micromatr[39][50] = 9'b111111111;
assign micromatr[39][51] = 9'b111111111;
assign micromatr[39][52] = 9'b111111111;
assign micromatr[39][53] = 9'b111111111;
assign micromatr[39][54] = 9'b111111111;
assign micromatr[39][55] = 9'b111111111;
assign micromatr[39][56] = 9'b111111111;
assign micromatr[39][57] = 9'b111111111;
assign micromatr[39][58] = 9'b111111111;
assign micromatr[39][59] = 9'b111111111;
assign micromatr[39][60] = 9'b111111111;
assign micromatr[39][61] = 9'b111111111;
assign micromatr[39][62] = 9'b111111111;
assign micromatr[39][63] = 9'b111111111;
assign micromatr[39][64] = 9'b111111111;
assign micromatr[39][65] = 9'b111111111;
assign micromatr[39][66] = 9'b111111111;
assign micromatr[39][67] = 9'b111111111;
assign micromatr[39][68] = 9'b111111111;
assign micromatr[39][69] = 9'b111111111;
assign micromatr[39][70] = 9'b111111111;
assign micromatr[39][71] = 9'b111111111;
assign micromatr[39][72] = 9'b111111111;
assign micromatr[39][73] = 9'b111111111;
assign micromatr[39][74] = 9'b111111111;
assign micromatr[39][75] = 9'b111111111;
assign micromatr[39][76] = 9'b111111111;
assign micromatr[39][77] = 9'b111111111;
assign micromatr[39][78] = 9'b111111111;
assign micromatr[39][79] = 9'b111111111;
assign micromatr[39][80] = 9'b111111111;
assign micromatr[39][81] = 9'b111111111;
assign micromatr[39][82] = 9'b111111111;
assign micromatr[39][83] = 9'b111111111;
assign micromatr[39][84] = 9'b111111111;
assign micromatr[39][85] = 9'b111111111;
assign micromatr[39][86] = 9'b111111111;
assign micromatr[39][87] = 9'b111111111;
assign micromatr[39][88] = 9'b111111111;
assign micromatr[39][89] = 9'b111111111;
assign micromatr[39][90] = 9'b111111111;
assign micromatr[39][91] = 9'b111111111;
assign micromatr[39][92] = 9'b111111111;
assign micromatr[39][93] = 9'b111111111;
assign micromatr[39][94] = 9'b111111111;
assign micromatr[39][95] = 9'b111111111;
assign micromatr[39][96] = 9'b111111111;
assign micromatr[39][97] = 9'b111111111;
assign micromatr[39][98] = 9'b111111111;
assign micromatr[39][99] = 9'b111111111;
assign micromatr[40][0] = 9'b111111111;
assign micromatr[40][1] = 9'b111111111;
assign micromatr[40][2] = 9'b111111111;
assign micromatr[40][3] = 9'b111111111;
assign micromatr[40][4] = 9'b111111111;
assign micromatr[40][5] = 9'b111111111;
assign micromatr[40][6] = 9'b111111111;
assign micromatr[40][7] = 9'b111111111;
assign micromatr[40][8] = 9'b111111111;
assign micromatr[40][9] = 9'b111111111;
assign micromatr[40][10] = 9'b111111111;
assign micromatr[40][11] = 9'b111111111;
assign micromatr[40][12] = 9'b111111111;
assign micromatr[40][13] = 9'b111111111;
assign micromatr[40][14] = 9'b111111111;
assign micromatr[40][15] = 9'b111111111;
assign micromatr[40][16] = 9'b111111111;
assign micromatr[40][17] = 9'b111111111;
assign micromatr[40][18] = 9'b111111111;
assign micromatr[40][19] = 9'b111111111;
assign micromatr[40][20] = 9'b111111111;
assign micromatr[40][21] = 9'b111111111;
assign micromatr[40][22] = 9'b111111111;
assign micromatr[40][23] = 9'b111111111;
assign micromatr[40][24] = 9'b111111111;
assign micromatr[40][25] = 9'b111111111;
assign micromatr[40][26] = 9'b111111111;
assign micromatr[40][27] = 9'b111111111;
assign micromatr[40][28] = 9'b111111111;
assign micromatr[40][29] = 9'b111111111;
assign micromatr[40][30] = 9'b111111111;
assign micromatr[40][31] = 9'b111111111;
assign micromatr[40][32] = 9'b111111111;
assign micromatr[40][33] = 9'b111111111;
assign micromatr[40][34] = 9'b111111111;
assign micromatr[40][35] = 9'b111111111;
assign micromatr[40][36] = 9'b111111111;
assign micromatr[40][37] = 9'b111111111;
assign micromatr[40][38] = 9'b111111111;
assign micromatr[40][39] = 9'b111111111;
assign micromatr[40][40] = 9'b111111111;
assign micromatr[40][41] = 9'b111111111;
assign micromatr[40][42] = 9'b111111111;
assign micromatr[40][43] = 9'b111111111;
assign micromatr[40][44] = 9'b111111111;
assign micromatr[40][45] = 9'b111111111;
assign micromatr[40][46] = 9'b111111111;
assign micromatr[40][47] = 9'b111111111;
assign micromatr[40][48] = 9'b111111111;
assign micromatr[40][49] = 9'b111111111;
assign micromatr[40][50] = 9'b111111111;
assign micromatr[40][51] = 9'b111111111;
assign micromatr[40][52] = 9'b111111111;
assign micromatr[40][53] = 9'b111111111;
assign micromatr[40][54] = 9'b111111111;
assign micromatr[40][55] = 9'b111111111;
assign micromatr[40][56] = 9'b111111111;
assign micromatr[40][57] = 9'b111111111;
assign micromatr[40][58] = 9'b111111111;
assign micromatr[40][59] = 9'b111111111;
assign micromatr[40][60] = 9'b111111111;
assign micromatr[40][61] = 9'b111111111;
assign micromatr[40][62] = 9'b111111111;
assign micromatr[40][63] = 9'b111111111;
assign micromatr[40][64] = 9'b111111111;
assign micromatr[40][65] = 9'b111111111;
assign micromatr[40][66] = 9'b111111111;
assign micromatr[40][67] = 9'b111111111;
assign micromatr[40][68] = 9'b111111111;
assign micromatr[40][69] = 9'b111111111;
assign micromatr[40][70] = 9'b111111111;
assign micromatr[40][71] = 9'b111111111;
assign micromatr[40][72] = 9'b111111111;
assign micromatr[40][73] = 9'b111111111;
assign micromatr[40][74] = 9'b111111111;
assign micromatr[40][75] = 9'b111111111;
assign micromatr[40][76] = 9'b111111111;
assign micromatr[40][77] = 9'b111111111;
assign micromatr[40][78] = 9'b111111111;
assign micromatr[40][79] = 9'b111111111;
assign micromatr[40][80] = 9'b111111111;
assign micromatr[40][81] = 9'b111111111;
assign micromatr[40][82] = 9'b111111111;
assign micromatr[40][83] = 9'b111111111;
assign micromatr[40][84] = 9'b111111111;
assign micromatr[40][85] = 9'b111111111;
assign micromatr[40][86] = 9'b111111111;
assign micromatr[40][87] = 9'b111111111;
assign micromatr[40][88] = 9'b111111111;
assign micromatr[40][89] = 9'b111111111;
assign micromatr[40][90] = 9'b111111111;
assign micromatr[40][91] = 9'b111111111;
assign micromatr[40][92] = 9'b111111111;
assign micromatr[40][93] = 9'b111111111;
assign micromatr[40][94] = 9'b111111111;
assign micromatr[40][95] = 9'b111111111;
assign micromatr[40][96] = 9'b111111111;
assign micromatr[40][97] = 9'b111111111;
assign micromatr[40][98] = 9'b111111111;
assign micromatr[40][99] = 9'b111111111;
assign micromatr[41][0] = 9'b111111111;
assign micromatr[41][1] = 9'b111111111;
assign micromatr[41][2] = 9'b111111111;
assign micromatr[41][3] = 9'b111111111;
assign micromatr[41][4] = 9'b111111111;
assign micromatr[41][5] = 9'b111111111;
assign micromatr[41][6] = 9'b111111111;
assign micromatr[41][7] = 9'b111111111;
assign micromatr[41][8] = 9'b111111111;
assign micromatr[41][9] = 9'b111111111;
assign micromatr[41][10] = 9'b111111111;
assign micromatr[41][11] = 9'b111111111;
assign micromatr[41][12] = 9'b111111111;
assign micromatr[41][13] = 9'b111111111;
assign micromatr[41][14] = 9'b111111111;
assign micromatr[41][15] = 9'b111111111;
assign micromatr[41][16] = 9'b111111111;
assign micromatr[41][17] = 9'b111111111;
assign micromatr[41][18] = 9'b111111111;
assign micromatr[41][19] = 9'b111111111;
assign micromatr[41][20] = 9'b111111111;
assign micromatr[41][21] = 9'b111111111;
assign micromatr[41][22] = 9'b111111111;
assign micromatr[41][23] = 9'b111111111;
assign micromatr[41][24] = 9'b111111111;
assign micromatr[41][25] = 9'b111111111;
assign micromatr[41][26] = 9'b111111111;
assign micromatr[41][27] = 9'b111111111;
assign micromatr[41][28] = 9'b111111111;
assign micromatr[41][29] = 9'b111111111;
assign micromatr[41][30] = 9'b111111111;
assign micromatr[41][31] = 9'b111111111;
assign micromatr[41][32] = 9'b111111111;
assign micromatr[41][33] = 9'b111111111;
assign micromatr[41][34] = 9'b111111111;
assign micromatr[41][35] = 9'b111111111;
assign micromatr[41][36] = 9'b111111111;
assign micromatr[41][37] = 9'b111111111;
assign micromatr[41][38] = 9'b111111111;
assign micromatr[41][39] = 9'b111111111;
assign micromatr[41][40] = 9'b111111111;
assign micromatr[41][41] = 9'b111111111;
assign micromatr[41][42] = 9'b111111111;
assign micromatr[41][43] = 9'b111111111;
assign micromatr[41][44] = 9'b111111111;
assign micromatr[41][45] = 9'b111111111;
assign micromatr[41][46] = 9'b111111111;
assign micromatr[41][47] = 9'b111111111;
assign micromatr[41][48] = 9'b111111111;
assign micromatr[41][49] = 9'b111111111;
assign micromatr[41][50] = 9'b111111111;
assign micromatr[41][51] = 9'b111111111;
assign micromatr[41][52] = 9'b111111111;
assign micromatr[41][53] = 9'b111111111;
assign micromatr[41][54] = 9'b111111111;
assign micromatr[41][55] = 9'b111111111;
assign micromatr[41][56] = 9'b111111111;
assign micromatr[41][57] = 9'b111111111;
assign micromatr[41][58] = 9'b111111111;
assign micromatr[41][59] = 9'b111111111;
assign micromatr[41][60] = 9'b111111111;
assign micromatr[41][61] = 9'b111111111;
assign micromatr[41][62] = 9'b111111111;
assign micromatr[41][63] = 9'b111111111;
assign micromatr[41][64] = 9'b111111111;
assign micromatr[41][65] = 9'b111111111;
assign micromatr[41][66] = 9'b111111111;
assign micromatr[41][67] = 9'b111111111;
assign micromatr[41][68] = 9'b111111111;
assign micromatr[41][69] = 9'b111111111;
assign micromatr[41][70] = 9'b111111111;
assign micromatr[41][71] = 9'b111111111;
assign micromatr[41][72] = 9'b111111111;
assign micromatr[41][73] = 9'b111111111;
assign micromatr[41][74] = 9'b111111111;
assign micromatr[41][75] = 9'b111111111;
assign micromatr[41][76] = 9'b111111111;
assign micromatr[41][77] = 9'b111111111;
assign micromatr[41][78] = 9'b111111111;
assign micromatr[41][79] = 9'b111111111;
assign micromatr[41][80] = 9'b111111111;
assign micromatr[41][81] = 9'b111111111;
assign micromatr[41][82] = 9'b111111111;
assign micromatr[41][83] = 9'b111111111;
assign micromatr[41][84] = 9'b111111111;
assign micromatr[41][85] = 9'b111111111;
assign micromatr[41][86] = 9'b111111111;
assign micromatr[41][87] = 9'b111111111;
assign micromatr[41][88] = 9'b111111111;
assign micromatr[41][89] = 9'b111111111;
assign micromatr[41][90] = 9'b111111111;
assign micromatr[41][91] = 9'b111111111;
assign micromatr[41][92] = 9'b111111111;
assign micromatr[41][93] = 9'b111111111;
assign micromatr[41][94] = 9'b111111111;
assign micromatr[41][95] = 9'b111111111;
assign micromatr[41][96] = 9'b111111111;
assign micromatr[41][97] = 9'b111111111;
assign micromatr[41][98] = 9'b111111111;
assign micromatr[41][99] = 9'b111111111;
assign micromatr[42][0] = 9'b111111111;
assign micromatr[42][1] = 9'b111111111;
assign micromatr[42][2] = 9'b111111111;
assign micromatr[42][3] = 9'b111111111;
assign micromatr[42][4] = 9'b111111111;
assign micromatr[42][5] = 9'b111111111;
assign micromatr[42][6] = 9'b111111111;
assign micromatr[42][7] = 9'b111111111;
assign micromatr[42][8] = 9'b111111111;
assign micromatr[42][9] = 9'b111111111;
assign micromatr[42][10] = 9'b111111111;
assign micromatr[42][11] = 9'b111111111;
assign micromatr[42][12] = 9'b111111111;
assign micromatr[42][13] = 9'b111111111;
assign micromatr[42][14] = 9'b111111111;
assign micromatr[42][15] = 9'b111111111;
assign micromatr[42][16] = 9'b111111111;
assign micromatr[42][17] = 9'b111111111;
assign micromatr[42][18] = 9'b111111111;
assign micromatr[42][19] = 9'b111111111;
assign micromatr[42][20] = 9'b111111111;
assign micromatr[42][21] = 9'b111111111;
assign micromatr[42][22] = 9'b111111111;
assign micromatr[42][23] = 9'b111111111;
assign micromatr[42][24] = 9'b111111111;
assign micromatr[42][25] = 9'b111111111;
assign micromatr[42][26] = 9'b111111111;
assign micromatr[42][27] = 9'b111111111;
assign micromatr[42][28] = 9'b111111111;
assign micromatr[42][29] = 9'b111111111;
assign micromatr[42][30] = 9'b111111111;
assign micromatr[42][31] = 9'b111111111;
assign micromatr[42][32] = 9'b111111111;
assign micromatr[42][33] = 9'b111111111;
assign micromatr[42][34] = 9'b111111111;
assign micromatr[42][35] = 9'b111111111;
assign micromatr[42][36] = 9'b111111111;
assign micromatr[42][37] = 9'b111111111;
assign micromatr[42][38] = 9'b111111111;
assign micromatr[42][39] = 9'b111111111;
assign micromatr[42][40] = 9'b111111111;
assign micromatr[42][41] = 9'b111111111;
assign micromatr[42][42] = 9'b111111111;
assign micromatr[42][43] = 9'b111111111;
assign micromatr[42][44] = 9'b111111111;
assign micromatr[42][45] = 9'b111111111;
assign micromatr[42][46] = 9'b111111111;
assign micromatr[42][47] = 9'b111111111;
assign micromatr[42][48] = 9'b111111111;
assign micromatr[42][49] = 9'b111111111;
assign micromatr[42][50] = 9'b111111111;
assign micromatr[42][51] = 9'b111111111;
assign micromatr[42][52] = 9'b111111111;
assign micromatr[42][53] = 9'b111111111;
assign micromatr[42][54] = 9'b111111111;
assign micromatr[42][55] = 9'b111111111;
assign micromatr[42][56] = 9'b111111111;
assign micromatr[42][57] = 9'b111111111;
assign micromatr[42][58] = 9'b111111111;
assign micromatr[42][59] = 9'b111111111;
assign micromatr[42][60] = 9'b111111111;
assign micromatr[42][61] = 9'b111111111;
assign micromatr[42][62] = 9'b111111111;
assign micromatr[42][63] = 9'b111111111;
assign micromatr[42][64] = 9'b111111111;
assign micromatr[42][65] = 9'b111111111;
assign micromatr[42][66] = 9'b111111111;
assign micromatr[42][67] = 9'b111111111;
assign micromatr[42][68] = 9'b111111111;
assign micromatr[42][69] = 9'b111111111;
assign micromatr[42][70] = 9'b111111111;
assign micromatr[42][71] = 9'b111111111;
assign micromatr[42][72] = 9'b111111111;
assign micromatr[42][73] = 9'b111111111;
assign micromatr[42][74] = 9'b111111111;
assign micromatr[42][75] = 9'b111111111;
assign micromatr[42][76] = 9'b111111111;
assign micromatr[42][77] = 9'b111111111;
assign micromatr[42][78] = 9'b111111111;
assign micromatr[42][79] = 9'b111111111;
assign micromatr[42][80] = 9'b111111111;
assign micromatr[42][81] = 9'b111111111;
assign micromatr[42][82] = 9'b111111111;
assign micromatr[42][83] = 9'b111111111;
assign micromatr[42][84] = 9'b111111111;
assign micromatr[42][85] = 9'b111111111;
assign micromatr[42][86] = 9'b111111111;
assign micromatr[42][87] = 9'b111111111;
assign micromatr[42][88] = 9'b111111111;
assign micromatr[42][89] = 9'b111111111;
assign micromatr[42][90] = 9'b111111111;
assign micromatr[42][91] = 9'b111111111;
assign micromatr[42][92] = 9'b111111111;
assign micromatr[42][93] = 9'b111111111;
assign micromatr[42][94] = 9'b111111111;
assign micromatr[42][95] = 9'b111111111;
assign micromatr[42][96] = 9'b111111111;
assign micromatr[42][97] = 9'b111111111;
assign micromatr[42][98] = 9'b111111111;
assign micromatr[42][99] = 9'b111111111;
assign micromatr[43][0] = 9'b111111111;
assign micromatr[43][1] = 9'b111111111;
assign micromatr[43][2] = 9'b111111111;
assign micromatr[43][3] = 9'b111111111;
assign micromatr[43][4] = 9'b111111111;
assign micromatr[43][5] = 9'b111111111;
assign micromatr[43][6] = 9'b111111111;
assign micromatr[43][7] = 9'b111111111;
assign micromatr[43][8] = 9'b111111111;
assign micromatr[43][9] = 9'b111111111;
assign micromatr[43][10] = 9'b111111111;
assign micromatr[43][11] = 9'b111111111;
assign micromatr[43][12] = 9'b111111111;
assign micromatr[43][13] = 9'b111111111;
assign micromatr[43][14] = 9'b111111111;
assign micromatr[43][15] = 9'b111111111;
assign micromatr[43][16] = 9'b111111111;
assign micromatr[43][17] = 9'b111111111;
assign micromatr[43][18] = 9'b111111111;
assign micromatr[43][19] = 9'b111111111;
assign micromatr[43][20] = 9'b111111111;
assign micromatr[43][21] = 9'b111111111;
assign micromatr[43][22] = 9'b111111111;
assign micromatr[43][23] = 9'b111111111;
assign micromatr[43][24] = 9'b111111111;
assign micromatr[43][25] = 9'b111111111;
assign micromatr[43][26] = 9'b111111111;
assign micromatr[43][27] = 9'b111111111;
assign micromatr[43][28] = 9'b111111111;
assign micromatr[43][29] = 9'b111111111;
assign micromatr[43][30] = 9'b111111111;
assign micromatr[43][31] = 9'b111111111;
assign micromatr[43][32] = 9'b111111111;
assign micromatr[43][33] = 9'b111111111;
assign micromatr[43][34] = 9'b111111111;
assign micromatr[43][35] = 9'b111111111;
assign micromatr[43][36] = 9'b111111111;
assign micromatr[43][37] = 9'b111111111;
assign micromatr[43][38] = 9'b111111111;
assign micromatr[43][39] = 9'b111111111;
assign micromatr[43][40] = 9'b111111111;
assign micromatr[43][41] = 9'b111111111;
assign micromatr[43][42] = 9'b111111111;
assign micromatr[43][43] = 9'b111111111;
assign micromatr[43][44] = 9'b111111111;
assign micromatr[43][45] = 9'b111111111;
assign micromatr[43][46] = 9'b111111111;
assign micromatr[43][47] = 9'b111111111;
assign micromatr[43][48] = 9'b111111111;
assign micromatr[43][49] = 9'b111111111;
assign micromatr[43][50] = 9'b111111111;
assign micromatr[43][51] = 9'b111111111;
assign micromatr[43][52] = 9'b111111111;
assign micromatr[43][53] = 9'b111111111;
assign micromatr[43][54] = 9'b111111111;
assign micromatr[43][55] = 9'b111111111;
assign micromatr[43][56] = 9'b111111111;
assign micromatr[43][57] = 9'b111111111;
assign micromatr[43][58] = 9'b111111111;
assign micromatr[43][59] = 9'b111111111;
assign micromatr[43][60] = 9'b111111111;
assign micromatr[43][61] = 9'b111111111;
assign micromatr[43][62] = 9'b111111111;
assign micromatr[43][63] = 9'b111111111;
assign micromatr[43][64] = 9'b111111111;
assign micromatr[43][65] = 9'b111111111;
assign micromatr[43][66] = 9'b111111111;
assign micromatr[43][67] = 9'b111111111;
assign micromatr[43][68] = 9'b111111111;
assign micromatr[43][69] = 9'b111111111;
assign micromatr[43][70] = 9'b111111111;
assign micromatr[43][71] = 9'b111111111;
assign micromatr[43][72] = 9'b111111111;
assign micromatr[43][73] = 9'b111111111;
assign micromatr[43][74] = 9'b111111111;
assign micromatr[43][75] = 9'b111111111;
assign micromatr[43][76] = 9'b111111111;
assign micromatr[43][77] = 9'b111111111;
assign micromatr[43][78] = 9'b111111111;
assign micromatr[43][79] = 9'b111111111;
assign micromatr[43][80] = 9'b111111111;
assign micromatr[43][81] = 9'b111111111;
assign micromatr[43][82] = 9'b111111111;
assign micromatr[43][83] = 9'b111111111;
assign micromatr[43][84] = 9'b111111111;
assign micromatr[43][85] = 9'b111111111;
assign micromatr[43][86] = 9'b111111111;
assign micromatr[43][87] = 9'b111111111;
assign micromatr[43][88] = 9'b111111111;
assign micromatr[43][89] = 9'b111111111;
assign micromatr[43][90] = 9'b111111111;
assign micromatr[43][91] = 9'b111111111;
assign micromatr[43][92] = 9'b111111111;
assign micromatr[43][93] = 9'b111111111;
assign micromatr[43][94] = 9'b111111111;
assign micromatr[43][95] = 9'b111111111;
assign micromatr[43][96] = 9'b111111111;
assign micromatr[43][97] = 9'b111111111;
assign micromatr[43][98] = 9'b111111111;
assign micromatr[43][99] = 9'b111111111;
assign micromatr[44][0] = 9'b111111111;
assign micromatr[44][1] = 9'b111111111;
assign micromatr[44][2] = 9'b111111111;
assign micromatr[44][3] = 9'b111111111;
assign micromatr[44][4] = 9'b111111111;
assign micromatr[44][5] = 9'b111111111;
assign micromatr[44][6] = 9'b111111111;
assign micromatr[44][7] = 9'b111111111;
assign micromatr[44][8] = 9'b111111111;
assign micromatr[44][9] = 9'b111111111;
assign micromatr[44][10] = 9'b111111111;
assign micromatr[44][11] = 9'b111111111;
assign micromatr[44][12] = 9'b111111111;
assign micromatr[44][13] = 9'b111111111;
assign micromatr[44][14] = 9'b111111111;
assign micromatr[44][15] = 9'b111111111;
assign micromatr[44][16] = 9'b111111111;
assign micromatr[44][17] = 9'b111111111;
assign micromatr[44][18] = 9'b111111111;
assign micromatr[44][19] = 9'b111111111;
assign micromatr[44][20] = 9'b111111111;
assign micromatr[44][21] = 9'b111111111;
assign micromatr[44][22] = 9'b111111111;
assign micromatr[44][23] = 9'b111111111;
assign micromatr[44][24] = 9'b111111111;
assign micromatr[44][25] = 9'b111111111;
assign micromatr[44][26] = 9'b111111111;
assign micromatr[44][27] = 9'b111111111;
assign micromatr[44][28] = 9'b111111111;
assign micromatr[44][29] = 9'b111111111;
assign micromatr[44][30] = 9'b111111111;
assign micromatr[44][31] = 9'b111111111;
assign micromatr[44][32] = 9'b111111111;
assign micromatr[44][33] = 9'b111111111;
assign micromatr[44][34] = 9'b111111111;
assign micromatr[44][35] = 9'b111111111;
assign micromatr[44][36] = 9'b111111111;
assign micromatr[44][37] = 9'b111111111;
assign micromatr[44][38] = 9'b111111111;
assign micromatr[44][39] = 9'b111111111;
assign micromatr[44][40] = 9'b111111111;
assign micromatr[44][41] = 9'b111111111;
assign micromatr[44][42] = 9'b111111111;
assign micromatr[44][43] = 9'b111111111;
assign micromatr[44][44] = 9'b111111111;
assign micromatr[44][45] = 9'b111111111;
assign micromatr[44][46] = 9'b111111111;
assign micromatr[44][47] = 9'b111111111;
assign micromatr[44][48] = 9'b111111111;
assign micromatr[44][49] = 9'b111111111;
assign micromatr[44][50] = 9'b111111111;
assign micromatr[44][51] = 9'b111111111;
assign micromatr[44][52] = 9'b111111111;
assign micromatr[44][53] = 9'b111111111;
assign micromatr[44][54] = 9'b111111111;
assign micromatr[44][55] = 9'b111111111;
assign micromatr[44][56] = 9'b111111111;
assign micromatr[44][57] = 9'b111111111;
assign micromatr[44][58] = 9'b111111111;
assign micromatr[44][59] = 9'b111111111;
assign micromatr[44][60] = 9'b111111111;
assign micromatr[44][61] = 9'b111111111;
assign micromatr[44][62] = 9'b111111111;
assign micromatr[44][63] = 9'b111111111;
assign micromatr[44][64] = 9'b111111111;
assign micromatr[44][65] = 9'b111111111;
assign micromatr[44][66] = 9'b111111111;
assign micromatr[44][67] = 9'b111111111;
assign micromatr[44][68] = 9'b111111111;
assign micromatr[44][69] = 9'b111111111;
assign micromatr[44][70] = 9'b111111111;
assign micromatr[44][71] = 9'b111111111;
assign micromatr[44][72] = 9'b111111111;
assign micromatr[44][73] = 9'b111111111;
assign micromatr[44][74] = 9'b111111111;
assign micromatr[44][75] = 9'b111111111;
assign micromatr[44][76] = 9'b111111111;
assign micromatr[44][77] = 9'b111111111;
assign micromatr[44][78] = 9'b111111111;
assign micromatr[44][79] = 9'b111111111;
assign micromatr[44][80] = 9'b111111111;
assign micromatr[44][81] = 9'b111111111;
assign micromatr[44][82] = 9'b111111111;
assign micromatr[44][83] = 9'b111111111;
assign micromatr[44][84] = 9'b111111111;
assign micromatr[44][85] = 9'b111111111;
assign micromatr[44][86] = 9'b111111111;
assign micromatr[44][87] = 9'b111111111;
assign micromatr[44][88] = 9'b111111111;
assign micromatr[44][89] = 9'b111111111;
assign micromatr[44][90] = 9'b111111111;
assign micromatr[44][91] = 9'b111111111;
assign micromatr[44][92] = 9'b111111111;
assign micromatr[44][93] = 9'b111111111;
assign micromatr[44][94] = 9'b111111111;
assign micromatr[44][95] = 9'b111111111;
assign micromatr[44][96] = 9'b111111111;
assign micromatr[44][97] = 9'b111111111;
assign micromatr[44][98] = 9'b111111111;
assign micromatr[44][99] = 9'b111111111;
assign micromatr[45][0] = 9'b111111111;
assign micromatr[45][1] = 9'b111111111;
assign micromatr[45][2] = 9'b111111111;
assign micromatr[45][3] = 9'b111111111;
assign micromatr[45][4] = 9'b111111111;
assign micromatr[45][5] = 9'b111111111;
assign micromatr[45][6] = 9'b111111111;
assign micromatr[45][7] = 9'b111111111;
assign micromatr[45][8] = 9'b111111111;
assign micromatr[45][9] = 9'b111111111;
assign micromatr[45][10] = 9'b111111111;
assign micromatr[45][11] = 9'b111111111;
assign micromatr[45][12] = 9'b111111111;
assign micromatr[45][13] = 9'b111111111;
assign micromatr[45][14] = 9'b111111111;
assign micromatr[45][15] = 9'b111111111;
assign micromatr[45][16] = 9'b111111111;
assign micromatr[45][17] = 9'b111111111;
assign micromatr[45][18] = 9'b111111111;
assign micromatr[45][19] = 9'b111111111;
assign micromatr[45][20] = 9'b111111111;
assign micromatr[45][21] = 9'b111111111;
assign micromatr[45][22] = 9'b111111111;
assign micromatr[45][23] = 9'b111111111;
assign micromatr[45][24] = 9'b111111111;
assign micromatr[45][25] = 9'b111111111;
assign micromatr[45][26] = 9'b111111111;
assign micromatr[45][27] = 9'b111111111;
assign micromatr[45][28] = 9'b111111111;
assign micromatr[45][29] = 9'b111111111;
assign micromatr[45][30] = 9'b111111111;
assign micromatr[45][31] = 9'b111111111;
assign micromatr[45][32] = 9'b111111111;
assign micromatr[45][33] = 9'b111111111;
assign micromatr[45][34] = 9'b111111111;
assign micromatr[45][35] = 9'b111111111;
assign micromatr[45][36] = 9'b111111111;
assign micromatr[45][37] = 9'b111111111;
assign micromatr[45][38] = 9'b111111111;
assign micromatr[45][39] = 9'b111111111;
assign micromatr[45][40] = 9'b111111111;
assign micromatr[45][41] = 9'b111111111;
assign micromatr[45][42] = 9'b111111111;
assign micromatr[45][43] = 9'b111111111;
assign micromatr[45][44] = 9'b111111111;
assign micromatr[45][45] = 9'b111111111;
assign micromatr[45][46] = 9'b111111111;
assign micromatr[45][47] = 9'b111111111;
assign micromatr[45][48] = 9'b111111111;
assign micromatr[45][49] = 9'b111111111;
assign micromatr[45][50] = 9'b111111111;
assign micromatr[45][51] = 9'b111111111;
assign micromatr[45][52] = 9'b111111111;
assign micromatr[45][53] = 9'b111111111;
assign micromatr[45][54] = 9'b111111111;
assign micromatr[45][55] = 9'b111111111;
assign micromatr[45][56] = 9'b111111111;
assign micromatr[45][57] = 9'b111111111;
assign micromatr[45][58] = 9'b111111111;
assign micromatr[45][59] = 9'b111111111;
assign micromatr[45][60] = 9'b111111111;
assign micromatr[45][61] = 9'b111111111;
assign micromatr[45][62] = 9'b111111111;
assign micromatr[45][63] = 9'b111111111;
assign micromatr[45][64] = 9'b111111111;
assign micromatr[45][65] = 9'b111111111;
assign micromatr[45][66] = 9'b111111111;
assign micromatr[45][67] = 9'b111111111;
assign micromatr[45][68] = 9'b111111111;
assign micromatr[45][69] = 9'b111111111;
assign micromatr[45][70] = 9'b111111111;
assign micromatr[45][71] = 9'b111111111;
assign micromatr[45][72] = 9'b111111111;
assign micromatr[45][73] = 9'b111111111;
assign micromatr[45][74] = 9'b111111111;
assign micromatr[45][75] = 9'b111111111;
assign micromatr[45][76] = 9'b111111111;
assign micromatr[45][77] = 9'b111111111;
assign micromatr[45][78] = 9'b111111111;
assign micromatr[45][79] = 9'b111111111;
assign micromatr[45][80] = 9'b111111111;
assign micromatr[45][81] = 9'b111111111;
assign micromatr[45][82] = 9'b111111111;
assign micromatr[45][83] = 9'b111111111;
assign micromatr[45][84] = 9'b111111111;
assign micromatr[45][85] = 9'b111111111;
assign micromatr[45][86] = 9'b111111111;
assign micromatr[45][87] = 9'b111111111;
assign micromatr[45][88] = 9'b111111111;
assign micromatr[45][89] = 9'b111111111;
assign micromatr[45][90] = 9'b111111111;
assign micromatr[45][91] = 9'b111111111;
assign micromatr[45][92] = 9'b111111111;
assign micromatr[45][93] = 9'b111111111;
assign micromatr[45][94] = 9'b111111111;
assign micromatr[45][95] = 9'b111111111;
assign micromatr[45][96] = 9'b111111111;
assign micromatr[45][97] = 9'b111111111;
assign micromatr[45][98] = 9'b111111111;
assign micromatr[45][99] = 9'b111111111;
assign micromatr[46][0] = 9'b111111111;
assign micromatr[46][1] = 9'b111111111;
assign micromatr[46][2] = 9'b111111111;
assign micromatr[46][3] = 9'b111111111;
assign micromatr[46][4] = 9'b111111111;
assign micromatr[46][5] = 9'b111111111;
assign micromatr[46][6] = 9'b111111111;
assign micromatr[46][7] = 9'b111111111;
assign micromatr[46][8] = 9'b111111111;
assign micromatr[46][9] = 9'b111111111;
assign micromatr[46][10] = 9'b111111111;
assign micromatr[46][11] = 9'b111111111;
assign micromatr[46][12] = 9'b111111111;
assign micromatr[46][13] = 9'b111111111;
assign micromatr[46][14] = 9'b111111111;
assign micromatr[46][15] = 9'b111111111;
assign micromatr[46][16] = 9'b111111111;
assign micromatr[46][17] = 9'b111111111;
assign micromatr[46][18] = 9'b111111111;
assign micromatr[46][19] = 9'b111111111;
assign micromatr[46][20] = 9'b111111111;
assign micromatr[46][21] = 9'b111111111;
assign micromatr[46][22] = 9'b111111111;
assign micromatr[46][23] = 9'b111111111;
assign micromatr[46][24] = 9'b111111111;
assign micromatr[46][25] = 9'b111111111;
assign micromatr[46][26] = 9'b111111111;
assign micromatr[46][27] = 9'b111111111;
assign micromatr[46][28] = 9'b111111111;
assign micromatr[46][29] = 9'b111111111;
assign micromatr[46][30] = 9'b111111111;
assign micromatr[46][31] = 9'b111111111;
assign micromatr[46][32] = 9'b111111111;
assign micromatr[46][33] = 9'b111111111;
assign micromatr[46][34] = 9'b111111111;
assign micromatr[46][35] = 9'b111111111;
assign micromatr[46][36] = 9'b111111111;
assign micromatr[46][37] = 9'b111111111;
assign micromatr[46][38] = 9'b111111111;
assign micromatr[46][39] = 9'b111111111;
assign micromatr[46][40] = 9'b111111111;
assign micromatr[46][41] = 9'b111111111;
assign micromatr[46][42] = 9'b111111111;
assign micromatr[46][43] = 9'b111111111;
assign micromatr[46][44] = 9'b111111111;
assign micromatr[46][45] = 9'b111111111;
assign micromatr[46][46] = 9'b111111111;
assign micromatr[46][47] = 9'b111111111;
assign micromatr[46][48] = 9'b111111111;
assign micromatr[46][49] = 9'b111111111;
assign micromatr[46][50] = 9'b111111111;
assign micromatr[46][51] = 9'b111111111;
assign micromatr[46][52] = 9'b111111111;
assign micromatr[46][53] = 9'b111111111;
assign micromatr[46][54] = 9'b111111111;
assign micromatr[46][55] = 9'b111111111;
assign micromatr[46][56] = 9'b111111111;
assign micromatr[46][57] = 9'b111111111;
assign micromatr[46][58] = 9'b111111111;
assign micromatr[46][59] = 9'b111111111;
assign micromatr[46][60] = 9'b111111111;
assign micromatr[46][61] = 9'b111111111;
assign micromatr[46][62] = 9'b111111111;
assign micromatr[46][63] = 9'b111111111;
assign micromatr[46][64] = 9'b111111111;
assign micromatr[46][65] = 9'b111111111;
assign micromatr[46][66] = 9'b111111111;
assign micromatr[46][67] = 9'b111111111;
assign micromatr[46][68] = 9'b111111111;
assign micromatr[46][69] = 9'b111111111;
assign micromatr[46][70] = 9'b111111111;
assign micromatr[46][71] = 9'b111111111;
assign micromatr[46][72] = 9'b111111111;
assign micromatr[46][73] = 9'b111111111;
assign micromatr[46][74] = 9'b111111111;
assign micromatr[46][75] = 9'b111111111;
assign micromatr[46][76] = 9'b111111111;
assign micromatr[46][77] = 9'b111111111;
assign micromatr[46][78] = 9'b111111111;
assign micromatr[46][79] = 9'b111111111;
assign micromatr[46][80] = 9'b111111111;
assign micromatr[46][81] = 9'b111111111;
assign micromatr[46][82] = 9'b111111111;
assign micromatr[46][83] = 9'b111111111;
assign micromatr[46][84] = 9'b111111111;
assign micromatr[46][85] = 9'b111111111;
assign micromatr[46][86] = 9'b111111111;
assign micromatr[46][87] = 9'b111111111;
assign micromatr[46][88] = 9'b111111111;
assign micromatr[46][89] = 9'b111111111;
assign micromatr[46][90] = 9'b111111111;
assign micromatr[46][91] = 9'b111111111;
assign micromatr[46][92] = 9'b111111111;
assign micromatr[46][93] = 9'b111111111;
assign micromatr[46][94] = 9'b111111111;
assign micromatr[46][95] = 9'b111111111;
assign micromatr[46][96] = 9'b111111111;
assign micromatr[46][97] = 9'b111111111;
assign micromatr[46][98] = 9'b111111111;
assign micromatr[46][99] = 9'b111111111;
assign micromatr[47][0] = 9'b111111111;
assign micromatr[47][1] = 9'b111111111;
assign micromatr[47][2] = 9'b111111111;
assign micromatr[47][3] = 9'b111111111;
assign micromatr[47][4] = 9'b111111111;
assign micromatr[47][5] = 9'b111111111;
assign micromatr[47][6] = 9'b111111111;
assign micromatr[47][7] = 9'b111111111;
assign micromatr[47][8] = 9'b111111111;
assign micromatr[47][9] = 9'b111111111;
assign micromatr[47][10] = 9'b111111111;
assign micromatr[47][11] = 9'b111111111;
assign micromatr[47][12] = 9'b111111111;
assign micromatr[47][13] = 9'b111111111;
assign micromatr[47][14] = 9'b111111111;
assign micromatr[47][15] = 9'b111111111;
assign micromatr[47][16] = 9'b111111111;
assign micromatr[47][17] = 9'b111111111;
assign micromatr[47][18] = 9'b111111111;
assign micromatr[47][19] = 9'b111111111;
assign micromatr[47][20] = 9'b111111111;
assign micromatr[47][21] = 9'b111111111;
assign micromatr[47][22] = 9'b111111111;
assign micromatr[47][23] = 9'b111111111;
assign micromatr[47][24] = 9'b111111111;
assign micromatr[47][25] = 9'b111111111;
assign micromatr[47][26] = 9'b111111111;
assign micromatr[47][27] = 9'b111111111;
assign micromatr[47][28] = 9'b111111111;
assign micromatr[47][29] = 9'b111111111;
assign micromatr[47][30] = 9'b111111111;
assign micromatr[47][31] = 9'b111111111;
assign micromatr[47][32] = 9'b111111111;
assign micromatr[47][33] = 9'b111111111;
assign micromatr[47][34] = 9'b111111111;
assign micromatr[47][35] = 9'b111111111;
assign micromatr[47][36] = 9'b111111111;
assign micromatr[47][37] = 9'b111111111;
assign micromatr[47][38] = 9'b111111111;
assign micromatr[47][39] = 9'b111111111;
assign micromatr[47][40] = 9'b111111111;
assign micromatr[47][41] = 9'b111111111;
assign micromatr[47][42] = 9'b111111111;
assign micromatr[47][43] = 9'b111111111;
assign micromatr[47][44] = 9'b111111111;
assign micromatr[47][45] = 9'b111111111;
assign micromatr[47][46] = 9'b111111111;
assign micromatr[47][47] = 9'b111111111;
assign micromatr[47][48] = 9'b111111111;
assign micromatr[47][49] = 9'b111111111;
assign micromatr[47][50] = 9'b111111111;
assign micromatr[47][51] = 9'b111111111;
assign micromatr[47][52] = 9'b111111111;
assign micromatr[47][53] = 9'b111111111;
assign micromatr[47][54] = 9'b111111111;
assign micromatr[47][55] = 9'b111111111;
assign micromatr[47][56] = 9'b111111111;
assign micromatr[47][57] = 9'b111111111;
assign micromatr[47][58] = 9'b111111111;
assign micromatr[47][59] = 9'b111111111;
assign micromatr[47][60] = 9'b111111111;
assign micromatr[47][61] = 9'b111111111;
assign micromatr[47][62] = 9'b111111111;
assign micromatr[47][63] = 9'b111111111;
assign micromatr[47][64] = 9'b111111111;
assign micromatr[47][65] = 9'b111111111;
assign micromatr[47][66] = 9'b111111111;
assign micromatr[47][67] = 9'b111111111;
assign micromatr[47][68] = 9'b111111111;
assign micromatr[47][69] = 9'b111111111;
assign micromatr[47][70] = 9'b111111111;
assign micromatr[47][71] = 9'b111111111;
assign micromatr[47][72] = 9'b111111111;
assign micromatr[47][73] = 9'b111111111;
assign micromatr[47][74] = 9'b111111111;
assign micromatr[47][75] = 9'b111111111;
assign micromatr[47][76] = 9'b111111111;
assign micromatr[47][77] = 9'b111111111;
assign micromatr[47][78] = 9'b111111111;
assign micromatr[47][79] = 9'b111111111;
assign micromatr[47][80] = 9'b111111111;
assign micromatr[47][81] = 9'b111111111;
assign micromatr[47][82] = 9'b111111111;
assign micromatr[47][83] = 9'b111111111;
assign micromatr[47][84] = 9'b111111111;
assign micromatr[47][85] = 9'b111111111;
assign micromatr[47][86] = 9'b111111111;
assign micromatr[47][87] = 9'b111111111;
assign micromatr[47][88] = 9'b111111111;
assign micromatr[47][89] = 9'b111111111;
assign micromatr[47][90] = 9'b111111111;
assign micromatr[47][91] = 9'b111111111;
assign micromatr[47][92] = 9'b111111111;
assign micromatr[47][93] = 9'b111111111;
assign micromatr[47][94] = 9'b111111111;
assign micromatr[47][95] = 9'b111111111;
assign micromatr[47][96] = 9'b111111111;
assign micromatr[47][97] = 9'b111111111;
assign micromatr[47][98] = 9'b111111111;
assign micromatr[47][99] = 9'b111111111;
assign micromatr[48][0] = 9'b111111111;
assign micromatr[48][1] = 9'b111111111;
assign micromatr[48][2] = 9'b111111111;
assign micromatr[48][3] = 9'b111111111;
assign micromatr[48][4] = 9'b111111111;
assign micromatr[48][5] = 9'b111111111;
assign micromatr[48][6] = 9'b111111111;
assign micromatr[48][7] = 9'b111111111;
assign micromatr[48][8] = 9'b111111111;
assign micromatr[48][9] = 9'b111111111;
assign micromatr[48][10] = 9'b111111111;
assign micromatr[48][11] = 9'b111111111;
assign micromatr[48][12] = 9'b111111111;
assign micromatr[48][13] = 9'b111111111;
assign micromatr[48][14] = 9'b111111111;
assign micromatr[48][15] = 9'b111111111;
assign micromatr[48][16] = 9'b111111111;
assign micromatr[48][17] = 9'b111111111;
assign micromatr[48][18] = 9'b111111111;
assign micromatr[48][19] = 9'b111111111;
assign micromatr[48][20] = 9'b111111111;
assign micromatr[48][21] = 9'b111111111;
assign micromatr[48][22] = 9'b111111111;
assign micromatr[48][23] = 9'b111111111;
assign micromatr[48][24] = 9'b111111111;
assign micromatr[48][25] = 9'b111111111;
assign micromatr[48][26] = 9'b111111111;
assign micromatr[48][27] = 9'b111111111;
assign micromatr[48][28] = 9'b111111111;
assign micromatr[48][29] = 9'b111111111;
assign micromatr[48][30] = 9'b111111111;
assign micromatr[48][31] = 9'b111111111;
assign micromatr[48][32] = 9'b111111111;
assign micromatr[48][33] = 9'b111111111;
assign micromatr[48][34] = 9'b111111111;
assign micromatr[48][35] = 9'b111111111;
assign micromatr[48][36] = 9'b111111111;
assign micromatr[48][37] = 9'b111111111;
assign micromatr[48][38] = 9'b111111111;
assign micromatr[48][39] = 9'b111111111;
assign micromatr[48][40] = 9'b111111111;
assign micromatr[48][41] = 9'b111111111;
assign micromatr[48][42] = 9'b111111111;
assign micromatr[48][43] = 9'b111111111;
assign micromatr[48][44] = 9'b111111111;
assign micromatr[48][45] = 9'b111111111;
assign micromatr[48][46] = 9'b111111111;
assign micromatr[48][47] = 9'b111111111;
assign micromatr[48][48] = 9'b111111111;
assign micromatr[48][49] = 9'b111111111;
assign micromatr[48][50] = 9'b111111111;
assign micromatr[48][51] = 9'b111111111;
assign micromatr[48][52] = 9'b111111111;
assign micromatr[48][53] = 9'b111111111;
assign micromatr[48][54] = 9'b111111111;
assign micromatr[48][55] = 9'b111111111;
assign micromatr[48][56] = 9'b111111111;
assign micromatr[48][57] = 9'b111111111;
assign micromatr[48][58] = 9'b111111111;
assign micromatr[48][59] = 9'b111111111;
assign micromatr[48][60] = 9'b111111111;
assign micromatr[48][61] = 9'b111111111;
assign micromatr[48][62] = 9'b111111111;
assign micromatr[48][63] = 9'b111111111;
assign micromatr[48][64] = 9'b111111111;
assign micromatr[48][65] = 9'b111111111;
assign micromatr[48][66] = 9'b111111111;
assign micromatr[48][67] = 9'b111111111;
assign micromatr[48][68] = 9'b111111111;
assign micromatr[48][69] = 9'b111111111;
assign micromatr[48][70] = 9'b111111111;
assign micromatr[48][71] = 9'b111111111;
assign micromatr[48][72] = 9'b111111111;
assign micromatr[48][73] = 9'b111111111;
assign micromatr[48][74] = 9'b111111111;
assign micromatr[48][75] = 9'b111111111;
assign micromatr[48][76] = 9'b111111111;
assign micromatr[48][77] = 9'b111111111;
assign micromatr[48][78] = 9'b111111111;
assign micromatr[48][79] = 9'b111111111;
assign micromatr[48][80] = 9'b111111111;
assign micromatr[48][81] = 9'b111111111;
assign micromatr[48][82] = 9'b111111111;
assign micromatr[48][83] = 9'b111111111;
assign micromatr[48][84] = 9'b111111111;
assign micromatr[48][85] = 9'b111111111;
assign micromatr[48][86] = 9'b111111111;
assign micromatr[48][87] = 9'b111111111;
assign micromatr[48][88] = 9'b111111111;
assign micromatr[48][89] = 9'b111111111;
assign micromatr[48][90] = 9'b111111111;
assign micromatr[48][91] = 9'b111111111;
assign micromatr[48][92] = 9'b111111111;
assign micromatr[48][93] = 9'b111111111;
assign micromatr[48][94] = 9'b111111111;
assign micromatr[48][95] = 9'b111111111;
assign micromatr[48][96] = 9'b111111111;
assign micromatr[48][97] = 9'b111111111;
assign micromatr[48][98] = 9'b111111111;
assign micromatr[48][99] = 9'b111111111;
assign micromatr[49][0] = 9'b111111111;
assign micromatr[49][1] = 9'b111111111;
assign micromatr[49][2] = 9'b111111111;
assign micromatr[49][3] = 9'b111111111;
assign micromatr[49][4] = 9'b111111111;
assign micromatr[49][5] = 9'b111111111;
assign micromatr[49][6] = 9'b111111111;
assign micromatr[49][7] = 9'b111111111;
assign micromatr[49][8] = 9'b111111111;
assign micromatr[49][9] = 9'b111111111;
assign micromatr[49][10] = 9'b111111111;
assign micromatr[49][11] = 9'b111111111;
assign micromatr[49][12] = 9'b111111111;
assign micromatr[49][13] = 9'b111111111;
assign micromatr[49][14] = 9'b111111111;
assign micromatr[49][15] = 9'b111111111;
assign micromatr[49][16] = 9'b111111111;
assign micromatr[49][17] = 9'b111111111;
assign micromatr[49][18] = 9'b111111111;
assign micromatr[49][19] = 9'b111111111;
assign micromatr[49][20] = 9'b111111111;
assign micromatr[49][21] = 9'b111111111;
assign micromatr[49][22] = 9'b111111111;
assign micromatr[49][23] = 9'b111111111;
assign micromatr[49][24] = 9'b111111111;
assign micromatr[49][25] = 9'b111111111;
assign micromatr[49][26] = 9'b111111111;
assign micromatr[49][27] = 9'b111111111;
assign micromatr[49][28] = 9'b111111111;
assign micromatr[49][29] = 9'b111111111;
assign micromatr[49][30] = 9'b111111111;
assign micromatr[49][31] = 9'b111111111;
assign micromatr[49][32] = 9'b111111111;
assign micromatr[49][33] = 9'b111111111;
assign micromatr[49][34] = 9'b111111111;
assign micromatr[49][35] = 9'b111111111;
assign micromatr[49][36] = 9'b111111111;
assign micromatr[49][37] = 9'b111111111;
assign micromatr[49][38] = 9'b111111111;
assign micromatr[49][39] = 9'b111111111;
assign micromatr[49][40] = 9'b111111111;
assign micromatr[49][41] = 9'b111111111;
assign micromatr[49][42] = 9'b111111111;
assign micromatr[49][43] = 9'b111111111;
assign micromatr[49][44] = 9'b111111111;
assign micromatr[49][45] = 9'b111111111;
assign micromatr[49][46] = 9'b111111111;
assign micromatr[49][47] = 9'b111111111;
assign micromatr[49][48] = 9'b111111111;
assign micromatr[49][49] = 9'b111111111;
assign micromatr[49][50] = 9'b111111111;
assign micromatr[49][51] = 9'b111111111;
assign micromatr[49][52] = 9'b111111111;
assign micromatr[49][53] = 9'b111111111;
assign micromatr[49][54] = 9'b111111111;
assign micromatr[49][55] = 9'b111111111;
assign micromatr[49][56] = 9'b111111111;
assign micromatr[49][57] = 9'b111111111;
assign micromatr[49][58] = 9'b111111111;
assign micromatr[49][59] = 9'b111111111;
assign micromatr[49][60] = 9'b111111111;
assign micromatr[49][61] = 9'b111111111;
assign micromatr[49][62] = 9'b111111111;
assign micromatr[49][63] = 9'b111111111;
assign micromatr[49][64] = 9'b111111111;
assign micromatr[49][65] = 9'b111111111;
assign micromatr[49][66] = 9'b111111111;
assign micromatr[49][67] = 9'b111111111;
assign micromatr[49][68] = 9'b111111111;
assign micromatr[49][69] = 9'b111111111;
assign micromatr[49][70] = 9'b111111111;
assign micromatr[49][71] = 9'b111111111;
assign micromatr[49][72] = 9'b111111111;
assign micromatr[49][73] = 9'b111111111;
assign micromatr[49][74] = 9'b111111111;
assign micromatr[49][75] = 9'b111111111;
assign micromatr[49][76] = 9'b111111111;
assign micromatr[49][77] = 9'b111111111;
assign micromatr[49][78] = 9'b111111111;
assign micromatr[49][79] = 9'b111111111;
assign micromatr[49][80] = 9'b111111111;
assign micromatr[49][81] = 9'b111111111;
assign micromatr[49][82] = 9'b111111111;
assign micromatr[49][83] = 9'b111111111;
assign micromatr[49][84] = 9'b111111111;
assign micromatr[49][85] = 9'b111111111;
assign micromatr[49][86] = 9'b111111111;
assign micromatr[49][87] = 9'b111111111;
assign micromatr[49][88] = 9'b111111111;
assign micromatr[49][89] = 9'b111111111;
assign micromatr[49][90] = 9'b111111111;
assign micromatr[49][91] = 9'b111111111;
assign micromatr[49][92] = 9'b111111111;
assign micromatr[49][93] = 9'b111111111;
assign micromatr[49][94] = 9'b111111111;
assign micromatr[49][95] = 9'b111111111;
assign micromatr[49][96] = 9'b111111111;
assign micromatr[49][97] = 9'b111111111;
assign micromatr[49][98] = 9'b111111111;
assign micromatr[49][99] = 9'b111111111;
//Total de Lineas = 5000
endmodule

