`timescale 1ns / 1ps
module cpo (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (f[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= f[vcount- posy][hcount- posx][7:5];
				green <= f[vcount- posy][hcount- posx][4:2];
            blue 	<= f[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 100;
parameter RESOLUCION_Y = 50;
wire [8:0] f[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign f[2][58] = 9'b100000000;
assign f[2][59] = 9'b100000000;
assign f[2][60] = 9'b100000000;
assign f[2][61] = 9'b100000000;
assign f[2][62] = 9'b100000000;
assign f[2][63] = 9'b100000000;
assign f[2][64] = 9'b100000000;
assign f[2][65] = 9'b100000000;
assign f[2][66] = 9'b100000000;
assign f[2][67] = 9'b100000000;
assign f[2][68] = 9'b100000000;
assign f[2][69] = 9'b100000000;
assign f[2][70] = 9'b100000000;
assign f[2][71] = 9'b100000000;
assign f[2][72] = 9'b100000000;
assign f[2][73] = 9'b100000000;
assign f[2][74] = 9'b100000000;
assign f[2][75] = 9'b100000000;
assign f[2][76] = 9'b100000000;
assign f[2][77] = 9'b100000000;
assign f[2][78] = 9'b100000000;
assign f[2][79] = 9'b100000000;
assign f[2][80] = 9'b100000000;
assign f[2][81] = 9'b100000000;
assign f[2][82] = 9'b100000000;
assign f[2][83] = 9'b100000000;
assign f[2][84] = 9'b100000000;
assign f[2][85] = 9'b100000000;
assign f[2][86] = 9'b100000000;
assign f[2][87] = 9'b100000000;
assign f[2][88] = 9'b100000000;
assign f[3][57] = 9'b100000000;
assign f[3][58] = 9'b101001001;
assign f[3][59] = 9'b101101101;
assign f[3][60] = 9'b110010001;
assign f[3][61] = 9'b110001101;
assign f[3][62] = 9'b110001101;
assign f[3][63] = 9'b110010001;
assign f[3][64] = 9'b110001101;
assign f[3][65] = 9'b101101101;
assign f[3][66] = 9'b110010001;
assign f[3][67] = 9'b110010001;
assign f[3][68] = 9'b110010001;
assign f[3][69] = 9'b110010001;
assign f[3][70] = 9'b110010001;
assign f[3][71] = 9'b110010001;
assign f[3][72] = 9'b110010001;
assign f[3][73] = 9'b110010001;
assign f[3][74] = 9'b110010001;
assign f[3][75] = 9'b110010001;
assign f[3][76] = 9'b110010001;
assign f[3][77] = 9'b110010001;
assign f[3][78] = 9'b110010001;
assign f[3][79] = 9'b110010001;
assign f[3][80] = 9'b110010001;
assign f[3][81] = 9'b110010001;
assign f[3][82] = 9'b110010001;
assign f[3][83] = 9'b110010001;
assign f[3][84] = 9'b110010001;
assign f[3][85] = 9'b110010001;
assign f[3][86] = 9'b110010001;
assign f[3][87] = 9'b110010001;
assign f[3][88] = 9'b101101101;
assign f[3][89] = 9'b100100100;
assign f[3][90] = 9'b100000000;
assign f[4][56] = 9'b100000000;
assign f[4][57] = 9'b110010001;
assign f[4][58] = 9'b111111111;
assign f[4][59] = 9'b111111111;
assign f[4][60] = 9'b111111111;
assign f[4][61] = 9'b111111111;
assign f[4][62] = 9'b111111111;
assign f[4][63] = 9'b111111111;
assign f[4][64] = 9'b111111111;
assign f[4][65] = 9'b111111111;
assign f[4][66] = 9'b111111111;
assign f[4][67] = 9'b111111111;
assign f[4][68] = 9'b111111111;
assign f[4][69] = 9'b111111111;
assign f[4][70] = 9'b111111111;
assign f[4][71] = 9'b111111111;
assign f[4][72] = 9'b111111111;
assign f[4][73] = 9'b111111111;
assign f[4][74] = 9'b111111111;
assign f[4][75] = 9'b111111111;
assign f[4][76] = 9'b111111111;
assign f[4][77] = 9'b111111111;
assign f[4][78] = 9'b111111111;
assign f[4][79] = 9'b111111111;
assign f[4][80] = 9'b111111111;
assign f[4][81] = 9'b111111111;
assign f[4][82] = 9'b111111111;
assign f[4][83] = 9'b111111111;
assign f[4][84] = 9'b111111111;
assign f[4][85] = 9'b111111111;
assign f[4][86] = 9'b111111111;
assign f[4][87] = 9'b111111111;
assign f[4][88] = 9'b111111111;
assign f[4][89] = 9'b111111111;
assign f[4][90] = 9'b100100100;
assign f[5][56] = 9'b100000000;
assign f[5][57] = 9'b110110110;
assign f[5][58] = 9'b111111111;
assign f[5][59] = 9'b111111111;
assign f[5][60] = 9'b111111111;
assign f[5][61] = 9'b111111111;
assign f[5][62] = 9'b111111111;
assign f[5][63] = 9'b111111111;
assign f[5][64] = 9'b111111111;
assign f[5][65] = 9'b111111111;
assign f[5][66] = 9'b111111111;
assign f[5][67] = 9'b111111111;
assign f[5][68] = 9'b111111111;
assign f[5][69] = 9'b111111111;
assign f[5][70] = 9'b111111111;
assign f[5][71] = 9'b111111111;
assign f[5][72] = 9'b111111111;
assign f[5][73] = 9'b111111111;
assign f[5][74] = 9'b111111111;
assign f[5][75] = 9'b111111111;
assign f[5][76] = 9'b111111111;
assign f[5][77] = 9'b111111111;
assign f[5][78] = 9'b111111111;
assign f[5][79] = 9'b111111111;
assign f[5][80] = 9'b111111111;
assign f[5][81] = 9'b111111111;
assign f[5][82] = 9'b111111111;
assign f[5][83] = 9'b111111111;
assign f[5][84] = 9'b111111111;
assign f[5][85] = 9'b111111111;
assign f[5][86] = 9'b111111111;
assign f[5][87] = 9'b111111111;
assign f[5][88] = 9'b111111111;
assign f[5][89] = 9'b111111111;
assign f[5][90] = 9'b101001001;
assign f[6][56] = 9'b100000000;
assign f[6][57] = 9'b110110110;
assign f[6][58] = 9'b111111111;
assign f[6][59] = 9'b111111111;
assign f[6][60] = 9'b111111111;
assign f[6][61] = 9'b111111111;
assign f[6][62] = 9'b111111111;
assign f[6][63] = 9'b111111111;
assign f[6][64] = 9'b111111111;
assign f[6][65] = 9'b111111111;
assign f[6][66] = 9'b111111111;
assign f[6][67] = 9'b111111111;
assign f[6][68] = 9'b111111111;
assign f[6][69] = 9'b111111111;
assign f[6][70] = 9'b111111111;
assign f[6][71] = 9'b111111111;
assign f[6][72] = 9'b111111111;
assign f[6][73] = 9'b111111111;
assign f[6][74] = 9'b111111111;
assign f[6][75] = 9'b111111111;
assign f[6][76] = 9'b111111111;
assign f[6][77] = 9'b111111111;
assign f[6][78] = 9'b111111111;
assign f[6][79] = 9'b111111111;
assign f[6][80] = 9'b111111111;
assign f[6][81] = 9'b111111111;
assign f[6][82] = 9'b111111111;
assign f[6][83] = 9'b111111111;
assign f[6][84] = 9'b111111111;
assign f[6][85] = 9'b111111111;
assign f[6][86] = 9'b111111111;
assign f[6][87] = 9'b111111111;
assign f[6][88] = 9'b111111111;
assign f[6][89] = 9'b111111111;
assign f[6][90] = 9'b101001001;
assign f[7][56] = 9'b100000000;
assign f[7][57] = 9'b110110110;
assign f[7][58] = 9'b111111111;
assign f[7][59] = 9'b111111111;
assign f[7][60] = 9'b111111111;
assign f[7][61] = 9'b101101101;
assign f[7][62] = 9'b101101101;
assign f[7][63] = 9'b111111111;
assign f[7][64] = 9'b111111111;
assign f[7][65] = 9'b110010001;
assign f[7][66] = 9'b111111111;
assign f[7][67] = 9'b111111111;
assign f[7][68] = 9'b111111111;
assign f[7][69] = 9'b111111111;
assign f[7][70] = 9'b111111111;
assign f[7][71] = 9'b111111111;
assign f[7][72] = 9'b101101101;
assign f[7][73] = 9'b101101101;
assign f[7][74] = 9'b111111111;
assign f[7][75] = 9'b111111111;
assign f[7][76] = 9'b110010010;
assign f[7][77] = 9'b111111111;
assign f[7][78] = 9'b111111111;
assign f[7][79] = 9'b111111111;
assign f[7][80] = 9'b111111111;
assign f[7][81] = 9'b111111111;
assign f[7][82] = 9'b111111111;
assign f[7][83] = 9'b111111111;
assign f[7][84] = 9'b111111111;
assign f[7][85] = 9'b111111111;
assign f[7][86] = 9'b111111111;
assign f[7][87] = 9'b111111111;
assign f[7][88] = 9'b111111111;
assign f[7][89] = 9'b111111111;
assign f[7][90] = 9'b101001001;
assign f[8][42] = 9'b100111101;
assign f[8][43] = 9'b100111101;
assign f[8][44] = 9'b100111101;
assign f[8][45] = 9'b100111101;
assign f[8][46] = 9'b100111101;
assign f[8][47] = 9'b100111101;
assign f[8][48] = 9'b100111101;
assign f[8][49] = 9'b100111101;
assign f[8][50] = 9'b100111101;
assign f[8][56] = 9'b100000000;
assign f[8][57] = 9'b110110110;
assign f[8][58] = 9'b111111111;
assign f[8][59] = 9'b111111111;
assign f[8][60] = 9'b111111111;
assign f[8][61] = 9'b101101101;
assign f[8][62] = 9'b110010010;
assign f[8][63] = 9'b111111111;
assign f[8][64] = 9'b111111111;
assign f[8][65] = 9'b110010001;
assign f[8][66] = 9'b111111111;
assign f[8][67] = 9'b111111111;
assign f[8][68] = 9'b111111111;
assign f[8][69] = 9'b111111111;
assign f[8][70] = 9'b111111111;
assign f[8][71] = 9'b111111111;
assign f[8][72] = 9'b101101101;
assign f[8][73] = 9'b110010001;
assign f[8][74] = 9'b110010001;
assign f[8][75] = 9'b111111111;
assign f[8][76] = 9'b110010001;
assign f[8][77] = 9'b111111111;
assign f[8][78] = 9'b111111111;
assign f[8][79] = 9'b111111111;
assign f[8][80] = 9'b110010001;
assign f[8][81] = 9'b110010001;
assign f[8][82] = 9'b111111111;
assign f[8][83] = 9'b110010010;
assign f[8][84] = 9'b101001001;
assign f[8][85] = 9'b111111111;
assign f[8][86] = 9'b111111111;
assign f[8][87] = 9'b111111111;
assign f[8][88] = 9'b111111111;
assign f[8][89] = 9'b111111111;
assign f[8][90] = 9'b101001001;
assign f[9][39] = 9'b100110101;
assign f[9][40] = 9'b100111101;
assign f[9][41] = 9'b100111101;
assign f[9][42] = 9'b100111101;
assign f[9][43] = 9'b100111101;
assign f[9][44] = 9'b100111101;
assign f[9][45] = 9'b100111101;
assign f[9][46] = 9'b100111101;
assign f[9][47] = 9'b100111101;
assign f[9][48] = 9'b100111101;
assign f[9][49] = 9'b100111101;
assign f[9][50] = 9'b100111101;
assign f[9][51] = 9'b100011101;
assign f[9][52] = 9'b100111101;
assign f[9][53] = 9'b100110101;
assign f[9][56] = 9'b100000000;
assign f[9][57] = 9'b110110110;
assign f[9][58] = 9'b111111111;
assign f[9][59] = 9'b111111111;
assign f[9][60] = 9'b111111111;
assign f[9][61] = 9'b101101101;
assign f[9][62] = 9'b111111111;
assign f[9][63] = 9'b111111111;
assign f[9][64] = 9'b111111111;
assign f[9][65] = 9'b110010001;
assign f[9][66] = 9'b111111111;
assign f[9][67] = 9'b111111111;
assign f[9][68] = 9'b111111111;
assign f[9][69] = 9'b111111111;
assign f[9][70] = 9'b111111111;
assign f[9][71] = 9'b111111111;
assign f[9][72] = 9'b101001001;
assign f[9][73] = 9'b110010001;
assign f[9][74] = 9'b111111111;
assign f[9][75] = 9'b111111111;
assign f[9][76] = 9'b110010001;
assign f[9][77] = 9'b111111111;
assign f[9][78] = 9'b111111111;
assign f[9][79] = 9'b111111111;
assign f[9][80] = 9'b101101101;
assign f[9][81] = 9'b101001001;
assign f[9][82] = 9'b111111111;
assign f[9][83] = 9'b110010001;
assign f[9][84] = 9'b101101101;
assign f[9][85] = 9'b110010001;
assign f[9][86] = 9'b111111111;
assign f[9][87] = 9'b111111111;
assign f[9][88] = 9'b111111111;
assign f[9][89] = 9'b111111111;
assign f[9][90] = 9'b101001001;
assign f[10][39] = 9'b100111101;
assign f[10][40] = 9'b100111101;
assign f[10][41] = 9'b100111101;
assign f[10][42] = 9'b100111101;
assign f[10][43] = 9'b100111101;
assign f[10][44] = 9'b100111101;
assign f[10][45] = 9'b100111101;
assign f[10][46] = 9'b100111101;
assign f[10][47] = 9'b100111101;
assign f[10][48] = 9'b100111101;
assign f[10][49] = 9'b100111101;
assign f[10][50] = 9'b100111101;
assign f[10][51] = 9'b100111101;
assign f[10][52] = 9'b100111101;
assign f[10][53] = 9'b100111101;
assign f[10][56] = 9'b100000000;
assign f[10][57] = 9'b110110110;
assign f[10][58] = 9'b111111111;
assign f[10][59] = 9'b111111111;
assign f[10][60] = 9'b111111111;
assign f[10][61] = 9'b101101101;
assign f[10][62] = 9'b110010001;
assign f[10][63] = 9'b111111111;
assign f[10][64] = 9'b111111111;
assign f[10][65] = 9'b110010001;
assign f[10][66] = 9'b110110110;
assign f[10][67] = 9'b111111111;
assign f[10][68] = 9'b111111111;
assign f[10][69] = 9'b111111111;
assign f[10][70] = 9'b111111111;
assign f[10][71] = 9'b111111111;
assign f[10][72] = 9'b101101101;
assign f[10][73] = 9'b111111111;
assign f[10][74] = 9'b111111111;
assign f[10][75] = 9'b111111111;
assign f[10][76] = 9'b110010001;
assign f[10][77] = 9'b110110110;
assign f[10][78] = 9'b111111111;
assign f[10][79] = 9'b111111111;
assign f[10][80] = 9'b100100100;
assign f[10][81] = 9'b101101101;
assign f[10][82] = 9'b111111111;
assign f[10][83] = 9'b110010001;
assign f[10][84] = 9'b110010001;
assign f[10][85] = 9'b110010001;
assign f[10][86] = 9'b111111111;
assign f[10][87] = 9'b111111111;
assign f[10][88] = 9'b111111111;
assign f[10][89] = 9'b111111111;
assign f[10][90] = 9'b101001001;
assign f[11][38] = 9'b100111101;
assign f[11][39] = 9'b100111101;
assign f[11][40] = 9'b100111101;
assign f[11][41] = 9'b100111101;
assign f[11][42] = 9'b100111101;
assign f[11][43] = 9'b100111101;
assign f[11][44] = 9'b100111101;
assign f[11][45] = 9'b100111101;
assign f[11][46] = 9'b100111101;
assign f[11][47] = 9'b110111111;
assign f[11][48] = 9'b111111111;
assign f[11][49] = 9'b111111111;
assign f[11][50] = 9'b111111111;
assign f[11][51] = 9'b111111111;
assign f[11][52] = 9'b101011101;
assign f[11][53] = 9'b100111101;
assign f[11][54] = 9'b100111101;
assign f[11][56] = 9'b100000000;
assign f[11][57] = 9'b110110110;
assign f[11][58] = 9'b111111111;
assign f[11][59] = 9'b111111111;
assign f[11][60] = 9'b111111111;
assign f[11][61] = 9'b111111111;
assign f[11][62] = 9'b110110110;
assign f[11][63] = 9'b111111111;
assign f[11][64] = 9'b111111111;
assign f[11][65] = 9'b111111111;
assign f[11][66] = 9'b111111111;
assign f[11][67] = 9'b111111111;
assign f[11][68] = 9'b111111111;
assign f[11][69] = 9'b111111111;
assign f[11][70] = 9'b111111111;
assign f[11][71] = 9'b111111111;
assign f[11][72] = 9'b111111111;
assign f[11][73] = 9'b111111111;
assign f[11][74] = 9'b111111111;
assign f[11][75] = 9'b111111111;
assign f[11][76] = 9'b111111111;
assign f[11][77] = 9'b111111111;
assign f[11][78] = 9'b111111111;
assign f[11][79] = 9'b111111111;
assign f[11][80] = 9'b111111111;
assign f[11][81] = 9'b111111111;
assign f[11][82] = 9'b111111111;
assign f[11][83] = 9'b111111111;
assign f[11][84] = 9'b111111111;
assign f[11][85] = 9'b111111111;
assign f[11][86] = 9'b111111111;
assign f[11][87] = 9'b111111111;
assign f[11][88] = 9'b111111111;
assign f[11][89] = 9'b111111111;
assign f[11][90] = 9'b101001001;
assign f[12][37] = 9'b100111101;
assign f[12][38] = 9'b100111101;
assign f[12][39] = 9'b100111101;
assign f[12][40] = 9'b100111101;
assign f[12][41] = 9'b100111101;
assign f[12][42] = 9'b100111101;
assign f[12][43] = 9'b100111101;
assign f[12][44] = 9'b100111101;
assign f[12][45] = 9'b100111101;
assign f[12][46] = 9'b100111101;
assign f[12][47] = 9'b111111111;
assign f[12][48] = 9'b111111111;
assign f[12][49] = 9'b111111111;
assign f[12][50] = 9'b111111111;
assign f[12][51] = 9'b111111111;
assign f[12][52] = 9'b101011101;
assign f[12][53] = 9'b100111101;
assign f[12][54] = 9'b100111101;
assign f[12][55] = 9'b100111101;
assign f[12][56] = 9'b100000100;
assign f[12][57] = 9'b110110010;
assign f[12][58] = 9'b111111111;
assign f[12][59] = 9'b111111111;
assign f[12][60] = 9'b111111111;
assign f[12][61] = 9'b111111111;
assign f[12][62] = 9'b111111111;
assign f[12][63] = 9'b111111111;
assign f[12][64] = 9'b111111111;
assign f[12][65] = 9'b111111111;
assign f[12][66] = 9'b111111111;
assign f[12][67] = 9'b111111111;
assign f[12][68] = 9'b111111111;
assign f[12][69] = 9'b111111111;
assign f[12][70] = 9'b111111111;
assign f[12][71] = 9'b111111111;
assign f[12][72] = 9'b111111111;
assign f[12][73] = 9'b111111111;
assign f[12][74] = 9'b111111111;
assign f[12][75] = 9'b111111111;
assign f[12][76] = 9'b111111111;
assign f[12][77] = 9'b111111111;
assign f[12][78] = 9'b111111111;
assign f[12][79] = 9'b111111111;
assign f[12][80] = 9'b111111111;
assign f[12][81] = 9'b111111111;
assign f[12][82] = 9'b111111111;
assign f[12][83] = 9'b111111111;
assign f[12][84] = 9'b111111111;
assign f[12][85] = 9'b111111111;
assign f[12][86] = 9'b111111111;
assign f[12][87] = 9'b111111111;
assign f[12][88] = 9'b111111111;
assign f[12][89] = 9'b111111111;
assign f[12][90] = 9'b101001001;
assign f[13][36] = 9'b100110101;
assign f[13][37] = 9'b100111101;
assign f[13][38] = 9'b100111101;
assign f[13][39] = 9'b100111101;
assign f[13][40] = 9'b100111101;
assign f[13][41] = 9'b100111101;
assign f[13][42] = 9'b100111101;
assign f[13][43] = 9'b100111101;
assign f[13][44] = 9'b100111101;
assign f[13][45] = 9'b100111101;
assign f[13][46] = 9'b100111101;
assign f[13][47] = 9'b110011111;
assign f[13][48] = 9'b111111111;
assign f[13][49] = 9'b111111111;
assign f[13][50] = 9'b111111111;
assign f[13][51] = 9'b111111111;
assign f[13][52] = 9'b101011101;
assign f[13][53] = 9'b100111101;
assign f[13][54] = 9'b100111101;
assign f[13][55] = 9'b100111101;
assign f[13][56] = 9'b100000100;
assign f[13][57] = 9'b110010001;
assign f[13][58] = 9'b111111111;
assign f[13][59] = 9'b111111111;
assign f[13][60] = 9'b111111111;
assign f[13][61] = 9'b111111111;
assign f[13][62] = 9'b111111111;
assign f[13][63] = 9'b111111111;
assign f[13][64] = 9'b111111111;
assign f[13][65] = 9'b111111111;
assign f[13][66] = 9'b111111111;
assign f[13][67] = 9'b111111111;
assign f[13][68] = 9'b111111111;
assign f[13][69] = 9'b111111111;
assign f[13][70] = 9'b111111111;
assign f[13][71] = 9'b111111111;
assign f[13][72] = 9'b111111111;
assign f[13][73] = 9'b111111111;
assign f[13][74] = 9'b111111111;
assign f[13][75] = 9'b111111111;
assign f[13][76] = 9'b111111111;
assign f[13][77] = 9'b111111111;
assign f[13][78] = 9'b111111111;
assign f[13][79] = 9'b111111111;
assign f[13][80] = 9'b111111111;
assign f[13][81] = 9'b111111111;
assign f[13][82] = 9'b111111111;
assign f[13][83] = 9'b111111111;
assign f[13][84] = 9'b111111111;
assign f[13][85] = 9'b111111111;
assign f[13][86] = 9'b111111111;
assign f[13][87] = 9'b111111111;
assign f[13][88] = 9'b111111111;
assign f[13][89] = 9'b111111111;
assign f[13][90] = 9'b101001000;
assign f[14][36] = 9'b100110101;
assign f[14][37] = 9'b100111101;
assign f[14][38] = 9'b100111101;
assign f[14][39] = 9'b100111101;
assign f[14][40] = 9'b100111101;
assign f[14][41] = 9'b100111101;
assign f[14][42] = 9'b100111101;
assign f[14][43] = 9'b100111101;
assign f[14][44] = 9'b100111101;
assign f[14][45] = 9'b100111101;
assign f[14][46] = 9'b100111101;
assign f[14][47] = 9'b100111101;
assign f[14][48] = 9'b100111101;
assign f[14][49] = 9'b100111101;
assign f[14][50] = 9'b100111101;
assign f[14][51] = 9'b100111101;
assign f[14][52] = 9'b100111101;
assign f[14][53] = 9'b100111101;
assign f[14][54] = 9'b100111101;
assign f[14][55] = 9'b100111101;
assign f[14][56] = 9'b100001001;
assign f[14][57] = 9'b100000000;
assign f[14][58] = 9'b101001001;
assign f[14][59] = 9'b110010001;
assign f[14][60] = 9'b110010001;
assign f[14][61] = 9'b110010001;
assign f[14][62] = 9'b110010001;
assign f[14][63] = 9'b110010001;
assign f[14][64] = 9'b110010001;
assign f[14][65] = 9'b110010001;
assign f[14][66] = 9'b110010001;
assign f[14][67] = 9'b111111111;
assign f[14][68] = 9'b111111111;
assign f[14][69] = 9'b111111111;
assign f[14][70] = 9'b111111111;
assign f[14][71] = 9'b111111111;
assign f[14][72] = 9'b111111111;
assign f[14][73] = 9'b111111111;
assign f[14][74] = 9'b111111111;
assign f[14][75] = 9'b110110110;
assign f[14][76] = 9'b110010001;
assign f[14][77] = 9'b110010001;
assign f[14][78] = 9'b110010001;
assign f[14][79] = 9'b110010001;
assign f[14][80] = 9'b110010001;
assign f[14][81] = 9'b110010001;
assign f[14][82] = 9'b110010001;
assign f[14][83] = 9'b110010001;
assign f[14][84] = 9'b110010001;
assign f[14][85] = 9'b110010001;
assign f[14][86] = 9'b110010001;
assign f[14][87] = 9'b110010001;
assign f[14][88] = 9'b101101101;
assign f[14][89] = 9'b100100100;
assign f[14][90] = 9'b100000000;
assign f[15][36] = 9'b100110101;
assign f[15][37] = 9'b100111101;
assign f[15][38] = 9'b100111101;
assign f[15][39] = 9'b100111101;
assign f[15][40] = 9'b100111101;
assign f[15][41] = 9'b100111101;
assign f[15][42] = 9'b100111101;
assign f[15][43] = 9'b100111101;
assign f[15][44] = 9'b100111101;
assign f[15][45] = 9'b100111101;
assign f[15][46] = 9'b100111101;
assign f[15][47] = 9'b101001101;
assign f[15][48] = 9'b101010101;
assign f[15][49] = 9'b101011101;
assign f[15][50] = 9'b100011101;
assign f[15][51] = 9'b100111101;
assign f[15][52] = 9'b100111101;
assign f[15][53] = 9'b100111101;
assign f[15][54] = 9'b100111101;
assign f[15][55] = 9'b100111101;
assign f[15][58] = 9'b100000000;
assign f[15][59] = 9'b100000000;
assign f[15][60] = 9'b100000000;
assign f[15][61] = 9'b100000000;
assign f[15][62] = 9'b100000000;
assign f[15][63] = 9'b100000000;
assign f[15][64] = 9'b100000000;
assign f[15][65] = 9'b100000000;
assign f[15][66] = 9'b100000000;
assign f[15][67] = 9'b110010010;
assign f[15][68] = 9'b111111111;
assign f[15][69] = 9'b111111111;
assign f[15][70] = 9'b111111111;
assign f[15][71] = 9'b111111111;
assign f[15][72] = 9'b111111111;
assign f[15][73] = 9'b110010010;
assign f[15][74] = 9'b101001000;
assign f[15][75] = 9'b100000000;
assign f[15][76] = 9'b100000000;
assign f[15][77] = 9'b100000000;
assign f[15][78] = 9'b100000000;
assign f[15][79] = 9'b100000000;
assign f[15][80] = 9'b100000000;
assign f[15][81] = 9'b100000000;
assign f[15][82] = 9'b100000000;
assign f[15][83] = 9'b100000000;
assign f[15][84] = 9'b100000000;
assign f[15][85] = 9'b100000000;
assign f[15][86] = 9'b100000000;
assign f[15][87] = 9'b100000000;
assign f[15][88] = 9'b100000000;
assign f[16][36] = 9'b100110101;
assign f[16][37] = 9'b100111101;
assign f[16][38] = 9'b100111101;
assign f[16][39] = 9'b100111101;
assign f[16][40] = 9'b100111101;
assign f[16][41] = 9'b100111101;
assign f[16][42] = 9'b100111101;
assign f[16][43] = 9'b100111101;
assign f[16][44] = 9'b100111101;
assign f[16][45] = 9'b100111101;
assign f[16][46] = 9'b100111101;
assign f[16][47] = 9'b101100100;
assign f[16][48] = 9'b111110001;
assign f[16][49] = 9'b110011111;
assign f[16][50] = 9'b100011101;
assign f[16][51] = 9'b100111101;
assign f[16][52] = 9'b100111101;
assign f[16][53] = 9'b100111101;
assign f[16][54] = 9'b100111101;
assign f[16][55] = 9'b100111101;
assign f[16][56] = 9'b100110101;
assign f[16][66] = 9'b100000000;
assign f[16][67] = 9'b110010010;
assign f[16][68] = 9'b111111111;
assign f[16][69] = 9'b111111111;
assign f[16][70] = 9'b111111111;
assign f[16][71] = 9'b110010001;
assign f[16][72] = 9'b100100100;
assign f[16][73] = 9'b100000000;
assign f[17][36] = 9'b100110101;
assign f[17][37] = 9'b100111101;
assign f[17][38] = 9'b100111101;
assign f[17][39] = 9'b100111101;
assign f[17][40] = 9'b100111101;
assign f[17][41] = 9'b100111101;
assign f[17][42] = 9'b100111101;
assign f[17][43] = 9'b100111101;
assign f[17][44] = 9'b100111101;
assign f[17][45] = 9'b100111101;
assign f[17][46] = 9'b100111101;
assign f[17][47] = 9'b100111101;
assign f[17][48] = 9'b101101101;
assign f[17][49] = 9'b110000000;
assign f[17][50] = 9'b110001000;
assign f[17][51] = 9'b110111111;
assign f[17][52] = 9'b101011101;
assign f[17][53] = 9'b100111101;
assign f[17][54] = 9'b100111101;
assign f[17][55] = 9'b100111101;
assign f[17][56] = 9'b100111101;
assign f[17][57] = 9'b100110101;
assign f[17][66] = 9'b100000000;
assign f[17][67] = 9'b110110110;
assign f[17][68] = 9'b111111111;
assign f[17][69] = 9'b101101101;
assign f[17][70] = 9'b100100100;
assign f[17][71] = 9'b100000000;
assign f[18][36] = 9'b100111101;
assign f[18][37] = 9'b100111101;
assign f[18][38] = 9'b100110001;
assign f[18][39] = 9'b100110001;
assign f[18][40] = 9'b100110101;
assign f[18][41] = 9'b100111101;
assign f[18][42] = 9'b100111101;
assign f[18][43] = 9'b100111101;
assign f[18][44] = 9'b100111101;
assign f[18][45] = 9'b100111101;
assign f[18][46] = 9'b100111101;
assign f[18][47] = 9'b100111101;
assign f[18][48] = 9'b101010001;
assign f[18][49] = 9'b101001000;
assign f[18][50] = 9'b101101101;
assign f[18][51] = 9'b101111110;
assign f[18][52] = 9'b100111101;
assign f[18][53] = 9'b100111101;
assign f[18][54] = 9'b100111101;
assign f[18][55] = 9'b100111101;
assign f[18][56] = 9'b100111101;
assign f[18][57] = 9'b100111101;
assign f[18][58] = 9'b100111101;
assign f[18][59] = 9'b100110101;
assign f[18][66] = 9'b100000000;
assign f[18][67] = 9'b101001000;
assign f[18][68] = 9'b100100100;
assign f[18][69] = 9'b100000000;
assign f[19][36] = 9'b100111101;
assign f[19][37] = 9'b100111101;
assign f[19][38] = 9'b100100000;
assign f[19][39] = 9'b100100000;
assign f[19][40] = 9'b100101101;
assign f[19][41] = 9'b100111101;
assign f[19][42] = 9'b100111101;
assign f[19][43] = 9'b100111101;
assign f[19][44] = 9'b100111101;
assign f[19][45] = 9'b100111101;
assign f[19][46] = 9'b100111101;
assign f[19][47] = 9'b100111101;
assign f[19][48] = 9'b100111101;
assign f[19][49] = 9'b100011101;
assign f[19][50] = 9'b100011101;
assign f[19][51] = 9'b100011101;
assign f[19][52] = 9'b100011101;
assign f[19][53] = 9'b100111101;
assign f[19][54] = 9'b100111101;
assign f[19][55] = 9'b100111101;
assign f[19][56] = 9'b100111101;
assign f[19][57] = 9'b100111101;
assign f[19][58] = 9'b100111101;
assign f[19][59] = 9'b100111101;
assign f[19][66] = 9'b100000000;
assign f[19][67] = 9'b100000000;
assign f[20][36] = 9'b100110001;
assign f[20][37] = 9'b100101000;
assign f[20][38] = 9'b100100000;
assign f[20][39] = 9'b100100000;
assign f[20][40] = 9'b100100100;
assign f[20][41] = 9'b101001000;
assign f[20][42] = 9'b110010001;
assign f[20][43] = 9'b100111101;
assign f[20][44] = 9'b100111101;
assign f[20][45] = 9'b100111101;
assign f[20][46] = 9'b100111101;
assign f[20][47] = 9'b100111101;
assign f[20][48] = 9'b100111101;
assign f[20][49] = 9'b101011101;
assign f[20][50] = 9'b110110001;
assign f[20][51] = 9'b110010001;
assign f[20][52] = 9'b110010001;
assign f[20][53] = 9'b110010001;
assign f[20][54] = 9'b110010001;
assign f[20][55] = 9'b110110001;
assign f[20][56] = 9'b101101000;
assign f[20][57] = 9'b101101000;
assign f[20][58] = 9'b101101000;
assign f[20][59] = 9'b101101000;
assign f[21][36] = 9'b100101000;
assign f[21][37] = 9'b100100000;
assign f[21][38] = 9'b100100000;
assign f[21][39] = 9'b100100000;
assign f[21][40] = 9'b100100000;
assign f[21][41] = 9'b101000000;
assign f[21][42] = 9'b110001001;
assign f[21][43] = 9'b100110001;
assign f[21][44] = 9'b100110001;
assign f[21][45] = 9'b100110001;
assign f[21][46] = 9'b100110001;
assign f[21][47] = 9'b100110001;
assign f[21][48] = 9'b100010001;
assign f[21][49] = 9'b101001101;
assign f[21][50] = 9'b110001001;
assign f[21][51] = 9'b110001001;
assign f[21][52] = 9'b110001001;
assign f[21][53] = 9'b110001001;
assign f[21][54] = 9'b110001001;
assign f[21][55] = 9'b110001001;
assign f[21][56] = 9'b110000100;
assign f[21][57] = 9'b110000000;
assign f[21][58] = 9'b110000000;
assign f[21][59] = 9'b110000000;
assign f[22][35] = 9'b100100000;
assign f[22][36] = 9'b100100000;
assign f[22][37] = 9'b100100000;
assign f[22][38] = 9'b100100000;
assign f[22][39] = 9'b100100000;
assign f[22][40] = 9'b100100000;
assign f[22][41] = 9'b100000000;
assign f[22][42] = 9'b100000000;
assign f[22][43] = 9'b100000000;
assign f[22][44] = 9'b100000000;
assign f[22][45] = 9'b100000000;
assign f[22][46] = 9'b100000000;
assign f[22][47] = 9'b100000000;
assign f[22][48] = 9'b100000000;
assign f[22][49] = 9'b100000000;
assign f[22][50] = 9'b100000000;
assign f[22][51] = 9'b100000000;
assign f[22][52] = 9'b100000000;
assign f[22][53] = 9'b100000000;
assign f[22][54] = 9'b100000000;
assign f[22][55] = 9'b100000000;
assign f[22][56] = 9'b101100100;
assign f[22][57] = 9'b110000100;
assign f[22][58] = 9'b110000100;
assign f[22][59] = 9'b110000100;
assign f[23][34] = 9'b100100100;
assign f[23][35] = 9'b100100000;
assign f[23][36] = 9'b101100100;
assign f[23][37] = 9'b110101101;
assign f[23][38] = 9'b110001101;
assign f[23][39] = 9'b101000100;
assign f[23][40] = 9'b100100000;
assign f[23][41] = 9'b101000100;
assign f[23][42] = 9'b110001101;
assign f[23][43] = 9'b110001101;
assign f[23][44] = 9'b101000100;
assign f[23][45] = 9'b100000000;
assign f[23][46] = 9'b100000000;
assign f[23][47] = 9'b100000000;
assign f[23][48] = 9'b100000000;
assign f[23][49] = 9'b101000100;
assign f[23][50] = 9'b110001101;
assign f[23][51] = 9'b100000000;
assign f[23][52] = 9'b100000000;
assign f[23][53] = 9'b100000000;
assign f[23][54] = 9'b100000000;
assign f[23][55] = 9'b100000000;
assign f[23][56] = 9'b101000100;
assign f[23][57] = 9'b101100101;
assign f[23][58] = 9'b101100101;
assign f[23][59] = 9'b101100101;
assign f[24][34] = 9'b100100000;
assign f[24][35] = 9'b100100000;
assign f[24][36] = 9'b101101000;
assign f[24][37] = 9'b111110001;
assign f[24][38] = 9'b111110001;
assign f[24][39] = 9'b101101000;
assign f[24][40] = 9'b100100000;
assign f[24][41] = 9'b101000100;
assign f[24][42] = 9'b111110001;
assign f[24][43] = 9'b111110001;
assign f[24][44] = 9'b101101000;
assign f[24][45] = 9'b100000000;
assign f[24][46] = 9'b100000000;
assign f[24][47] = 9'b100000000;
assign f[24][48] = 9'b100000000;
assign f[24][49] = 9'b101001000;
assign f[24][50] = 9'b111101101;
assign f[24][51] = 9'b100100000;
assign f[24][52] = 9'b100000000;
assign f[24][53] = 9'b100000000;
assign f[24][54] = 9'b100000000;
assign f[24][55] = 9'b100000000;
assign f[25][34] = 9'b100100000;
assign f[25][35] = 9'b100100000;
assign f[25][36] = 9'b101101000;
assign f[25][37] = 9'b111110001;
assign f[25][38] = 9'b111110001;
assign f[25][39] = 9'b111110001;
assign f[25][40] = 9'b101101000;
assign f[25][41] = 9'b101000100;
assign f[25][42] = 9'b111110001;
assign f[25][43] = 9'b111110001;
assign f[25][44] = 9'b101001000;
assign f[25][45] = 9'b100000000;
assign f[25][46] = 9'b100000000;
assign f[25][47] = 9'b100000000;
assign f[25][48] = 9'b100000000;
assign f[25][49] = 9'b101000100;
assign f[25][50] = 9'b110101101;
assign f[25][51] = 9'b100000000;
assign f[25][52] = 9'b100000000;
assign f[25][53] = 9'b100000000;
assign f[25][54] = 9'b100000000;
assign f[25][55] = 9'b100000000;
assign f[26][34] = 9'b100100000;
assign f[26][35] = 9'b100100000;
assign f[26][36] = 9'b101000100;
assign f[26][37] = 9'b101101000;
assign f[26][38] = 9'b111110001;
assign f[26][39] = 9'b111110001;
assign f[26][40] = 9'b101101000;
assign f[26][41] = 9'b101000100;
assign f[26][42] = 9'b111110001;
assign f[26][43] = 9'b111110001;
assign f[26][44] = 9'b110001101;
assign f[26][45] = 9'b110001001;
assign f[26][46] = 9'b110001001;
assign f[26][47] = 9'b110001001;
assign f[26][48] = 9'b110001001;
assign f[26][49] = 9'b110001101;
assign f[26][50] = 9'b111101101;
assign f[26][51] = 9'b110001001;
assign f[26][52] = 9'b110001001;
assign f[26][53] = 9'b110001001;
assign f[26][54] = 9'b110001001;
assign f[26][55] = 9'b110001101;
assign f[27][34] = 9'b100100000;
assign f[27][35] = 9'b100100000;
assign f[27][36] = 9'b100100000;
assign f[27][37] = 9'b100100000;
assign f[27][38] = 9'b110101101;
assign f[27][39] = 9'b111110001;
assign f[27][40] = 9'b101101000;
assign f[27][41] = 9'b101000100;
assign f[27][42] = 9'b111110001;
assign f[27][43] = 9'b111110001;
assign f[27][44] = 9'b111110001;
assign f[27][45] = 9'b111110001;
assign f[27][46] = 9'b111110001;
assign f[27][47] = 9'b111110001;
assign f[27][48] = 9'b111110001;
assign f[27][49] = 9'b111110001;
assign f[27][50] = 9'b111110001;
assign f[27][51] = 9'b111101101;
assign f[27][52] = 9'b111110001;
assign f[27][53] = 9'b111110001;
assign f[27][54] = 9'b111110001;
assign f[27][55] = 9'b111110001;
assign f[28][34] = 9'b100100000;
assign f[28][35] = 9'b100100000;
assign f[28][36] = 9'b100100000;
assign f[28][37] = 9'b100100000;
assign f[28][38] = 9'b100100000;
assign f[28][39] = 9'b110101101;
assign f[28][40] = 9'b101101000;
assign f[28][41] = 9'b101000100;
assign f[28][42] = 9'b111110001;
assign f[28][43] = 9'b111110001;
assign f[28][44] = 9'b111110001;
assign f[28][45] = 9'b111110001;
assign f[28][46] = 9'b111110001;
assign f[28][47] = 9'b111110001;
assign f[28][48] = 9'b111110001;
assign f[28][49] = 9'b111110001;
assign f[28][50] = 9'b111110001;
assign f[28][51] = 9'b111110001;
assign f[28][52] = 9'b111110001;
assign f[28][53] = 9'b111110001;
assign f[28][54] = 9'b111110001;
assign f[28][55] = 9'b111110001;
assign f[29][34] = 9'b100100000;
assign f[29][35] = 9'b100100000;
assign f[29][36] = 9'b100100000;
assign f[29][37] = 9'b100100000;
assign f[29][38] = 9'b100100000;
assign f[29][39] = 9'b110101101;
assign f[29][40] = 9'b110001101;
assign f[29][41] = 9'b101101000;
assign f[29][42] = 9'b111110001;
assign f[29][43] = 9'b111110001;
assign f[29][44] = 9'b111110001;
assign f[29][45] = 9'b111110001;
assign f[29][46] = 9'b111110001;
assign f[29][47] = 9'b111110001;
assign f[29][48] = 9'b111110001;
assign f[29][49] = 9'b110001101;
assign f[29][50] = 9'b101000100;
assign f[29][51] = 9'b101000100;
assign f[29][52] = 9'b110001101;
assign f[29][53] = 9'b111110001;
assign f[29][54] = 9'b111110001;
assign f[29][55] = 9'b111110001;
assign f[30][34] = 9'b100100100;
assign f[30][35] = 9'b100100000;
assign f[30][36] = 9'b100100000;
assign f[30][37] = 9'b100100000;
assign f[30][38] = 9'b100100000;
assign f[30][39] = 9'b110001101;
assign f[30][40] = 9'b110101101;
assign f[30][41] = 9'b110001000;
assign f[30][42] = 9'b111101101;
assign f[30][43] = 9'b111110001;
assign f[30][44] = 9'b111110001;
assign f[30][45] = 9'b111110001;
assign f[30][46] = 9'b111110001;
assign f[30][47] = 9'b111110001;
assign f[30][48] = 9'b111110001;
assign f[30][49] = 9'b110001001;
assign f[30][50] = 9'b100000000;
assign f[30][51] = 9'b100000000;
assign f[30][52] = 9'b110001101;
assign f[30][53] = 9'b111110001;
assign f[30][54] = 9'b111110001;
assign f[30][55] = 9'b111110001;
assign f[31][35] = 9'b100100000;
assign f[31][36] = 9'b101000000;
assign f[31][37] = 9'b100100000;
assign f[31][38] = 9'b100100000;
assign f[31][39] = 9'b110001101;
assign f[31][40] = 9'b110101101;
assign f[31][41] = 9'b110001000;
assign f[31][42] = 9'b110001000;
assign f[31][43] = 9'b111101101;
assign f[31][44] = 9'b111110001;
assign f[31][45] = 9'b111110001;
assign f[31][46] = 9'b111110001;
assign f[31][47] = 9'b111110001;
assign f[31][48] = 9'b111110001;
assign f[31][49] = 9'b111110001;
assign f[31][50] = 9'b111110001;
assign f[31][51] = 9'b111110001;
assign f[31][52] = 9'b111110001;
assign f[31][53] = 9'b111110001;
assign f[31][54] = 9'b111110001;
assign f[31][55] = 9'b111110001;
assign f[32][35] = 9'b100100100;
assign f[32][36] = 9'b100100100;
assign f[32][37] = 9'b100100000;
assign f[32][38] = 9'b100100000;
assign f[32][39] = 9'b110001101;
assign f[32][40] = 9'b110101101;
assign f[32][41] = 9'b110001000;
assign f[32][42] = 9'b110001000;
assign f[32][43] = 9'b110001101;
assign f[32][44] = 9'b111101101;
assign f[32][45] = 9'b111110001;
assign f[32][46] = 9'b111110001;
assign f[32][47] = 9'b110101101;
assign f[32][48] = 9'b110001101;
assign f[32][49] = 9'b110101101;
assign f[32][50] = 9'b110101101;
assign f[32][51] = 9'b110101101;
assign f[32][52] = 9'b110101101;
assign f[32][53] = 9'b110001101;
assign f[32][54] = 9'b110101101;
assign f[32][55] = 9'b111110001;
assign f[33][36] = 9'b100100100;
assign f[33][37] = 9'b100100000;
assign f[33][38] = 9'b100100000;
assign f[33][39] = 9'b110001101;
assign f[33][40] = 9'b110101101;
assign f[33][41] = 9'b110001000;
assign f[33][42] = 9'b110001000;
assign f[33][43] = 9'b101101000;
assign f[33][44] = 9'b110001101;
assign f[33][45] = 9'b111110001;
assign f[33][46] = 9'b111110001;
assign f[33][47] = 9'b110001000;
assign f[33][48] = 9'b101101000;
assign f[33][49] = 9'b101101000;
assign f[33][50] = 9'b101101000;
assign f[33][51] = 9'b101101000;
assign f[33][52] = 9'b101101000;
assign f[33][53] = 9'b101101000;
assign f[33][54] = 9'b110001000;
assign f[33][55] = 9'b111110001;
assign f[34][38] = 9'b100100000;
assign f[34][39] = 9'b110001101;
assign f[34][40] = 9'b111110001;
assign f[34][41] = 9'b110101101;
assign f[34][42] = 9'b110001000;
assign f[34][43] = 9'b110001000;
assign f[34][44] = 9'b110001000;
assign f[34][45] = 9'b110001101;
assign f[34][46] = 9'b111110001;
assign f[34][47] = 9'b110001000;
assign f[34][48] = 9'b100100000;
assign f[34][49] = 9'b100000000;
assign f[34][50] = 9'b100000000;
assign f[34][51] = 9'b100000000;
assign f[34][52] = 9'b100000000;
assign f[34][53] = 9'b100100100;
assign f[34][54] = 9'b110001101;
assign f[34][55] = 9'b111110001;
assign f[35][38] = 9'b100100000;
assign f[35][39] = 9'b110001101;
assign f[35][40] = 9'b111110001;
assign f[35][41] = 9'b111101101;
assign f[35][42] = 9'b110001101;
assign f[35][43] = 9'b110001000;
assign f[35][44] = 9'b110001000;
assign f[35][45] = 9'b110001000;
assign f[35][46] = 9'b110101101;
assign f[35][47] = 9'b110001000;
assign f[35][48] = 9'b101101000;
assign f[35][49] = 9'b101000100;
assign f[35][50] = 9'b100100100;
assign f[35][51] = 9'b100100100;
assign f[35][52] = 9'b101000100;
assign f[35][53] = 9'b101101000;
assign f[35][54] = 9'b110001000;
assign f[35][55] = 9'b110101101;
assign f[36][38] = 9'b100100000;
assign f[36][39] = 9'b110001101;
assign f[36][40] = 9'b111110001;
assign f[36][41] = 9'b111110001;
assign f[36][42] = 9'b111110001;
assign f[36][43] = 9'b110001000;
assign f[36][44] = 9'b110001000;
assign f[36][45] = 9'b110001000;
assign f[36][46] = 9'b110001000;
assign f[36][47] = 9'b110001000;
assign f[36][48] = 9'b111101101;
assign f[36][49] = 9'b111101101;
assign f[36][50] = 9'b110001000;
assign f[36][51] = 9'b110001000;
assign f[36][52] = 9'b111110001;
assign f[36][53] = 9'b110101101;
assign f[36][54] = 9'b110001000;
assign f[36][55] = 9'b110001000;
assign f[37][39] = 9'b110101101;
assign f[37][40] = 9'b111110001;
assign f[37][41] = 9'b111110001;
assign f[37][42] = 9'b111110001;
assign f[37][43] = 9'b111110001;
assign f[37][44] = 9'b110001001;
assign f[37][45] = 9'b101101000;
assign f[37][46] = 9'b110001000;
assign f[37][47] = 9'b110001000;
assign f[37][48] = 9'b110101101;
assign f[37][49] = 9'b111110001;
assign f[37][50] = 9'b111101101;
assign f[37][51] = 9'b111101101;
assign f[37][52] = 9'b111110001;
assign f[37][53] = 9'b110101101;
assign f[37][54] = 9'b110001000;
assign f[37][55] = 9'b110001000;
assign f[38][39] = 9'b111110001;
assign f[38][40] = 9'b111110001;
assign f[38][41] = 9'b111110001;
assign f[38][42] = 9'b111110001;
assign f[38][43] = 9'b111110001;
assign f[38][44] = 9'b110101101;
assign f[38][45] = 9'b110001000;
assign f[38][46] = 9'b110001000;
assign f[38][47] = 9'b110001000;
assign f[38][48] = 9'b110001101;
assign f[38][49] = 9'b110101101;
assign f[38][50] = 9'b110101101;
assign f[38][51] = 9'b110101101;
assign f[38][52] = 9'b110101101;
assign f[38][53] = 9'b110001101;
assign f[38][54] = 9'b110001000;
assign f[38][55] = 9'b101101001;
assign f[39][39] = 9'b110110001;
assign f[39][40] = 9'b111110001;
assign f[39][41] = 9'b111110001;
assign f[39][42] = 9'b111110001;
assign f[39][43] = 9'b111110001;
assign f[39][44] = 9'b111110001;
assign f[39][45] = 9'b111101101;
assign f[39][46] = 9'b110001000;
assign f[39][47] = 9'b110001000;
assign f[39][48] = 9'b110001000;
assign f[39][49] = 9'b110001000;
assign f[39][50] = 9'b110001000;
assign f[39][51] = 9'b110001000;
assign f[39][52] = 9'b110001000;
assign f[39][53] = 9'b110001000;
assign f[39][54] = 9'b101101001;
assign f[40][39] = 9'b111110001;
assign f[40][40] = 9'b111110001;
assign f[40][41] = 9'b111110001;
assign f[40][42] = 9'b111110001;
assign f[40][43] = 9'b111110001;
assign f[40][44] = 9'b111110001;
assign f[40][45] = 9'b111110001;
assign f[40][46] = 9'b111101101;
assign f[40][47] = 9'b111101101;
assign f[40][48] = 9'b111101101;
assign f[40][49] = 9'b111101101;
assign f[40][50] = 9'b111101101;
assign f[40][51] = 9'b111101101;
assign f[40][52] = 9'b110001101;
assign f[41][38] = 9'b100110001;
assign f[41][39] = 9'b101110001;
assign f[41][40] = 9'b110010001;
assign f[41][41] = 9'b110010001;
assign f[41][42] = 9'b110010001;
assign f[41][43] = 9'b110001101;
assign f[41][44] = 9'b110101101;
assign f[41][45] = 9'b111101101;
assign f[41][46] = 9'b111101101;
assign f[41][47] = 9'b111101101;
assign f[41][48] = 9'b110010001;
assign f[41][49] = 9'b110010001;
assign f[41][50] = 9'b110010001;
assign f[41][51] = 9'b110010001;
assign f[41][52] = 9'b101010001;
assign f[42][38] = 9'b100110001;
assign f[42][39] = 9'b100010001;
assign f[42][40] = 9'b100010001;
assign f[42][41] = 9'b100010001;
assign f[42][42] = 9'b100010001;
assign f[42][43] = 9'b100101101;
assign f[42][44] = 9'b110001001;
assign f[42][45] = 9'b110101001;
assign f[42][46] = 9'b110101001;
assign f[42][47] = 9'b110101001;
assign f[42][48] = 9'b101001101;
assign f[42][49] = 9'b100010001;
assign f[42][50] = 9'b100010001;
assign f[42][51] = 9'b100010001;
assign f[42][52] = 9'b100110001;
assign f[42][53] = 9'b100110001;
assign f[43][30] = 9'b110111111;
assign f[43][31] = 9'b111111111;
assign f[43][32] = 9'b101110111;
assign f[43][33] = 9'b100001111;
assign f[43][34] = 9'b100110001;
assign f[43][35] = 9'b100110001;
assign f[43][36] = 9'b100110001;
assign f[43][37] = 9'b100110001;
assign f[43][38] = 9'b100110001;
assign f[43][39] = 9'b100110001;
assign f[43][40] = 9'b100110001;
assign f[43][41] = 9'b100110001;
assign f[43][42] = 9'b100110001;
assign f[43][43] = 9'b100110001;
assign f[43][44] = 9'b100110001;
assign f[43][45] = 9'b101010001;
assign f[43][46] = 9'b101010001;
assign f[43][47] = 9'b101010001;
assign f[43][48] = 9'b100110001;
assign f[43][49] = 9'b100110001;
assign f[43][50] = 9'b100110001;
assign f[43][51] = 9'b100110001;
assign f[43][52] = 9'b100110001;
assign f[43][53] = 9'b100110001;
assign f[43][54] = 9'b100110001;
assign f[43][55] = 9'b100110001;
assign f[43][56] = 9'b100110001;
assign f[43][57] = 9'b100001101;
assign f[43][58] = 9'b100110011;
assign f[43][59] = 9'b111111111;
assign f[43][60] = 9'b111111111;
assign f[44][30] = 9'b111111111;
assign f[44][31] = 9'b111111111;
assign f[44][32] = 9'b110011111;
assign f[44][33] = 9'b100001111;
assign f[44][34] = 9'b100110001;
assign f[44][35] = 9'b100110001;
assign f[44][36] = 9'b100110001;
assign f[44][37] = 9'b100110001;
assign f[44][38] = 9'b100110001;
assign f[44][39] = 9'b100110001;
assign f[44][40] = 9'b100110001;
assign f[44][41] = 9'b100110001;
assign f[44][42] = 9'b100110001;
assign f[44][43] = 9'b100110001;
assign f[44][44] = 9'b100110001;
assign f[44][45] = 9'b100010001;
assign f[44][46] = 9'b100010001;
assign f[44][47] = 9'b100010001;
assign f[44][48] = 9'b100110001;
assign f[44][49] = 9'b100110001;
assign f[44][50] = 9'b100110001;
assign f[44][51] = 9'b100110001;
assign f[44][52] = 9'b100110001;
assign f[44][53] = 9'b100110001;
assign f[44][54] = 9'b100110001;
assign f[44][55] = 9'b100110001;
assign f[44][56] = 9'b100110001;
assign f[44][57] = 9'b100010010;
assign f[44][58] = 9'b100110011;
assign f[44][59] = 9'b111111111;
assign f[44][60] = 9'b111111111;
assign f[44][61] = 9'b110111111;
assign f[45][30] = 9'b111111111;
assign f[45][31] = 9'b111111111;
assign f[45][32] = 9'b110010111;
assign f[45][33] = 9'b100001111;
assign f[45][34] = 9'b100110001;
assign f[45][35] = 9'b100110001;
assign f[45][36] = 9'b100110001;
assign f[45][37] = 9'b100110001;
assign f[45][38] = 9'b100110001;
assign f[45][39] = 9'b100110001;
assign f[45][40] = 9'b100110001;
assign f[45][41] = 9'b100110001;
assign f[45][42] = 9'b100110001;
assign f[45][43] = 9'b100110001;
assign f[45][44] = 9'b100110001;
assign f[45][45] = 9'b100110001;
assign f[45][46] = 9'b100110001;
assign f[45][47] = 9'b100110001;
assign f[45][48] = 9'b100110001;
assign f[45][49] = 9'b100110001;
assign f[45][50] = 9'b100110001;
assign f[45][51] = 9'b100110001;
assign f[45][52] = 9'b100010001;
assign f[45][53] = 9'b100010001;
assign f[45][54] = 9'b100110001;
assign f[45][55] = 9'b100110001;
assign f[45][56] = 9'b100110001;
assign f[45][57] = 9'b100001101;
assign f[45][58] = 9'b100110011;
assign f[45][59] = 9'b111111111;
assign f[45][60] = 9'b111111111;
assign f[45][61] = 9'b110111111;
assign f[46][30] = 9'b111111111;
assign f[46][31] = 9'b111111111;
assign f[46][32] = 9'b110011111;
assign f[46][33] = 9'b100001111;
assign f[46][34] = 9'b100110001;
assign f[46][35] = 9'b100110001;
assign f[46][36] = 9'b100110001;
assign f[46][37] = 9'b100110001;
assign f[46][38] = 9'b100110001;
assign f[46][39] = 9'b100110001;
assign f[46][40] = 9'b100110001;
assign f[46][41] = 9'b100110001;
assign f[46][42] = 9'b100110001;
assign f[46][43] = 9'b100110001;
assign f[46][44] = 9'b100110001;
assign f[46][45] = 9'b100110001;
assign f[46][46] = 9'b100110001;
assign f[46][47] = 9'b100110001;
assign f[46][48] = 9'b100110001;
assign f[46][49] = 9'b100110001;
assign f[46][50] = 9'b100110001;
assign f[46][51] = 9'b100010001;
assign f[46][52] = 9'b110011110;
assign f[46][53] = 9'b101111110;
assign f[46][54] = 9'b100010001;
assign f[46][55] = 9'b100110001;
assign f[46][56] = 9'b100110001;
assign f[46][57] = 9'b100010001;
assign f[46][58] = 9'b100110011;
assign f[46][59] = 9'b111111111;
assign f[46][60] = 9'b111111111;
assign f[46][61] = 9'b110111111;
assign f[47][30] = 9'b111111111;
assign f[47][31] = 9'b111111111;
assign f[47][32] = 9'b110010111;
assign f[47][33] = 9'b100001111;
assign f[47][34] = 9'b100110001;
assign f[47][35] = 9'b100110001;
assign f[47][36] = 9'b100110001;
assign f[47][37] = 9'b100110001;
assign f[47][38] = 9'b100110001;
assign f[47][39] = 9'b100110001;
assign f[47][40] = 9'b100110001;
assign f[47][41] = 9'b100110001;
assign f[47][42] = 9'b100110001;
assign f[47][43] = 9'b100110001;
assign f[47][44] = 9'b100110001;
assign f[47][45] = 9'b100110001;
assign f[47][46] = 9'b100110001;
assign f[47][47] = 9'b100110001;
assign f[47][48] = 9'b100110001;
assign f[47][49] = 9'b100110001;
assign f[47][50] = 9'b100110001;
assign f[47][51] = 9'b100010001;
assign f[47][52] = 9'b111111111;
assign f[47][53] = 9'b110111111;
assign f[47][54] = 9'b100010001;
assign f[47][55] = 9'b100110001;
assign f[47][56] = 9'b100110001;
assign f[47][57] = 9'b100010001;
assign f[47][58] = 9'b101010011;
assign f[47][59] = 9'b111111111;
assign f[47][60] = 9'b111111111;
assign f[47][61] = 9'b110111111;
//Total de Lineas = 1350
endmodule

