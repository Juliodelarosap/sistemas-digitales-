`timescale 1ns / 1ps
module nombre (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (no[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= no[vcount- posy][hcount- posx][7:5];
				green <= no[vcount- posy][hcount- posx][4:2];
            blue 	<= no[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 150;
parameter RESOLUCION_Y = 50;
wire [8:0] no[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign no[15][32] = 9'b111111111;
assign no[15][33] = 9'b111111111;
assign no[15][34] = 9'b111111111;
assign no[15][35] = 9'b111111111;
assign no[15][42] = 9'b111111111;
assign no[15][43] = 9'b111111111;
assign no[15][44] = 9'b111111111;
assign no[15][45] = 9'b111111111;
assign no[15][46] = 9'b111111111;
assign no[15][50] = 9'b111111111;
assign no[15][51] = 9'b111111111;
assign no[15][52] = 9'b111111111;
assign no[15][53] = 9'b111111111;
assign no[15][54] = 9'b111111111;
assign no[15][55] = 9'b111111111;
assign no[15][56] = 9'b111111111;
assign no[15][57] = 9'b111111111;
assign no[15][58] = 9'b111111111;
assign no[15][59] = 9'b111111111;
assign no[15][60] = 9'b111111111;
assign no[15][75] = 9'b111111111;
assign no[15][76] = 9'b111111111;
assign no[15][77] = 9'b111111111;
assign no[15][78] = 9'b111111111;
assign no[15][88] = 9'b111111111;
assign no[15][89] = 9'b111111111;
assign no[15][90] = 9'b111111111;
assign no[15][91] = 9'b111111111;
assign no[15][110] = 9'b111111111;
assign no[15][111] = 9'b111111111;
assign no[15][112] = 9'b111111111;
assign no[15][113] = 9'b111111111;
assign no[15][114] = 9'b111111111;
assign no[15][123] = 9'b111111111;
assign no[15][124] = 9'b111111111;
assign no[15][125] = 9'b111111111;
assign no[15][126] = 9'b111111111;
assign no[15][127] = 9'b111111111;
assign no[15][128] = 9'b111111111;
assign no[15][135] = 9'b111111111;
assign no[15][136] = 9'b111111111;
assign no[16][14] = 9'b111111111;
assign no[16][15] = 9'b111111111;
assign no[16][16] = 9'b111111111;
assign no[16][17] = 9'b111111111;
assign no[16][18] = 9'b111111111;
assign no[16][19] = 9'b111111111;
assign no[16][20] = 9'b111111111;
assign no[16][21] = 9'b111111111;
assign no[16][22] = 9'b111111111;
assign no[16][23] = 9'b111111111;
assign no[16][24] = 9'b111111111;
assign no[16][25] = 9'b111111111;
assign no[16][26] = 9'b111111111;
assign no[16][27] = 9'b111111111;
assign no[16][28] = 9'b111111111;
assign no[16][29] = 9'b111111111;
assign no[16][31] = 9'b111111111;
assign no[16][32] = 9'b111111111;
assign no[16][33] = 9'b111111111;
assign no[16][34] = 9'b111111111;
assign no[16][35] = 9'b111111111;
assign no[16][36] = 9'b111111111;
assign no[16][42] = 9'b111111111;
assign no[16][43] = 9'b111111111;
assign no[16][44] = 9'b111111111;
assign no[16][45] = 9'b111111111;
assign no[16][46] = 9'b111111111;
assign no[16][49] = 9'b111111111;
assign no[16][50] = 9'b111111111;
assign no[16][51] = 9'b111111111;
assign no[16][52] = 9'b111111111;
assign no[16][53] = 9'b111111111;
assign no[16][54] = 9'b111111111;
assign no[16][55] = 9'b111111111;
assign no[16][56] = 9'b111111111;
assign no[16][57] = 9'b111111111;
assign no[16][58] = 9'b111111111;
assign no[16][59] = 9'b111111111;
assign no[16][60] = 9'b111111111;
assign no[16][61] = 9'b111111111;
assign no[16][70] = 9'b111111111;
assign no[16][71] = 9'b111111111;
assign no[16][72] = 9'b111111111;
assign no[16][73] = 9'b111111111;
assign no[16][74] = 9'b111111111;
assign no[16][75] = 9'b111111111;
assign no[16][76] = 9'b111111111;
assign no[16][77] = 9'b111111111;
assign no[16][78] = 9'b111111111;
assign no[16][79] = 9'b111111111;
assign no[16][80] = 9'b111111111;
assign no[16][81] = 9'b111111111;
assign no[16][82] = 9'b111111111;
assign no[16][83] = 9'b111111111;
assign no[16][88] = 9'b111111111;
assign no[16][89] = 9'b111111111;
assign no[16][90] = 9'b111111111;
assign no[16][91] = 9'b111111111;
assign no[16][92] = 9'b111111111;
assign no[16][109] = 9'b111111111;
assign no[16][110] = 9'b111111111;
assign no[16][111] = 9'b111111111;
assign no[16][112] = 9'b111111111;
assign no[16][113] = 9'b111111111;
assign no[16][114] = 9'b111111111;
assign no[16][115] = 9'b111111111;
assign no[16][123] = 9'b111111111;
assign no[16][124] = 9'b111111111;
assign no[16][125] = 9'b111111111;
assign no[16][126] = 9'b111111111;
assign no[16][127] = 9'b111111111;
assign no[16][128] = 9'b111111111;
assign no[16][129] = 9'b111111111;
assign no[16][135] = 9'b111111111;
assign no[16][136] = 9'b111111111;
assign no[16][137] = 9'b111111111;
assign no[16][138] = 9'b111111111;
assign no[17][14] = 9'b111111111;
assign no[17][15] = 9'b111111111;
assign no[17][16] = 9'b111111111;
assign no[17][17] = 9'b111111111;
assign no[17][18] = 9'b111111111;
assign no[17][19] = 9'b111111111;
assign no[17][20] = 9'b111111111;
assign no[17][21] = 9'b111111111;
assign no[17][22] = 9'b111111111;
assign no[17][23] = 9'b111111111;
assign no[17][24] = 9'b111111111;
assign no[17][25] = 9'b111111111;
assign no[17][26] = 9'b111111111;
assign no[17][27] = 9'b111111111;
assign no[17][28] = 9'b111111111;
assign no[17][29] = 9'b111111111;
assign no[17][31] = 9'b111111111;
assign no[17][32] = 9'b111111111;
assign no[17][33] = 9'b111111111;
assign no[17][34] = 9'b111111111;
assign no[17][35] = 9'b111111111;
assign no[17][36] = 9'b111111111;
assign no[17][42] = 9'b111111111;
assign no[17][43] = 9'b111111111;
assign no[17][44] = 9'b111111111;
assign no[17][45] = 9'b111111111;
assign no[17][46] = 9'b111111111;
assign no[17][49] = 9'b111111111;
assign no[17][50] = 9'b111111111;
assign no[17][51] = 9'b111111111;
assign no[17][52] = 9'b111111111;
assign no[17][53] = 9'b111111111;
assign no[17][54] = 9'b111111111;
assign no[17][55] = 9'b111111111;
assign no[17][56] = 9'b111111111;
assign no[17][57] = 9'b111111111;
assign no[17][58] = 9'b111111111;
assign no[17][59] = 9'b111111111;
assign no[17][60] = 9'b111111111;
assign no[17][61] = 9'b111111111;
assign no[17][70] = 9'b111111111;
assign no[17][71] = 9'b111111111;
assign no[17][72] = 9'b111111111;
assign no[17][73] = 9'b111111111;
assign no[17][74] = 9'b111111111;
assign no[17][75] = 9'b111111111;
assign no[17][76] = 9'b111111111;
assign no[17][77] = 9'b111111111;
assign no[17][78] = 9'b111111111;
assign no[17][79] = 9'b111111111;
assign no[17][80] = 9'b111111111;
assign no[17][81] = 9'b111111111;
assign no[17][82] = 9'b111111111;
assign no[17][83] = 9'b111111111;
assign no[17][84] = 9'b111111111;
assign no[17][88] = 9'b111111111;
assign no[17][89] = 9'b111111111;
assign no[17][90] = 9'b111111111;
assign no[17][91] = 9'b111111111;
assign no[17][92] = 9'b111111111;
assign no[17][109] = 9'b111111111;
assign no[17][110] = 9'b111111111;
assign no[17][111] = 9'b111111111;
assign no[17][112] = 9'b111111111;
assign no[17][113] = 9'b111111111;
assign no[17][114] = 9'b111111111;
assign no[17][115] = 9'b111111111;
assign no[17][123] = 9'b111111111;
assign no[17][124] = 9'b111111111;
assign no[17][125] = 9'b111111111;
assign no[17][126] = 9'b111111111;
assign no[17][127] = 9'b111111111;
assign no[17][128] = 9'b111111111;
assign no[17][129] = 9'b111111111;
assign no[17][130] = 9'b111111111;
assign no[17][135] = 9'b111111111;
assign no[17][136] = 9'b111111111;
assign no[17][137] = 9'b111111111;
assign no[17][138] = 9'b111111111;
assign no[18][15] = 9'b111111111;
assign no[18][16] = 9'b111111111;
assign no[18][17] = 9'b111111111;
assign no[18][18] = 9'b111111111;
assign no[18][19] = 9'b111111111;
assign no[18][20] = 9'b111111111;
assign no[18][21] = 9'b111111111;
assign no[18][22] = 9'b111111111;
assign no[18][23] = 9'b111111111;
assign no[18][24] = 9'b111111111;
assign no[18][25] = 9'b111111111;
assign no[18][26] = 9'b111111111;
assign no[18][27] = 9'b111111111;
assign no[18][28] = 9'b111111111;
assign no[18][29] = 9'b111111111;
assign no[18][31] = 9'b111111111;
assign no[18][32] = 9'b111111111;
assign no[18][33] = 9'b111111111;
assign no[18][34] = 9'b111111111;
assign no[18][35] = 9'b111111111;
assign no[18][36] = 9'b111111111;
assign no[18][42] = 9'b111111111;
assign no[18][43] = 9'b111111111;
assign no[18][44] = 9'b111111111;
assign no[18][45] = 9'b111111111;
assign no[18][46] = 9'b111111111;
assign no[18][49] = 9'b111111111;
assign no[18][50] = 9'b111111111;
assign no[18][51] = 9'b111111111;
assign no[18][52] = 9'b111111111;
assign no[18][53] = 9'b111111111;
assign no[18][54] = 9'b111111111;
assign no[18][56] = 9'b111111111;
assign no[18][70] = 9'b111111111;
assign no[18][71] = 9'b111111111;
assign no[18][72] = 9'b111111111;
assign no[18][73] = 9'b111111111;
assign no[18][74] = 9'b111111111;
assign no[18][75] = 9'b111111111;
assign no[18][76] = 9'b111111111;
assign no[18][77] = 9'b111111111;
assign no[18][78] = 9'b111111111;
assign no[18][79] = 9'b111111111;
assign no[18][80] = 9'b111111111;
assign no[18][81] = 9'b111111111;
assign no[18][82] = 9'b111111111;
assign no[18][83] = 9'b111111111;
assign no[18][84] = 9'b111111111;
assign no[18][88] = 9'b111111111;
assign no[18][89] = 9'b111111111;
assign no[18][90] = 9'b111111111;
assign no[18][91] = 9'b111111111;
assign no[18][92] = 9'b111111111;
assign no[18][108] = 9'b111111111;
assign no[18][109] = 9'b111111111;
assign no[18][110] = 9'b111111111;
assign no[18][111] = 9'b111111111;
assign no[18][112] = 9'b111111111;
assign no[18][113] = 9'b111111111;
assign no[18][114] = 9'b111111111;
assign no[18][115] = 9'b111111111;
assign no[18][116] = 9'b111111111;
assign no[18][123] = 9'b111111111;
assign no[18][124] = 9'b111111111;
assign no[18][125] = 9'b111111111;
assign no[18][126] = 9'b111111111;
assign no[18][127] = 9'b111111111;
assign no[18][128] = 9'b111111111;
assign no[18][129] = 9'b111111111;
assign no[18][130] = 9'b111111111;
assign no[18][135] = 9'b111111111;
assign no[18][136] = 9'b111111111;
assign no[18][137] = 9'b111111111;
assign no[18][138] = 9'b111111111;
assign no[19][20] = 9'b111111111;
assign no[19][21] = 9'b111111111;
assign no[19][22] = 9'b111111111;
assign no[19][23] = 9'b111111111;
assign no[19][24] = 9'b111111111;
assign no[19][31] = 9'b111111111;
assign no[19][32] = 9'b111111111;
assign no[19][33] = 9'b111111111;
assign no[19][34] = 9'b111111111;
assign no[19][35] = 9'b111111111;
assign no[19][36] = 9'b111111111;
assign no[19][42] = 9'b111111111;
assign no[19][43] = 9'b111111111;
assign no[19][44] = 9'b111111111;
assign no[19][45] = 9'b111111111;
assign no[19][46] = 9'b111111111;
assign no[19][49] = 9'b111111111;
assign no[19][50] = 9'b111111111;
assign no[19][51] = 9'b111111111;
assign no[19][52] = 9'b111111111;
assign no[19][53] = 9'b111111111;
assign no[19][70] = 9'b111111111;
assign no[19][71] = 9'b111111111;
assign no[19][72] = 9'b111111111;
assign no[19][73] = 9'b111111111;
assign no[19][74] = 9'b111111111;
assign no[19][75] = 9'b111111111;
assign no[19][80] = 9'b111111111;
assign no[19][81] = 9'b111111111;
assign no[19][82] = 9'b111111111;
assign no[19][83] = 9'b111111111;
assign no[19][84] = 9'b111111111;
assign no[19][85] = 9'b111111111;
assign no[19][88] = 9'b111111111;
assign no[19][89] = 9'b111111111;
assign no[19][90] = 9'b111111111;
assign no[19][91] = 9'b111111111;
assign no[19][92] = 9'b111111111;
assign no[19][107] = 9'b111111111;
assign no[19][108] = 9'b111111111;
assign no[19][109] = 9'b111111111;
assign no[19][110] = 9'b111111111;
assign no[19][111] = 9'b111111111;
assign no[19][112] = 9'b111111111;
assign no[19][113] = 9'b111111111;
assign no[19][114] = 9'b111111111;
assign no[19][115] = 9'b111111111;
assign no[19][116] = 9'b111111111;
assign no[19][123] = 9'b111111111;
assign no[19][124] = 9'b111111111;
assign no[19][125] = 9'b111111111;
assign no[19][126] = 9'b111111111;
assign no[19][127] = 9'b111111111;
assign no[19][128] = 9'b111111111;
assign no[19][129] = 9'b111111111;
assign no[19][130] = 9'b111111111;
assign no[19][135] = 9'b111111111;
assign no[19][136] = 9'b111111111;
assign no[19][137] = 9'b111111111;
assign no[19][138] = 9'b111111111;
assign no[20][20] = 9'b111111111;
assign no[20][21] = 9'b111111111;
assign no[20][22] = 9'b111111111;
assign no[20][23] = 9'b111111111;
assign no[20][24] = 9'b111111111;
assign no[20][31] = 9'b111111111;
assign no[20][32] = 9'b111111111;
assign no[20][33] = 9'b111111111;
assign no[20][34] = 9'b111111111;
assign no[20][35] = 9'b111111111;
assign no[20][36] = 9'b111111111;
assign no[20][42] = 9'b111111111;
assign no[20][43] = 9'b111111111;
assign no[20][44] = 9'b111111111;
assign no[20][45] = 9'b111111111;
assign no[20][46] = 9'b111111111;
assign no[20][49] = 9'b111111111;
assign no[20][50] = 9'b111111111;
assign no[20][51] = 9'b111111111;
assign no[20][52] = 9'b111111111;
assign no[20][53] = 9'b111111111;
assign no[20][71] = 9'b111111111;
assign no[20][72] = 9'b111111111;
assign no[20][73] = 9'b111111111;
assign no[20][74] = 9'b111111111;
assign no[20][75] = 9'b111111111;
assign no[20][80] = 9'b111111111;
assign no[20][81] = 9'b111111111;
assign no[20][82] = 9'b111111111;
assign no[20][83] = 9'b111111111;
assign no[20][84] = 9'b111111111;
assign no[20][85] = 9'b111111111;
assign no[20][88] = 9'b111111111;
assign no[20][89] = 9'b111111111;
assign no[20][90] = 9'b111111111;
assign no[20][91] = 9'b111111111;
assign no[20][92] = 9'b111111111;
assign no[20][107] = 9'b111111111;
assign no[20][109] = 9'b111111111;
assign no[20][110] = 9'b111111111;
assign no[20][113] = 9'b111111111;
assign no[20][114] = 9'b111111111;
assign no[20][115] = 9'b111111111;
assign no[20][116] = 9'b111111111;
assign no[20][122] = 9'b111111111;
assign no[20][123] = 9'b111111111;
assign no[20][124] = 9'b111111111;
assign no[20][125] = 9'b111111111;
assign no[20][126] = 9'b111111111;
assign no[20][127] = 9'b111111111;
assign no[20][128] = 9'b111111111;
assign no[20][129] = 9'b111111111;
assign no[20][130] = 9'b111111111;
assign no[20][131] = 9'b111111111;
assign no[20][135] = 9'b111111111;
assign no[20][136] = 9'b111111111;
assign no[20][137] = 9'b111111111;
assign no[20][138] = 9'b111111111;
assign no[21][20] = 9'b111111111;
assign no[21][21] = 9'b111111111;
assign no[21][22] = 9'b111111111;
assign no[21][23] = 9'b111111111;
assign no[21][24] = 9'b111111111;
assign no[21][31] = 9'b111111111;
assign no[21][32] = 9'b111111111;
assign no[21][33] = 9'b111111111;
assign no[21][34] = 9'b111111111;
assign no[21][35] = 9'b111111111;
assign no[21][36] = 9'b111111111;
assign no[21][42] = 9'b111111111;
assign no[21][43] = 9'b111111111;
assign no[21][44] = 9'b111111111;
assign no[21][45] = 9'b111111111;
assign no[21][46] = 9'b111111111;
assign no[21][49] = 9'b111111111;
assign no[21][50] = 9'b111111111;
assign no[21][51] = 9'b111111111;
assign no[21][52] = 9'b111111111;
assign no[21][53] = 9'b111111111;
assign no[21][70] = 9'b111111111;
assign no[21][71] = 9'b111111111;
assign no[21][72] = 9'b111111111;
assign no[21][73] = 9'b111111111;
assign no[21][74] = 9'b111111111;
assign no[21][75] = 9'b111111111;
assign no[21][80] = 9'b111111111;
assign no[21][81] = 9'b111111111;
assign no[21][82] = 9'b111111111;
assign no[21][83] = 9'b111111111;
assign no[21][84] = 9'b111111111;
assign no[21][85] = 9'b111111111;
assign no[21][88] = 9'b111111111;
assign no[21][89] = 9'b111111111;
assign no[21][90] = 9'b111111111;
assign no[21][91] = 9'b111111111;
assign no[21][92] = 9'b111111111;
assign no[21][107] = 9'b111111111;
assign no[21][110] = 9'b111111111;
assign no[21][113] = 9'b111111111;
assign no[21][114] = 9'b111111111;
assign no[21][115] = 9'b111111111;
assign no[21][116] = 9'b111111111;
assign no[21][117] = 9'b111111111;
assign no[21][123] = 9'b111111111;
assign no[21][124] = 9'b111111111;
assign no[21][125] = 9'b111111111;
assign no[21][126] = 9'b111111111;
assign no[21][127] = 9'b111111111;
assign no[21][128] = 9'b111111111;
assign no[21][129] = 9'b111111111;
assign no[21][130] = 9'b111111111;
assign no[21][131] = 9'b111111111;
assign no[21][135] = 9'b111111111;
assign no[21][136] = 9'b111111111;
assign no[21][137] = 9'b111111111;
assign no[21][138] = 9'b111111111;
assign no[22][20] = 9'b111111111;
assign no[22][21] = 9'b111111111;
assign no[22][22] = 9'b111111111;
assign no[22][23] = 9'b111111111;
assign no[22][24] = 9'b111111111;
assign no[22][31] = 9'b111111111;
assign no[22][32] = 9'b111111111;
assign no[22][33] = 9'b111111111;
assign no[22][34] = 9'b111111111;
assign no[22][35] = 9'b111111111;
assign no[22][36] = 9'b111111111;
assign no[22][37] = 9'b111111111;
assign no[22][38] = 9'b111111111;
assign no[22][41] = 9'b111111111;
assign no[22][42] = 9'b111111111;
assign no[22][43] = 9'b111111111;
assign no[22][44] = 9'b111111111;
assign no[22][45] = 9'b111111111;
assign no[22][46] = 9'b111111111;
assign no[22][49] = 9'b111111111;
assign no[22][50] = 9'b111111111;
assign no[22][51] = 9'b111111111;
assign no[22][52] = 9'b111111111;
assign no[22][53] = 9'b111111111;
assign no[22][54] = 9'b111111111;
assign no[22][55] = 9'b111111111;
assign no[22][56] = 9'b111111111;
assign no[22][57] = 9'b111111111;
assign no[22][58] = 9'b111111111;
assign no[22][59] = 9'b111111111;
assign no[22][60] = 9'b111111111;
assign no[22][70] = 9'b111111111;
assign no[22][71] = 9'b111111111;
assign no[22][72] = 9'b111111111;
assign no[22][73] = 9'b111111111;
assign no[22][74] = 9'b111111111;
assign no[22][75] = 9'b111111111;
assign no[22][80] = 9'b111111111;
assign no[22][81] = 9'b111111111;
assign no[22][82] = 9'b111111111;
assign no[22][83] = 9'b111111111;
assign no[22][84] = 9'b111111111;
assign no[22][85] = 9'b111111111;
assign no[22][88] = 9'b111111111;
assign no[22][89] = 9'b111111111;
assign no[22][90] = 9'b111111111;
assign no[22][91] = 9'b111111111;
assign no[22][92] = 9'b111111111;
assign no[22][107] = 9'b111111111;
assign no[22][108] = 9'b111111111;
assign no[22][109] = 9'b111111111;
assign no[22][113] = 9'b111111111;
assign no[22][114] = 9'b111111111;
assign no[22][115] = 9'b111111111;
assign no[22][116] = 9'b111111111;
assign no[22][117] = 9'b111111111;
assign no[22][123] = 9'b111111111;
assign no[22][124] = 9'b111111111;
assign no[22][125] = 9'b111111111;
assign no[22][126] = 9'b111111111;
assign no[22][128] = 9'b111111111;
assign no[22][129] = 9'b111111111;
assign no[22][130] = 9'b111111111;
assign no[22][131] = 9'b111111111;
assign no[22][132] = 9'b111111111;
assign no[22][135] = 9'b111111111;
assign no[22][136] = 9'b111111111;
assign no[22][137] = 9'b111111111;
assign no[22][138] = 9'b111111111;
assign no[23][20] = 9'b111111111;
assign no[23][21] = 9'b111111111;
assign no[23][22] = 9'b111111111;
assign no[23][23] = 9'b111111111;
assign no[23][24] = 9'b111111111;
assign no[23][31] = 9'b111111111;
assign no[23][32] = 9'b111111111;
assign no[23][33] = 9'b111111111;
assign no[23][34] = 9'b111111111;
assign no[23][35] = 9'b111111111;
assign no[23][36] = 9'b111111111;
assign no[23][37] = 9'b111111111;
assign no[23][38] = 9'b111111111;
assign no[23][39] = 9'b111111111;
assign no[23][40] = 9'b111111111;
assign no[23][41] = 9'b111111111;
assign no[23][42] = 9'b111111111;
assign no[23][43] = 9'b111111111;
assign no[23][44] = 9'b111111111;
assign no[23][45] = 9'b111111111;
assign no[23][46] = 9'b111111111;
assign no[23][49] = 9'b111111111;
assign no[23][50] = 9'b111111111;
assign no[23][51] = 9'b111111111;
assign no[23][52] = 9'b111111111;
assign no[23][53] = 9'b111111111;
assign no[23][54] = 9'b111111111;
assign no[23][55] = 9'b111111111;
assign no[23][56] = 9'b111111111;
assign no[23][57] = 9'b111111111;
assign no[23][58] = 9'b111111111;
assign no[23][59] = 9'b111111111;
assign no[23][60] = 9'b111111111;
assign no[23][71] = 9'b111111111;
assign no[23][72] = 9'b111111111;
assign no[23][73] = 9'b111111111;
assign no[23][74] = 9'b111111111;
assign no[23][75] = 9'b111111111;
assign no[23][76] = 9'b111111111;
assign no[23][77] = 9'b111111111;
assign no[23][78] = 9'b111111111;
assign no[23][79] = 9'b111111111;
assign no[23][80] = 9'b111111111;
assign no[23][81] = 9'b111111111;
assign no[23][82] = 9'b111111111;
assign no[23][83] = 9'b111111111;
assign no[23][84] = 9'b111111111;
assign no[23][88] = 9'b111111111;
assign no[23][89] = 9'b111111111;
assign no[23][90] = 9'b111111111;
assign no[23][91] = 9'b111111111;
assign no[23][92] = 9'b111111111;
assign no[23][107] = 9'b111111111;
assign no[23][109] = 9'b111111111;
assign no[23][113] = 9'b111111111;
assign no[23][114] = 9'b111111111;
assign no[23][115] = 9'b111111111;
assign no[23][116] = 9'b111111111;
assign no[23][117] = 9'b111111111;
assign no[23][118] = 9'b111111111;
assign no[23][122] = 9'b111111111;
assign no[23][123] = 9'b111111111;
assign no[23][124] = 9'b111111111;
assign no[23][125] = 9'b111111111;
assign no[23][126] = 9'b111111111;
assign no[23][128] = 9'b111111111;
assign no[23][129] = 9'b111111111;
assign no[23][130] = 9'b111111111;
assign no[23][131] = 9'b111111111;
assign no[23][132] = 9'b111111111;
assign no[23][135] = 9'b111111111;
assign no[23][136] = 9'b111111111;
assign no[23][137] = 9'b111111111;
assign no[23][138] = 9'b111111111;
assign no[24][20] = 9'b111111111;
assign no[24][21] = 9'b111111111;
assign no[24][22] = 9'b111111111;
assign no[24][23] = 9'b111111111;
assign no[24][24] = 9'b111111111;
assign no[24][31] = 9'b111111111;
assign no[24][32] = 9'b111111111;
assign no[24][33] = 9'b111111111;
assign no[24][34] = 9'b111111111;
assign no[24][35] = 9'b111111111;
assign no[24][36] = 9'b111111111;
assign no[24][37] = 9'b111111111;
assign no[24][38] = 9'b111111111;
assign no[24][39] = 9'b111111111;
assign no[24][40] = 9'b111111111;
assign no[24][41] = 9'b111111111;
assign no[24][42] = 9'b111111111;
assign no[24][43] = 9'b111111111;
assign no[24][44] = 9'b111111111;
assign no[24][45] = 9'b111111111;
assign no[24][46] = 9'b111111111;
assign no[24][49] = 9'b111111111;
assign no[24][50] = 9'b111111111;
assign no[24][51] = 9'b111111111;
assign no[24][52] = 9'b111111111;
assign no[24][53] = 9'b111111111;
assign no[24][54] = 9'b111111111;
assign no[24][55] = 9'b111111111;
assign no[24][56] = 9'b111111111;
assign no[24][57] = 9'b111111111;
assign no[24][58] = 9'b111111111;
assign no[24][59] = 9'b111111111;
assign no[24][60] = 9'b111111111;
assign no[24][71] = 9'b111111111;
assign no[24][72] = 9'b111111111;
assign no[24][73] = 9'b111111111;
assign no[24][74] = 9'b111111111;
assign no[24][75] = 9'b111111111;
assign no[24][76] = 9'b111111111;
assign no[24][77] = 9'b111111111;
assign no[24][78] = 9'b111111111;
assign no[24][79] = 9'b111111111;
assign no[24][80] = 9'b111111111;
assign no[24][81] = 9'b111111111;
assign no[24][82] = 9'b111111111;
assign no[24][83] = 9'b111111111;
assign no[24][84] = 9'b111111111;
assign no[24][88] = 9'b111111111;
assign no[24][89] = 9'b111111111;
assign no[24][90] = 9'b111111111;
assign no[24][91] = 9'b111111111;
assign no[24][92] = 9'b111111111;
assign no[24][106] = 9'b111111111;
assign no[24][107] = 9'b111111111;
assign no[24][108] = 9'b111111111;
assign no[24][109] = 9'b111111111;
assign no[24][114] = 9'b111111111;
assign no[24][115] = 9'b111111111;
assign no[24][116] = 9'b111111111;
assign no[24][117] = 9'b111111111;
assign no[24][118] = 9'b111111111;
assign no[24][123] = 9'b111111111;
assign no[24][124] = 9'b111111111;
assign no[24][125] = 9'b111111111;
assign no[24][126] = 9'b111111111;
assign no[24][129] = 9'b111111111;
assign no[24][130] = 9'b111111111;
assign no[24][131] = 9'b111111111;
assign no[24][132] = 9'b111111111;
assign no[24][135] = 9'b111111111;
assign no[24][136] = 9'b111111111;
assign no[24][137] = 9'b111111111;
assign no[24][138] = 9'b111111111;
assign no[25][20] = 9'b111111111;
assign no[25][21] = 9'b111111111;
assign no[25][22] = 9'b111111111;
assign no[25][23] = 9'b111111111;
assign no[25][24] = 9'b111111111;
assign no[25][31] = 9'b111111111;
assign no[25][32] = 9'b111111111;
assign no[25][33] = 9'b111111111;
assign no[25][34] = 9'b111111111;
assign no[25][35] = 9'b111111111;
assign no[25][36] = 9'b111111111;
assign no[25][41] = 9'b111111111;
assign no[25][42] = 9'b111111111;
assign no[25][43] = 9'b111111111;
assign no[25][44] = 9'b111111111;
assign no[25][45] = 9'b111111111;
assign no[25][46] = 9'b111111111;
assign no[25][49] = 9'b111111111;
assign no[25][50] = 9'b111111111;
assign no[25][51] = 9'b111111111;
assign no[25][52] = 9'b111111111;
assign no[25][53] = 9'b111111111;
assign no[25][54] = 9'b111111111;
assign no[25][70] = 9'b111111111;
assign no[25][71] = 9'b111111111;
assign no[25][72] = 9'b111111111;
assign no[25][73] = 9'b111111111;
assign no[25][74] = 9'b111111111;
assign no[25][75] = 9'b111111111;
assign no[25][76] = 9'b111111111;
assign no[25][77] = 9'b111111111;
assign no[25][78] = 9'b111111111;
assign no[25][79] = 9'b111111111;
assign no[25][80] = 9'b111111111;
assign no[25][81] = 9'b111111111;
assign no[25][82] = 9'b111111111;
assign no[25][88] = 9'b111111111;
assign no[25][89] = 9'b111111111;
assign no[25][90] = 9'b111111111;
assign no[25][91] = 9'b111111111;
assign no[25][92] = 9'b111111111;
assign no[25][106] = 9'b111111111;
assign no[25][107] = 9'b111111111;
assign no[25][108] = 9'b111111111;
assign no[25][109] = 9'b111111111;
assign no[25][114] = 9'b111111111;
assign no[25][115] = 9'b111111111;
assign no[25][116] = 9'b111111111;
assign no[25][117] = 9'b111111111;
assign no[25][118] = 9'b111111111;
assign no[25][123] = 9'b111111111;
assign no[25][124] = 9'b111111111;
assign no[25][125] = 9'b111111111;
assign no[25][126] = 9'b111111111;
assign no[25][132] = 9'b111111111;
assign no[25][133] = 9'b111111111;
assign no[25][135] = 9'b111111111;
assign no[25][136] = 9'b111111111;
assign no[25][137] = 9'b111111111;
assign no[25][138] = 9'b111111111;
assign no[26][20] = 9'b111111111;
assign no[26][21] = 9'b111111111;
assign no[26][22] = 9'b111111111;
assign no[26][23] = 9'b111111111;
assign no[26][24] = 9'b111111111;
assign no[26][31] = 9'b111111111;
assign no[26][32] = 9'b111111111;
assign no[26][33] = 9'b111111111;
assign no[26][34] = 9'b111111111;
assign no[26][35] = 9'b111111111;
assign no[26][36] = 9'b111111111;
assign no[26][42] = 9'b111111111;
assign no[26][43] = 9'b111111111;
assign no[26][44] = 9'b111111111;
assign no[26][45] = 9'b111111111;
assign no[26][46] = 9'b111111111;
assign no[26][49] = 9'b111111111;
assign no[26][50] = 9'b111111111;
assign no[26][51] = 9'b111111111;
assign no[26][52] = 9'b111111111;
assign no[26][53] = 9'b111111111;
assign no[26][71] = 9'b111111111;
assign no[26][72] = 9'b111111111;
assign no[26][73] = 9'b111111111;
assign no[26][74] = 9'b111111111;
assign no[26][75] = 9'b111111111;
assign no[26][88] = 9'b111111111;
assign no[26][90] = 9'b111111111;
assign no[26][91] = 9'b111111111;
assign no[26][92] = 9'b111111111;
assign no[26][105] = 9'b111111111;
assign no[26][106] = 9'b111111111;
assign no[26][107] = 9'b111111111;
assign no[26][108] = 9'b111111111;
assign no[26][109] = 9'b111111111;
assign no[26][111] = 9'b111111111;
assign no[26][112] = 9'b111111111;
assign no[26][113] = 9'b111111111;
assign no[26][114] = 9'b111111111;
assign no[26][115] = 9'b111111111;
assign no[26][116] = 9'b111111111;
assign no[26][117] = 9'b111111111;
assign no[26][118] = 9'b111111111;
assign no[26][119] = 9'b111111111;
assign no[26][122] = 9'b111111111;
assign no[26][123] = 9'b111111111;
assign no[26][124] = 9'b111111111;
assign no[26][125] = 9'b111111111;
assign no[26][126] = 9'b111111111;
assign no[26][129] = 9'b111111111;
assign no[26][130] = 9'b111111111;
assign no[26][131] = 9'b111111111;
assign no[26][132] = 9'b111111111;
assign no[26][133] = 9'b111111111;
assign no[26][135] = 9'b111111111;
assign no[26][136] = 9'b111111111;
assign no[26][137] = 9'b111111111;
assign no[26][138] = 9'b111111111;
assign no[27][20] = 9'b111111111;
assign no[27][21] = 9'b111111111;
assign no[27][22] = 9'b111111111;
assign no[27][23] = 9'b111111111;
assign no[27][24] = 9'b111111111;
assign no[27][31] = 9'b111111111;
assign no[27][32] = 9'b111111111;
assign no[27][33] = 9'b111111111;
assign no[27][34] = 9'b111111111;
assign no[27][35] = 9'b111111111;
assign no[27][36] = 9'b111111111;
assign no[27][42] = 9'b111111111;
assign no[27][43] = 9'b111111111;
assign no[27][44] = 9'b111111111;
assign no[27][45] = 9'b111111111;
assign no[27][46] = 9'b111111111;
assign no[27][49] = 9'b111111111;
assign no[27][50] = 9'b111111111;
assign no[27][51] = 9'b111111111;
assign no[27][52] = 9'b111111111;
assign no[27][53] = 9'b111111111;
assign no[27][70] = 9'b111111111;
assign no[27][71] = 9'b111111111;
assign no[27][72] = 9'b111111111;
assign no[27][73] = 9'b111111111;
assign no[27][74] = 9'b111111111;
assign no[27][75] = 9'b111111111;
assign no[27][88] = 9'b111111111;
assign no[27][89] = 9'b111111111;
assign no[27][90] = 9'b111111111;
assign no[27][91] = 9'b111111111;
assign no[27][92] = 9'b111111111;
assign no[27][104] = 9'b111111111;
assign no[27][105] = 9'b111111111;
assign no[27][106] = 9'b111111111;
assign no[27][107] = 9'b111111111;
assign no[27][108] = 9'b111111111;
assign no[27][109] = 9'b111111111;
assign no[27][110] = 9'b111111111;
assign no[27][111] = 9'b111111111;
assign no[27][112] = 9'b111111111;
assign no[27][113] = 9'b111111111;
assign no[27][114] = 9'b111111111;
assign no[27][115] = 9'b111111111;
assign no[27][116] = 9'b111111111;
assign no[27][117] = 9'b111111111;
assign no[27][118] = 9'b111111111;
assign no[27][119] = 9'b111111111;
assign no[27][122] = 9'b111111111;
assign no[27][123] = 9'b111111111;
assign no[27][124] = 9'b111111111;
assign no[27][125] = 9'b111111111;
assign no[27][126] = 9'b111111111;
assign no[27][130] = 9'b111111111;
assign no[27][131] = 9'b111111111;
assign no[27][132] = 9'b111111111;
assign no[27][133] = 9'b111111111;
assign no[27][134] = 9'b111111111;
assign no[27][135] = 9'b111111111;
assign no[27][136] = 9'b111111111;
assign no[27][137] = 9'b111111111;
assign no[27][138] = 9'b111111111;
assign no[28][20] = 9'b111111111;
assign no[28][21] = 9'b111111111;
assign no[28][22] = 9'b111111111;
assign no[28][23] = 9'b111111111;
assign no[28][24] = 9'b111111111;
assign no[28][31] = 9'b111111111;
assign no[28][32] = 9'b111111111;
assign no[28][33] = 9'b111111111;
assign no[28][34] = 9'b111111111;
assign no[28][35] = 9'b111111111;
assign no[28][36] = 9'b111111111;
assign no[28][42] = 9'b111111111;
assign no[28][43] = 9'b111111111;
assign no[28][44] = 9'b111111111;
assign no[28][45] = 9'b111111111;
assign no[28][46] = 9'b111111111;
assign no[28][49] = 9'b111111111;
assign no[28][50] = 9'b111111111;
assign no[28][51] = 9'b111111111;
assign no[28][52] = 9'b111111111;
assign no[28][53] = 9'b111111111;
assign no[28][70] = 9'b111111111;
assign no[28][71] = 9'b111111111;
assign no[28][72] = 9'b111111111;
assign no[28][73] = 9'b111111111;
assign no[28][74] = 9'b111111111;
assign no[28][75] = 9'b111111111;
assign no[28][88] = 9'b111111111;
assign no[28][89] = 9'b111111111;
assign no[28][90] = 9'b111111111;
assign no[28][91] = 9'b111111111;
assign no[28][92] = 9'b111111111;
assign no[28][104] = 9'b111111111;
assign no[28][105] = 9'b111111111;
assign no[28][106] = 9'b111111111;
assign no[28][107] = 9'b111111111;
assign no[28][108] = 9'b111111111;
assign no[28][109] = 9'b111111111;
assign no[28][110] = 9'b111111111;
assign no[28][111] = 9'b111111111;
assign no[28][112] = 9'b111111111;
assign no[28][113] = 9'b111111111;
assign no[28][114] = 9'b111111111;
assign no[28][115] = 9'b111111111;
assign no[28][116] = 9'b111111111;
assign no[28][117] = 9'b111111111;
assign no[28][118] = 9'b111111111;
assign no[28][119] = 9'b111111111;
assign no[28][122] = 9'b111111111;
assign no[28][123] = 9'b111111111;
assign no[28][124] = 9'b111111111;
assign no[28][125] = 9'b111111111;
assign no[28][126] = 9'b111111111;
assign no[28][130] = 9'b111111111;
assign no[28][131] = 9'b111111111;
assign no[28][132] = 9'b111111111;
assign no[28][133] = 9'b111111111;
assign no[28][134] = 9'b111111111;
assign no[28][135] = 9'b111111111;
assign no[28][136] = 9'b111111111;
assign no[28][137] = 9'b111111111;
assign no[28][138] = 9'b111111111;
assign no[29][20] = 9'b111111111;
assign no[29][21] = 9'b111111111;
assign no[29][22] = 9'b111111111;
assign no[29][23] = 9'b111111111;
assign no[29][24] = 9'b111111111;
assign no[29][31] = 9'b111111111;
assign no[29][32] = 9'b111111111;
assign no[29][33] = 9'b111111111;
assign no[29][34] = 9'b111111111;
assign no[29][35] = 9'b111111111;
assign no[29][36] = 9'b111111111;
assign no[29][42] = 9'b111111111;
assign no[29][43] = 9'b111111111;
assign no[29][44] = 9'b111111111;
assign no[29][45] = 9'b111111111;
assign no[29][46] = 9'b111111111;
assign no[29][49] = 9'b111111111;
assign no[29][50] = 9'b111111111;
assign no[29][51] = 9'b111111111;
assign no[29][52] = 9'b111111111;
assign no[29][53] = 9'b111111111;
assign no[29][70] = 9'b111111111;
assign no[29][71] = 9'b111111111;
assign no[29][72] = 9'b111111111;
assign no[29][73] = 9'b111111111;
assign no[29][74] = 9'b111111111;
assign no[29][75] = 9'b111111111;
assign no[29][88] = 9'b111111111;
assign no[29][89] = 9'b111111111;
assign no[29][90] = 9'b111111111;
assign no[29][91] = 9'b111111111;
assign no[29][92] = 9'b111111111;
assign no[29][103] = 9'b111111111;
assign no[29][104] = 9'b111111111;
assign no[29][105] = 9'b111111111;
assign no[29][106] = 9'b111111111;
assign no[29][107] = 9'b111111111;
assign no[29][115] = 9'b111111111;
assign no[29][116] = 9'b111111111;
assign no[29][117] = 9'b111111111;
assign no[29][118] = 9'b111111111;
assign no[29][119] = 9'b111111111;
assign no[29][120] = 9'b111111111;
assign no[29][122] = 9'b111111111;
assign no[29][123] = 9'b111111111;
assign no[29][124] = 9'b111111111;
assign no[29][125] = 9'b111111111;
assign no[29][126] = 9'b111111111;
assign no[29][131] = 9'b111111111;
assign no[29][132] = 9'b111111111;
assign no[29][133] = 9'b111111111;
assign no[29][134] = 9'b111111111;
assign no[29][135] = 9'b111111111;
assign no[29][136] = 9'b111111111;
assign no[29][137] = 9'b111111111;
assign no[29][138] = 9'b111111111;
assign no[30][20] = 9'b111111111;
assign no[30][21] = 9'b111111111;
assign no[30][22] = 9'b111111111;
assign no[30][23] = 9'b111111111;
assign no[30][24] = 9'b111111111;
assign no[30][31] = 9'b111111111;
assign no[30][32] = 9'b111111111;
assign no[30][33] = 9'b111111111;
assign no[30][34] = 9'b111111111;
assign no[30][35] = 9'b111111111;
assign no[30][36] = 9'b111111111;
assign no[30][42] = 9'b111111111;
assign no[30][43] = 9'b111111111;
assign no[30][44] = 9'b111111111;
assign no[30][45] = 9'b111111111;
assign no[30][46] = 9'b111111111;
assign no[30][49] = 9'b111111111;
assign no[30][50] = 9'b111111111;
assign no[30][51] = 9'b111111111;
assign no[30][52] = 9'b111111111;
assign no[30][53] = 9'b111111111;
assign no[30][54] = 9'b111111111;
assign no[30][55] = 9'b111111111;
assign no[30][56] = 9'b111111111;
assign no[30][57] = 9'b111111111;
assign no[30][58] = 9'b111111111;
assign no[30][59] = 9'b111111111;
assign no[30][60] = 9'b111111111;
assign no[30][61] = 9'b111111111;
assign no[30][70] = 9'b111111111;
assign no[30][71] = 9'b111111111;
assign no[30][72] = 9'b111111111;
assign no[30][73] = 9'b111111111;
assign no[30][74] = 9'b111111111;
assign no[30][75] = 9'b111111111;
assign no[30][88] = 9'b111111111;
assign no[30][89] = 9'b111111111;
assign no[30][90] = 9'b111111111;
assign no[30][91] = 9'b111111111;
assign no[30][92] = 9'b111111111;
assign no[30][93] = 9'b111111111;
assign no[30][94] = 9'b111111111;
assign no[30][95] = 9'b111111111;
assign no[30][96] = 9'b111111111;
assign no[30][97] = 9'b111111111;
assign no[30][98] = 9'b111111111;
assign no[30][99] = 9'b111111111;
assign no[30][103] = 9'b111111111;
assign no[30][104] = 9'b111111111;
assign no[30][105] = 9'b111111111;
assign no[30][106] = 9'b111111111;
assign no[30][107] = 9'b111111111;
assign no[30][115] = 9'b111111111;
assign no[30][116] = 9'b111111111;
assign no[30][117] = 9'b111111111;
assign no[30][118] = 9'b111111111;
assign no[30][119] = 9'b111111111;
assign no[30][120] = 9'b111111111;
assign no[30][122] = 9'b111111111;
assign no[30][123] = 9'b111111111;
assign no[30][124] = 9'b111111111;
assign no[30][125] = 9'b111111111;
assign no[30][126] = 9'b111111111;
assign no[30][131] = 9'b111111111;
assign no[30][132] = 9'b111111111;
assign no[30][133] = 9'b111111111;
assign no[30][134] = 9'b111111111;
assign no[30][135] = 9'b111111111;
assign no[30][136] = 9'b111111111;
assign no[30][137] = 9'b111111111;
assign no[30][138] = 9'b111111111;
assign no[31][20] = 9'b111111111;
assign no[31][21] = 9'b111111111;
assign no[31][22] = 9'b111111111;
assign no[31][23] = 9'b111111111;
assign no[31][24] = 9'b111111111;
assign no[31][31] = 9'b111111111;
assign no[31][32] = 9'b111111111;
assign no[31][33] = 9'b111111111;
assign no[31][34] = 9'b111111111;
assign no[31][35] = 9'b111111111;
assign no[31][36] = 9'b111111111;
assign no[31][42] = 9'b111111111;
assign no[31][43] = 9'b111111111;
assign no[31][44] = 9'b111111111;
assign no[31][45] = 9'b111111111;
assign no[31][46] = 9'b111111111;
assign no[31][49] = 9'b111111111;
assign no[31][50] = 9'b111111111;
assign no[31][51] = 9'b111111111;
assign no[31][52] = 9'b111111111;
assign no[31][53] = 9'b111111111;
assign no[31][54] = 9'b111111111;
assign no[31][55] = 9'b111111111;
assign no[31][56] = 9'b111111111;
assign no[31][57] = 9'b111111111;
assign no[31][58] = 9'b111111111;
assign no[31][59] = 9'b111111111;
assign no[31][60] = 9'b111111111;
assign no[31][61] = 9'b111111111;
assign no[31][70] = 9'b111111111;
assign no[31][71] = 9'b111111111;
assign no[31][72] = 9'b111111111;
assign no[31][73] = 9'b111111111;
assign no[31][74] = 9'b111111111;
assign no[31][75] = 9'b111111111;
assign no[31][88] = 9'b111111111;
assign no[31][89] = 9'b111111111;
assign no[31][90] = 9'b111111111;
assign no[31][91] = 9'b111111111;
assign no[31][92] = 9'b111111111;
assign no[31][93] = 9'b111111111;
assign no[31][94] = 9'b111111111;
assign no[31][95] = 9'b111111111;
assign no[31][96] = 9'b111111111;
assign no[31][97] = 9'b111111111;
assign no[31][98] = 9'b111111111;
assign no[31][99] = 9'b111111111;
assign no[31][103] = 9'b111111111;
assign no[31][104] = 9'b111111111;
assign no[31][105] = 9'b111111111;
assign no[31][106] = 9'b111111111;
assign no[31][107] = 9'b111111111;
assign no[31][116] = 9'b111111111;
assign no[31][117] = 9'b111111111;
assign no[31][118] = 9'b111111111;
assign no[31][119] = 9'b111111111;
assign no[31][120] = 9'b111111111;
assign no[31][122] = 9'b111111111;
assign no[31][123] = 9'b111111111;
assign no[31][124] = 9'b111111111;
assign no[31][125] = 9'b111111111;
assign no[31][126] = 9'b111111111;
assign no[31][131] = 9'b111111111;
assign no[31][132] = 9'b111111111;
assign no[31][133] = 9'b111111111;
assign no[31][134] = 9'b111111111;
assign no[31][135] = 9'b111111111;
assign no[31][136] = 9'b111111111;
assign no[31][137] = 9'b111111111;
assign no[31][138] = 9'b111111111;
assign no[32][20] = 9'b111111111;
assign no[32][21] = 9'b111111111;
assign no[32][22] = 9'b111111111;
assign no[32][23] = 9'b111111111;
assign no[32][24] = 9'b111111111;
assign no[32][31] = 9'b111111111;
assign no[32][32] = 9'b111111111;
assign no[32][33] = 9'b111111111;
assign no[32][34] = 9'b111111111;
assign no[32][35] = 9'b111111111;
assign no[32][42] = 9'b111111111;
assign no[32][43] = 9'b111111111;
assign no[32][44] = 9'b111111111;
assign no[32][45] = 9'b111111111;
assign no[32][46] = 9'b111111111;
assign no[32][49] = 9'b111111111;
assign no[32][50] = 9'b111111111;
assign no[32][51] = 9'b111111111;
assign no[32][52] = 9'b111111111;
assign no[32][53] = 9'b111111111;
assign no[32][54] = 9'b111111111;
assign no[32][55] = 9'b111111111;
assign no[32][56] = 9'b111111111;
assign no[32][57] = 9'b111111111;
assign no[32][58] = 9'b111111111;
assign no[32][59] = 9'b111111111;
assign no[32][60] = 9'b111111111;
assign no[32][61] = 9'b111111111;
assign no[32][71] = 9'b111111111;
assign no[32][72] = 9'b111111111;
assign no[32][73] = 9'b111111111;
assign no[32][74] = 9'b111111111;
assign no[32][75] = 9'b111111111;
assign no[32][88] = 9'b111111111;
assign no[32][89] = 9'b111111111;
assign no[32][90] = 9'b111111111;
assign no[32][91] = 9'b111111111;
assign no[32][92] = 9'b111111111;
assign no[32][93] = 9'b111111111;
assign no[32][94] = 9'b111111111;
assign no[32][95] = 9'b111111111;
assign no[32][96] = 9'b111111111;
assign no[32][97] = 9'b111111111;
assign no[32][98] = 9'b111111111;
assign no[32][99] = 9'b111111111;
assign no[32][103] = 9'b111111111;
assign no[32][104] = 9'b111111111;
assign no[32][105] = 9'b111111111;
assign no[32][106] = 9'b111111111;
assign no[32][116] = 9'b111111111;
assign no[32][117] = 9'b111111111;
assign no[32][118] = 9'b111111111;
assign no[32][119] = 9'b111111111;
assign no[32][120] = 9'b111111111;
assign no[32][123] = 9'b111111111;
assign no[32][124] = 9'b111111111;
assign no[32][125] = 9'b111111111;
assign no[32][126] = 9'b111111111;
assign no[32][132] = 9'b111111111;
assign no[32][133] = 9'b111111111;
assign no[32][134] = 9'b111111111;
assign no[32][135] = 9'b111111111;
assign no[32][136] = 9'b111111111;
assign no[32][137] = 9'b111111111;
assign no[32][138] = 9'b111111111;
//Total de Lineas = 1167
endmodule

