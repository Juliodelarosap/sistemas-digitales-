`timescale 1ns / 1ps
module f1_alonzo (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (F[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= F[vcount- posy][hcount- posx][7:5];
				green <= F[vcount- posy][hcount- posx][4:2];
            blue 	<= F[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 40;
parameter RESOLUCION_Y = 60;
wire [8:0] F[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign F[0][9] = 9'b100000000;
assign F[0][10] = 9'b100000000;
assign F[0][29] = 9'b100000000;
assign F[0][30] = 9'b100000000;
assign F[1][8] = 9'b100000000;
assign F[1][9] = 9'b100100100;
assign F[1][10] = 9'b100000000;
assign F[1][11] = 9'b100000000;
assign F[1][28] = 9'b100000000;
assign F[1][29] = 9'b100000000;
assign F[1][30] = 9'b100100100;
assign F[1][31] = 9'b100000000;
assign F[2][8] = 9'b100000000;
assign F[2][9] = 9'b100101000;
assign F[2][10] = 9'b100000000;
assign F[2][11] = 9'b100000000;
assign F[2][12] = 9'b100000000;
assign F[2][13] = 9'b100000100;
assign F[2][14] = 9'b101001000;
assign F[2][15] = 9'b101000100;
assign F[2][16] = 9'b100000000;
assign F[2][17] = 9'b100000000;
assign F[2][18] = 9'b100100100;
assign F[2][19] = 9'b100100100;
assign F[2][20] = 9'b100000000;
assign F[2][21] = 9'b100000000;
assign F[2][22] = 9'b100000000;
assign F[2][23] = 9'b101000100;
assign F[2][24] = 9'b100000000;
assign F[2][25] = 9'b100100100;
assign F[2][26] = 9'b100000100;
assign F[2][27] = 9'b100000100;
assign F[2][28] = 9'b100000000;
assign F[2][29] = 9'b100000000;
assign F[2][30] = 9'b100101000;
assign F[2][31] = 9'b100000000;
assign F[3][8] = 9'b100000000;
assign F[3][9] = 9'b101011100;
assign F[3][10] = 9'b100101000;
assign F[3][11] = 9'b100000100;
assign F[3][12] = 9'b100001000;
assign F[3][13] = 9'b100101001;
assign F[3][14] = 9'b110010110;
assign F[3][15] = 9'b101110001;
assign F[3][16] = 9'b100001000;
assign F[3][17] = 9'b100001000;
assign F[3][18] = 9'b101110001;
assign F[3][19] = 9'b101001101;
assign F[3][20] = 9'b100000100;
assign F[3][21] = 9'b100001000;
assign F[3][22] = 9'b100001000;
assign F[3][23] = 9'b101110001;
assign F[3][24] = 9'b100001000;
assign F[3][25] = 9'b101110001;
assign F[3][26] = 9'b100110001;
assign F[3][27] = 9'b100010001;
assign F[3][28] = 9'b100001000;
assign F[3][29] = 9'b100101000;
assign F[3][30] = 9'b101011100;
assign F[3][31] = 9'b100000000;
assign F[4][8] = 9'b100000000;
assign F[4][9] = 9'b101011100;
assign F[4][10] = 9'b100101000;
assign F[4][11] = 9'b100000100;
assign F[4][12] = 9'b100001000;
assign F[4][13] = 9'b100001000;
assign F[4][14] = 9'b100000100;
assign F[4][15] = 9'b100000100;
assign F[4][16] = 9'b100001000;
assign F[4][17] = 9'b100000100;
assign F[4][18] = 9'b100000100;
assign F[4][19] = 9'b100000100;
assign F[4][20] = 9'b100100100;
assign F[4][21] = 9'b100100100;
assign F[4][22] = 9'b100000100;
assign F[4][23] = 9'b100000100;
assign F[4][24] = 9'b100001000;
assign F[4][25] = 9'b100000100;
assign F[4][26] = 9'b100001000;
assign F[4][27] = 9'b100010001;
assign F[4][28] = 9'b100001000;
assign F[4][29] = 9'b100101000;
assign F[4][30] = 9'b101011100;
assign F[4][31] = 9'b100000000;
assign F[5][8] = 9'b100000000;
assign F[5][9] = 9'b101111100;
assign F[5][10] = 9'b100101000;
assign F[5][11] = 9'b100000100;
assign F[5][12] = 9'b100001101;
assign F[5][13] = 9'b100001000;
assign F[5][14] = 9'b100001000;
assign F[5][15] = 9'b100001000;
assign F[5][16] = 9'b100100100;
assign F[5][17] = 9'b100100100;
assign F[5][18] = 9'b100100100;
assign F[5][19] = 9'b100100100;
assign F[5][20] = 9'b100100100;
assign F[5][21] = 9'b100100100;
assign F[5][22] = 9'b100100100;
assign F[5][23] = 9'b100100100;
assign F[5][24] = 9'b100001000;
assign F[5][25] = 9'b100001000;
assign F[5][26] = 9'b100001000;
assign F[5][27] = 9'b100001101;
assign F[5][28] = 9'b100001000;
assign F[5][29] = 9'b100101000;
assign F[5][30] = 9'b101111100;
assign F[5][31] = 9'b100000000;
assign F[6][2] = 9'b100000000;
assign F[6][3] = 9'b100000000;
assign F[6][4] = 9'b100000000;
assign F[6][5] = 9'b100000000;
assign F[6][6] = 9'b100000000;
assign F[6][8] = 9'b100000000;
assign F[6][9] = 9'b100101000;
assign F[6][10] = 9'b100000100;
assign F[6][11] = 9'b100000000;
assign F[6][12] = 9'b100000100;
assign F[6][13] = 9'b100000100;
assign F[6][14] = 9'b100000100;
assign F[6][15] = 9'b100000000;
assign F[6][16] = 9'b100000000;
assign F[6][17] = 9'b100000000;
assign F[6][18] = 9'b100000000;
assign F[6][19] = 9'b100000000;
assign F[6][20] = 9'b100000000;
assign F[6][21] = 9'b100000000;
assign F[6][22] = 9'b100000000;
assign F[6][23] = 9'b100000000;
assign F[6][24] = 9'b100000000;
assign F[6][25] = 9'b100000100;
assign F[6][26] = 9'b100000100;
assign F[6][27] = 9'b100000100;
assign F[6][28] = 9'b100000100;
assign F[6][29] = 9'b100000100;
assign F[6][30] = 9'b100101100;
assign F[6][31] = 9'b100000000;
assign F[6][33] = 9'b100000000;
assign F[6][34] = 9'b100000000;
assign F[6][35] = 9'b100000000;
assign F[6][36] = 9'b100000000;
assign F[6][37] = 9'b100000000;
assign F[7][1] = 9'b100000000;
assign F[7][2] = 9'b100000000;
assign F[7][3] = 9'b100000000;
assign F[7][4] = 9'b100000000;
assign F[7][5] = 9'b100000000;
assign F[7][6] = 9'b100000000;
assign F[7][7] = 9'b100000000;
assign F[7][10] = 9'b100000000;
assign F[7][11] = 9'b100000000;
assign F[7][12] = 9'b100100000;
assign F[7][13] = 9'b100100000;
assign F[7][14] = 9'b100100000;
assign F[7][15] = 9'b100000000;
assign F[7][16] = 9'b100000000;
assign F[7][17] = 9'b100000000;
assign F[7][18] = 9'b100000000;
assign F[7][19] = 9'b100000000;
assign F[7][20] = 9'b100000000;
assign F[7][21] = 9'b100000000;
assign F[7][22] = 9'b100000000;
assign F[7][23] = 9'b100000000;
assign F[7][24] = 9'b100000000;
assign F[7][25] = 9'b100100000;
assign F[7][26] = 9'b100100000;
assign F[7][27] = 9'b100100000;
assign F[7][28] = 9'b100000000;
assign F[7][29] = 9'b100000000;
assign F[7][32] = 9'b100000000;
assign F[7][33] = 9'b100000000;
assign F[7][34] = 9'b100000000;
assign F[7][35] = 9'b100000000;
assign F[7][36] = 9'b100000000;
assign F[7][37] = 9'b100000000;
assign F[7][38] = 9'b100000000;
assign F[8][0] = 9'b100000000;
assign F[8][1] = 9'b100000000;
assign F[8][2] = 9'b100100100;
assign F[8][3] = 9'b100100100;
assign F[8][4] = 9'b100100100;
assign F[8][5] = 9'b100100100;
assign F[8][6] = 9'b100100100;
assign F[8][7] = 9'b100000000;
assign F[8][8] = 9'b100000000;
assign F[8][12] = 9'b100000000;
assign F[8][13] = 9'b100000000;
assign F[8][14] = 9'b100000000;
assign F[8][15] = 9'b100000000;
assign F[8][16] = 9'b100000000;
assign F[8][17] = 9'b100000000;
assign F[8][18] = 9'b100000000;
assign F[8][19] = 9'b100000000;
assign F[8][20] = 9'b100000000;
assign F[8][21] = 9'b100000000;
assign F[8][22] = 9'b100000000;
assign F[8][23] = 9'b100000000;
assign F[8][24] = 9'b100000000;
assign F[8][25] = 9'b100000000;
assign F[8][26] = 9'b100000000;
assign F[8][27] = 9'b100000000;
assign F[8][31] = 9'b100000000;
assign F[8][32] = 9'b100000000;
assign F[8][33] = 9'b100100100;
assign F[8][34] = 9'b100100100;
assign F[8][35] = 9'b100100100;
assign F[8][36] = 9'b100100100;
assign F[8][37] = 9'b100100100;
assign F[8][38] = 9'b100000000;
assign F[8][39] = 9'b100000000;
assign F[9][0] = 9'b100000000;
assign F[9][1] = 9'b100000000;
assign F[9][2] = 9'b100100100;
assign F[9][3] = 9'b100000000;
assign F[9][4] = 9'b100000000;
assign F[9][5] = 9'b100000000;
assign F[9][6] = 9'b100100100;
assign F[9][7] = 9'b100000000;
assign F[9][8] = 9'b100000000;
assign F[9][9] = 9'b100000000;
assign F[9][10] = 9'b100000000;
assign F[9][11] = 9'b100000000;
assign F[9][12] = 9'b100000000;
assign F[9][13] = 9'b100000000;
assign F[9][14] = 9'b100000000;
assign F[9][15] = 9'b100000000;
assign F[9][16] = 9'b100000000;
assign F[9][17] = 9'b100000000;
assign F[9][18] = 9'b100000000;
assign F[9][19] = 9'b100000000;
assign F[9][20] = 9'b100000000;
assign F[9][21] = 9'b100000000;
assign F[9][22] = 9'b100000000;
assign F[9][23] = 9'b100000000;
assign F[9][24] = 9'b100000000;
assign F[9][25] = 9'b100000000;
assign F[9][26] = 9'b100000000;
assign F[9][27] = 9'b100000000;
assign F[9][28] = 9'b100000000;
assign F[9][29] = 9'b100000000;
assign F[9][30] = 9'b100000000;
assign F[9][31] = 9'b100000000;
assign F[9][32] = 9'b100000000;
assign F[9][33] = 9'b100100100;
assign F[9][34] = 9'b100000000;
assign F[9][35] = 9'b100000000;
assign F[9][36] = 9'b100000000;
assign F[9][37] = 9'b100100100;
assign F[9][38] = 9'b100000000;
assign F[9][39] = 9'b100000000;
assign F[10][0] = 9'b100000000;
assign F[10][1] = 9'b100000000;
assign F[10][2] = 9'b100100100;
assign F[10][3] = 9'b100000000;
assign F[10][4] = 9'b100000000;
assign F[10][5] = 9'b100000000;
assign F[10][6] = 9'b100100100;
assign F[10][7] = 9'b100000000;
assign F[10][8] = 9'b100000000;
assign F[10][9] = 9'b100000000;
assign F[10][10] = 9'b100100100;
assign F[10][11] = 9'b100000000;
assign F[10][12] = 9'b100000000;
assign F[10][13] = 9'b100000000;
assign F[10][14] = 9'b100000000;
assign F[10][15] = 9'b100000000;
assign F[10][16] = 9'b100000000;
assign F[10][17] = 9'b100000000;
assign F[10][18] = 9'b100000000;
assign F[10][19] = 9'b100000000;
assign F[10][20] = 9'b100000000;
assign F[10][21] = 9'b100000000;
assign F[10][22] = 9'b100000000;
assign F[10][23] = 9'b100000000;
assign F[10][24] = 9'b100000000;
assign F[10][25] = 9'b100000000;
assign F[10][26] = 9'b100000000;
assign F[10][27] = 9'b100000000;
assign F[10][28] = 9'b100000000;
assign F[10][29] = 9'b100100100;
assign F[10][30] = 9'b100000000;
assign F[10][31] = 9'b100000000;
assign F[10][32] = 9'b100000000;
assign F[10][33] = 9'b100100100;
assign F[10][34] = 9'b100000000;
assign F[10][35] = 9'b100000000;
assign F[10][36] = 9'b100000000;
assign F[10][37] = 9'b100100100;
assign F[10][38] = 9'b100000000;
assign F[10][39] = 9'b100000000;
assign F[11][0] = 9'b100000000;
assign F[11][1] = 9'b100000000;
assign F[11][2] = 9'b100100100;
assign F[11][3] = 9'b100000000;
assign F[11][4] = 9'b100000000;
assign F[11][5] = 9'b100000000;
assign F[11][6] = 9'b100100100;
assign F[11][7] = 9'b100000000;
assign F[11][8] = 9'b100000000;
assign F[11][9] = 9'b100000000;
assign F[11][10] = 9'b100000000;
assign F[11][11] = 9'b100100100;
assign F[11][12] = 9'b100100100;
assign F[11][13] = 9'b100000000;
assign F[11][14] = 9'b100000000;
assign F[11][15] = 9'b100000100;
assign F[11][16] = 9'b100000100;
assign F[11][17] = 9'b100000100;
assign F[11][18] = 9'b100000100;
assign F[11][19] = 9'b100000000;
assign F[11][20] = 9'b100000000;
assign F[11][21] = 9'b100000100;
assign F[11][22] = 9'b100000100;
assign F[11][23] = 9'b100000100;
assign F[11][24] = 9'b100000100;
assign F[11][25] = 9'b100000000;
assign F[11][26] = 9'b100000000;
assign F[11][27] = 9'b100100100;
assign F[11][28] = 9'b100100100;
assign F[11][29] = 9'b100000000;
assign F[11][30] = 9'b100000000;
assign F[11][31] = 9'b100000000;
assign F[11][32] = 9'b100000000;
assign F[11][33] = 9'b100100100;
assign F[11][34] = 9'b100000000;
assign F[11][35] = 9'b100000000;
assign F[11][36] = 9'b100000000;
assign F[11][37] = 9'b100100100;
assign F[11][38] = 9'b100000000;
assign F[11][39] = 9'b100000000;
assign F[12][0] = 9'b100000000;
assign F[12][1] = 9'b100000000;
assign F[12][2] = 9'b100100100;
assign F[12][3] = 9'b100100100;
assign F[12][4] = 9'b100100100;
assign F[12][5] = 9'b100100100;
assign F[12][6] = 9'b100100100;
assign F[12][7] = 9'b100000000;
assign F[12][8] = 9'b100000000;
assign F[12][11] = 9'b100000000;
assign F[12][12] = 9'b100000000;
assign F[12][13] = 9'b100100100;
assign F[12][14] = 9'b100100100;
assign F[12][15] = 9'b100000000;
assign F[12][16] = 9'b100000100;
assign F[12][17] = 9'b100000100;
assign F[12][18] = 9'b100000100;
assign F[12][19] = 9'b100000000;
assign F[12][20] = 9'b100000000;
assign F[12][21] = 9'b100000100;
assign F[12][22] = 9'b100000100;
assign F[12][23] = 9'b100000100;
assign F[12][24] = 9'b100000000;
assign F[12][25] = 9'b100100100;
assign F[12][26] = 9'b100100100;
assign F[12][27] = 9'b100000000;
assign F[12][28] = 9'b100000000;
assign F[12][31] = 9'b100000000;
assign F[12][32] = 9'b100000000;
assign F[12][33] = 9'b100100100;
assign F[12][34] = 9'b100100100;
assign F[12][35] = 9'b100100100;
assign F[12][36] = 9'b100100100;
assign F[12][37] = 9'b100100100;
assign F[12][38] = 9'b100000000;
assign F[12][39] = 9'b100000000;
assign F[13][1] = 9'b100000000;
assign F[13][2] = 9'b100000000;
assign F[13][3] = 9'b100000000;
assign F[13][4] = 9'b100000000;
assign F[13][5] = 9'b100000000;
assign F[13][6] = 9'b100000000;
assign F[13][7] = 9'b100000000;
assign F[13][9] = 9'b100000000;
assign F[13][10] = 9'b100000000;
assign F[13][11] = 9'b100100100;
assign F[13][12] = 9'b100100100;
assign F[13][13] = 9'b100000000;
assign F[13][14] = 9'b100100000;
assign F[13][15] = 9'b100000000;
assign F[13][16] = 9'b100000100;
assign F[13][17] = 9'b100000100;
assign F[13][18] = 9'b101001001;
assign F[13][19] = 9'b100100100;
assign F[13][20] = 9'b100100100;
assign F[13][21] = 9'b101001001;
assign F[13][22] = 9'b100000100;
assign F[13][23] = 9'b100000100;
assign F[13][24] = 9'b100000000;
assign F[13][25] = 9'b100100000;
assign F[13][26] = 9'b100000000;
assign F[13][27] = 9'b100100100;
assign F[13][28] = 9'b100100100;
assign F[13][29] = 9'b100000000;
assign F[13][30] = 9'b100000000;
assign F[13][32] = 9'b100000000;
assign F[13][33] = 9'b100000000;
assign F[13][34] = 9'b100000000;
assign F[13][35] = 9'b100000000;
assign F[13][36] = 9'b100000000;
assign F[13][37] = 9'b100000000;
assign F[13][38] = 9'b100000000;
assign F[14][8] = 9'b100000000;
assign F[14][9] = 9'b100000000;
assign F[14][10] = 9'b100100100;
assign F[14][11] = 9'b100100100;
assign F[14][12] = 9'b100100100;
assign F[14][13] = 9'b100100100;
assign F[14][14] = 9'b100000000;
assign F[14][15] = 9'b100000100;
assign F[14][16] = 9'b100001000;
assign F[14][17] = 9'b100001000;
assign F[14][18] = 9'b101010001;
assign F[14][19] = 9'b101110110;
assign F[14][20] = 9'b110111111;
assign F[14][21] = 9'b110011111;
assign F[14][22] = 9'b100001100;
assign F[14][23] = 9'b100001101;
assign F[14][24] = 9'b100000100;
assign F[14][25] = 9'b100000000;
assign F[14][26] = 9'b100100100;
assign F[14][27] = 9'b100100100;
assign F[14][28] = 9'b100100100;
assign F[14][29] = 9'b100100100;
assign F[14][30] = 9'b100000000;
assign F[14][31] = 9'b100000000;
assign F[15][5] = 9'b100000000;
assign F[15][6] = 9'b100000000;
assign F[15][7] = 9'b100000000;
assign F[15][8] = 9'b100100100;
assign F[15][9] = 9'b100100100;
assign F[15][10] = 9'b100100100;
assign F[15][11] = 9'b100100100;
assign F[15][12] = 9'b100100100;
assign F[15][13] = 9'b100100000;
assign F[15][14] = 9'b100000000;
assign F[15][15] = 9'b100001000;
assign F[15][16] = 9'b100001101;
assign F[15][17] = 9'b100001000;
assign F[15][18] = 9'b110111110;
assign F[15][19] = 9'b110011111;
assign F[15][20] = 9'b101110001;
assign F[15][21] = 9'b101010001;
assign F[15][22] = 9'b100010001;
assign F[15][23] = 9'b100010001;
assign F[15][24] = 9'b100010001;
assign F[15][25] = 9'b100000000;
assign F[15][26] = 9'b100100000;
assign F[15][27] = 9'b100100100;
assign F[15][28] = 9'b100100100;
assign F[15][29] = 9'b100100100;
assign F[15][30] = 9'b100100100;
assign F[15][31] = 9'b100100100;
assign F[15][32] = 9'b100000000;
assign F[15][33] = 9'b100000000;
assign F[15][34] = 9'b100000000;
assign F[16][4] = 9'b100000000;
assign F[16][5] = 9'b100000000;
assign F[16][6] = 9'b100100100;
assign F[16][7] = 9'b100100100;
assign F[16][8] = 9'b100100100;
assign F[16][9] = 9'b100100100;
assign F[16][10] = 9'b100100100;
assign F[16][11] = 9'b100100100;
assign F[16][12] = 9'b100100100;
assign F[16][13] = 9'b100100000;
assign F[16][14] = 9'b100000000;
assign F[16][15] = 9'b100001000;
assign F[16][16] = 9'b100001100;
assign F[16][17] = 9'b100001101;
assign F[16][18] = 9'b101010001;
assign F[16][19] = 9'b110011101;
assign F[16][20] = 9'b110011101;
assign F[16][21] = 9'b101010101;
assign F[16][22] = 9'b100001101;
assign F[16][23] = 9'b100001101;
assign F[16][24] = 9'b100010001;
assign F[16][25] = 9'b100000000;
assign F[16][26] = 9'b100100000;
assign F[16][27] = 9'b100100100;
assign F[16][28] = 9'b100100100;
assign F[16][29] = 9'b100100100;
assign F[16][30] = 9'b100100100;
assign F[16][31] = 9'b100100100;
assign F[16][32] = 9'b100100100;
assign F[16][33] = 9'b100100100;
assign F[16][34] = 9'b100000000;
assign F[16][35] = 9'b100000000;
assign F[17][4] = 9'b100000000;
assign F[17][5] = 9'b100000000;
assign F[17][6] = 9'b100100100;
assign F[17][7] = 9'b101001001;
assign F[17][8] = 9'b100100100;
assign F[17][9] = 9'b100100100;
assign F[17][10] = 9'b100100100;
assign F[17][11] = 9'b100100100;
assign F[17][12] = 9'b100100100;
assign F[17][13] = 9'b100100000;
assign F[17][14] = 9'b100000000;
assign F[17][15] = 9'b100001000;
assign F[17][16] = 9'b100001000;
assign F[17][17] = 9'b100001000;
assign F[17][18] = 9'b100001000;
assign F[17][19] = 9'b100111100;
assign F[17][20] = 9'b100111100;
assign F[17][21] = 9'b100001101;
assign F[17][22] = 9'b100001000;
assign F[17][23] = 9'b100001000;
assign F[17][24] = 9'b100010001;
assign F[17][25] = 9'b100000000;
assign F[17][26] = 9'b100100000;
assign F[17][27] = 9'b100100100;
assign F[17][28] = 9'b100100100;
assign F[17][29] = 9'b100100100;
assign F[17][30] = 9'b100100100;
assign F[17][31] = 9'b100100100;
assign F[17][32] = 9'b100100100;
assign F[17][33] = 9'b100100100;
assign F[17][34] = 9'b100000000;
assign F[17][35] = 9'b100000000;
assign F[18][4] = 9'b100000000;
assign F[18][5] = 9'b100100100;
assign F[18][6] = 9'b110010001;
assign F[18][7] = 9'b110010001;
assign F[18][8] = 9'b100100100;
assign F[18][9] = 9'b100100100;
assign F[18][10] = 9'b100100100;
assign F[18][11] = 9'b100100100;
assign F[18][12] = 9'b100100100;
assign F[18][13] = 9'b100000000;
assign F[18][14] = 9'b100001000;
assign F[18][15] = 9'b100001000;
assign F[18][16] = 9'b100001000;
assign F[18][17] = 9'b100000100;
assign F[18][18] = 9'b100001101;
assign F[18][19] = 9'b101011100;
assign F[18][20] = 9'b101011100;
assign F[18][21] = 9'b100001101;
assign F[18][22] = 9'b100000100;
assign F[18][23] = 9'b100001000;
assign F[18][24] = 9'b100010001;
assign F[18][25] = 9'b100001000;
assign F[18][26] = 9'b100000000;
assign F[18][27] = 9'b100100100;
assign F[18][28] = 9'b100100100;
assign F[18][29] = 9'b100100100;
assign F[18][30] = 9'b100100100;
assign F[18][31] = 9'b100100100;
assign F[18][32] = 9'b101101101;
assign F[18][33] = 9'b100100100;
assign F[18][34] = 9'b100000000;
assign F[18][35] = 9'b100000000;
assign F[19][4] = 9'b100000000;
assign F[19][5] = 9'b100100100;
assign F[19][6] = 9'b101101101;
assign F[19][7] = 9'b100100100;
assign F[19][8] = 9'b100100100;
assign F[19][9] = 9'b100100100;
assign F[19][10] = 9'b100100100;
assign F[19][11] = 9'b100100100;
assign F[19][12] = 9'b100000000;
assign F[19][13] = 9'b100000100;
assign F[19][14] = 9'b100001101;
assign F[19][15] = 9'b100001000;
assign F[19][16] = 9'b100001000;
assign F[19][17] = 9'b100000100;
assign F[19][18] = 9'b100001101;
assign F[19][19] = 9'b101011100;
assign F[19][20] = 9'b101011100;
assign F[19][21] = 9'b100001101;
assign F[19][22] = 9'b100000100;
assign F[19][23] = 9'b100001000;
assign F[19][24] = 9'b100001000;
assign F[19][25] = 9'b100010001;
assign F[19][26] = 9'b100000100;
assign F[19][27] = 9'b100000000;
assign F[19][28] = 9'b100100100;
assign F[19][29] = 9'b100100100;
assign F[19][30] = 9'b100100100;
assign F[19][31] = 9'b100100100;
assign F[19][32] = 9'b110010001;
assign F[19][33] = 9'b110110110;
assign F[19][34] = 9'b100100100;
assign F[19][35] = 9'b100000000;
assign F[20][4] = 9'b100000000;
assign F[20][5] = 9'b100000000;
assign F[20][6] = 9'b100100100;
assign F[20][7] = 9'b110010010;
assign F[20][8] = 9'b100100100;
assign F[20][9] = 9'b100100100;
assign F[20][10] = 9'b100100100;
assign F[20][11] = 9'b100000000;
assign F[20][12] = 9'b100000100;
assign F[20][13] = 9'b100001101;
assign F[20][14] = 9'b100001000;
assign F[20][15] = 9'b100001000;
assign F[20][16] = 9'b100001000;
assign F[20][17] = 9'b100101101;
assign F[20][18] = 9'b100001101;
assign F[20][19] = 9'b100110100;
assign F[20][20] = 9'b100110100;
assign F[20][21] = 9'b100001101;
assign F[20][22] = 9'b100101101;
assign F[20][23] = 9'b100001000;
assign F[20][24] = 9'b100001000;
assign F[20][25] = 9'b100001101;
assign F[20][26] = 9'b100010001;
assign F[20][27] = 9'b100000100;
assign F[20][28] = 9'b100000000;
assign F[20][29] = 9'b100100100;
assign F[20][30] = 9'b100100100;
assign F[20][31] = 9'b100100100;
assign F[20][32] = 9'b110010001;
assign F[20][33] = 9'b101001001;
assign F[20][34] = 9'b100000000;
assign F[20][35] = 9'b100000000;
assign F[21][4] = 9'b100000000;
assign F[21][5] = 9'b100000000;
assign F[21][6] = 9'b100100100;
assign F[21][7] = 9'b100100100;
assign F[21][8] = 9'b100100100;
assign F[21][9] = 9'b100100100;
assign F[21][10] = 9'b100000000;
assign F[21][11] = 9'b100000100;
assign F[21][12] = 9'b100001000;
assign F[21][13] = 9'b100001000;
assign F[21][14] = 9'b100001000;
assign F[21][15] = 9'b100001000;
assign F[21][16] = 9'b100001000;
assign F[21][17] = 9'b111111111;
assign F[21][18] = 9'b101010001;
assign F[21][19] = 9'b100001000;
assign F[21][20] = 9'b100001000;
assign F[21][21] = 9'b101011110;
assign F[21][22] = 9'b111111111;
assign F[21][23] = 9'b100001000;
assign F[21][24] = 9'b100001000;
assign F[21][25] = 9'b100000100;
assign F[21][26] = 9'b100001101;
assign F[21][27] = 9'b100001100;
assign F[21][28] = 9'b100000100;
assign F[21][29] = 9'b100000000;
assign F[21][30] = 9'b100100100;
assign F[21][31] = 9'b100100100;
assign F[21][32] = 9'b110010001;
assign F[21][33] = 9'b101001000;
assign F[21][34] = 9'b100000000;
assign F[21][35] = 9'b100000000;
assign F[22][4] = 9'b100000000;
assign F[22][5] = 9'b100000000;
assign F[22][6] = 9'b100100100;
assign F[22][7] = 9'b100100100;
assign F[22][8] = 9'b100100100;
assign F[22][9] = 9'b100100100;
assign F[22][10] = 9'b100000000;
assign F[22][11] = 9'b100001000;
assign F[22][12] = 9'b100001101;
assign F[22][13] = 9'b100001000;
assign F[22][14] = 9'b100000100;
assign F[22][15] = 9'b100001000;
assign F[22][16] = 9'b111111111;
assign F[22][17] = 9'b101010001;
assign F[22][18] = 9'b100001101;
assign F[22][19] = 9'b100001000;
assign F[22][20] = 9'b100001000;
assign F[22][21] = 9'b100001101;
assign F[22][22] = 9'b101010001;
assign F[22][23] = 9'b111111111;
assign F[22][24] = 9'b100001000;
assign F[22][25] = 9'b100000100;
assign F[22][26] = 9'b100000100;
assign F[22][27] = 9'b100001101;
assign F[22][28] = 9'b100001000;
assign F[22][29] = 9'b100000000;
assign F[22][30] = 9'b100100100;
assign F[22][31] = 9'b100100100;
assign F[22][32] = 9'b101001001;
assign F[22][33] = 9'b100100100;
assign F[22][34] = 9'b100000000;
assign F[22][35] = 9'b100000000;
assign F[23][4] = 9'b100000000;
assign F[23][5] = 9'b100000000;
assign F[23][6] = 9'b100100100;
assign F[23][7] = 9'b100100100;
assign F[23][8] = 9'b100100100;
assign F[23][9] = 9'b100000000;
assign F[23][10] = 9'b100001000;
assign F[23][11] = 9'b100001101;
assign F[23][12] = 9'b100001000;
assign F[23][13] = 9'b100000100;
assign F[23][14] = 9'b100001000;
assign F[23][15] = 9'b100101000;
assign F[23][16] = 9'b110011110;
assign F[23][17] = 9'b100001101;
assign F[23][18] = 9'b100001000;
assign F[23][19] = 9'b100001000;
assign F[23][20] = 9'b100001000;
assign F[23][21] = 9'b100001000;
assign F[23][22] = 9'b100001101;
assign F[23][23] = 9'b110011110;
assign F[23][24] = 9'b100101000;
assign F[23][25] = 9'b100001000;
assign F[23][26] = 9'b100000100;
assign F[23][27] = 9'b100001000;
assign F[23][28] = 9'b100001101;
assign F[23][29] = 9'b100001000;
assign F[23][30] = 9'b100000000;
assign F[23][31] = 9'b100100100;
assign F[23][32] = 9'b100100100;
assign F[23][33] = 9'b100100100;
assign F[23][34] = 9'b100000000;
assign F[23][35] = 9'b100000000;
assign F[24][4] = 9'b100000000;
assign F[24][5] = 9'b100000000;
assign F[24][6] = 9'b100100100;
assign F[24][7] = 9'b100100100;
assign F[24][8] = 9'b100000000;
assign F[24][9] = 9'b100001000;
assign F[24][10] = 9'b100001000;
assign F[24][11] = 9'b100001000;
assign F[24][12] = 9'b100000100;
assign F[24][13] = 9'b100000100;
assign F[24][14] = 9'b100000100;
assign F[24][15] = 9'b100001000;
assign F[24][16] = 9'b100001101;
assign F[24][17] = 9'b100001100;
assign F[24][18] = 9'b100001000;
assign F[24][19] = 9'b100001000;
assign F[24][20] = 9'b100001000;
assign F[24][21] = 9'b100001000;
assign F[24][22] = 9'b100001100;
assign F[24][23] = 9'b100001101;
assign F[24][24] = 9'b100001000;
assign F[24][25] = 9'b100000100;
assign F[24][26] = 9'b100000100;
assign F[24][27] = 9'b100000100;
assign F[24][28] = 9'b100001000;
assign F[24][29] = 9'b100001000;
assign F[24][30] = 9'b100000100;
assign F[24][31] = 9'b100000000;
assign F[24][32] = 9'b100100100;
assign F[24][33] = 9'b100100100;
assign F[24][34] = 9'b100000000;
assign F[24][35] = 9'b100000000;
assign F[25][4] = 9'b100000000;
assign F[25][5] = 9'b100000000;
assign F[25][6] = 9'b100100100;
assign F[25][7] = 9'b100100100;
assign F[25][8] = 9'b100000000;
assign F[25][9] = 9'b100001000;
assign F[25][10] = 9'b100001000;
assign F[25][11] = 9'b100000100;
assign F[25][12] = 9'b100000100;
assign F[25][13] = 9'b100001000;
assign F[25][14] = 9'b100001000;
assign F[25][15] = 9'b100001000;
assign F[25][16] = 9'b100001101;
assign F[25][17] = 9'b100001101;
assign F[25][18] = 9'b100001000;
assign F[25][19] = 9'b100001000;
assign F[25][20] = 9'b100001000;
assign F[25][21] = 9'b100001000;
assign F[25][22] = 9'b100001101;
assign F[25][23] = 9'b100010001;
assign F[25][24] = 9'b100001000;
assign F[25][25] = 9'b100001000;
assign F[25][26] = 9'b100001000;
assign F[25][27] = 9'b100000100;
assign F[25][28] = 9'b100000100;
assign F[25][29] = 9'b100001000;
assign F[25][30] = 9'b100001000;
assign F[25][31] = 9'b100000000;
assign F[25][32] = 9'b100100100;
assign F[25][33] = 9'b100100100;
assign F[25][34] = 9'b100000000;
assign F[25][35] = 9'b100000000;
assign F[26][4] = 9'b100000000;
assign F[26][5] = 9'b100000000;
assign F[26][6] = 9'b100100100;
assign F[26][7] = 9'b100100100;
assign F[26][8] = 9'b100000000;
assign F[26][9] = 9'b100001000;
assign F[26][10] = 9'b100001000;
assign F[26][11] = 9'b100000100;
assign F[26][12] = 9'b100001000;
assign F[26][13] = 9'b100000100;
assign F[26][14] = 9'b100001000;
assign F[26][15] = 9'b100001000;
assign F[26][16] = 9'b100000100;
assign F[26][17] = 9'b100000100;
assign F[26][18] = 9'b100001000;
assign F[26][19] = 9'b100001000;
assign F[26][20] = 9'b100001000;
assign F[26][21] = 9'b100001000;
assign F[26][22] = 9'b100000100;
assign F[26][23] = 9'b100000100;
assign F[26][24] = 9'b100001101;
assign F[26][25] = 9'b100001000;
assign F[26][26] = 9'b100000100;
assign F[26][27] = 9'b100001000;
assign F[26][28] = 9'b100000100;
assign F[26][29] = 9'b100001000;
assign F[26][30] = 9'b100001000;
assign F[26][31] = 9'b100000000;
assign F[26][32] = 9'b100100100;
assign F[26][33] = 9'b100100100;
assign F[26][34] = 9'b100000000;
assign F[26][35] = 9'b100000000;
assign F[27][4] = 9'b100000000;
assign F[27][5] = 9'b100000000;
assign F[27][6] = 9'b100100100;
assign F[27][7] = 9'b100100100;
assign F[27][8] = 9'b100000000;
assign F[27][9] = 9'b100001000;
assign F[27][10] = 9'b100001000;
assign F[27][11] = 9'b100000100;
assign F[27][12] = 9'b100000100;
assign F[27][13] = 9'b100001000;
assign F[27][14] = 9'b100001000;
assign F[27][15] = 9'b100001000;
assign F[27][16] = 9'b100000000;
assign F[27][17] = 9'b100100000;
assign F[27][18] = 9'b100000000;
assign F[27][19] = 9'b100000000;
assign F[27][20] = 9'b100000000;
assign F[27][21] = 9'b100000000;
assign F[27][22] = 9'b100100000;
assign F[27][23] = 9'b100000000;
assign F[27][24] = 9'b100010001;
assign F[27][25] = 9'b100001000;
assign F[27][26] = 9'b100001000;
assign F[27][27] = 9'b100000100;
assign F[27][28] = 9'b100000100;
assign F[27][29] = 9'b100001000;
assign F[27][30] = 9'b100001000;
assign F[27][31] = 9'b100000000;
assign F[27][32] = 9'b100100100;
assign F[27][33] = 9'b100100100;
assign F[27][34] = 9'b100000000;
assign F[27][35] = 9'b100000000;
assign F[28][4] = 9'b100000000;
assign F[28][5] = 9'b100000000;
assign F[28][6] = 9'b100100100;
assign F[28][7] = 9'b100100100;
assign F[28][8] = 9'b100000000;
assign F[28][9] = 9'b100000100;
assign F[28][10] = 9'b100001000;
assign F[28][11] = 9'b100001000;
assign F[28][12] = 9'b100001000;
assign F[28][13] = 9'b100001000;
assign F[28][14] = 9'b100001000;
assign F[28][15] = 9'b100010001;
assign F[28][16] = 9'b100000000;
assign F[28][17] = 9'b100000000;
assign F[28][18] = 9'b100000000;
assign F[28][19] = 9'b100000000;
assign F[28][20] = 9'b100000000;
assign F[28][21] = 9'b100000000;
assign F[28][22] = 9'b100000000;
assign F[28][23] = 9'b100000000;
assign F[28][24] = 9'b100001101;
assign F[28][25] = 9'b100001101;
assign F[28][26] = 9'b100001000;
assign F[28][27] = 9'b100001000;
assign F[28][28] = 9'b100001000;
assign F[28][29] = 9'b100001000;
assign F[28][30] = 9'b100000100;
assign F[28][31] = 9'b100000000;
assign F[28][32] = 9'b100100100;
assign F[28][33] = 9'b100100100;
assign F[28][34] = 9'b100000000;
assign F[28][35] = 9'b100000000;
assign F[29][4] = 9'b100000000;
assign F[29][5] = 9'b100000000;
assign F[29][6] = 9'b100100100;
assign F[29][7] = 9'b100000000;
assign F[29][8] = 9'b100001000;
assign F[29][9] = 9'b100001000;
assign F[29][10] = 9'b100001000;
assign F[29][11] = 9'b100001000;
assign F[29][12] = 9'b100001000;
assign F[29][13] = 9'b100001000;
assign F[29][14] = 9'b100001101;
assign F[29][15] = 9'b100001101;
assign F[29][16] = 9'b100001000;
assign F[29][17] = 9'b100000000;
assign F[29][18] = 9'b100000000;
assign F[29][19] = 9'b100000000;
assign F[29][20] = 9'b100000000;
assign F[29][21] = 9'b100000000;
assign F[29][22] = 9'b100000000;
assign F[29][23] = 9'b100001000;
assign F[29][24] = 9'b100001101;
assign F[29][25] = 9'b100010001;
assign F[29][26] = 9'b100001000;
assign F[29][27] = 9'b100001000;
assign F[29][28] = 9'b100001000;
assign F[29][29] = 9'b100001000;
assign F[29][30] = 9'b100001000;
assign F[29][31] = 9'b100001000;
assign F[29][32] = 9'b100000000;
assign F[29][33] = 9'b100100100;
assign F[29][34] = 9'b100000000;
assign F[29][35] = 9'b100000000;
assign F[30][4] = 9'b100000000;
assign F[30][5] = 9'b100000000;
assign F[30][6] = 9'b100100100;
assign F[30][7] = 9'b100000000;
assign F[30][8] = 9'b100001000;
assign F[30][9] = 9'b100001000;
assign F[30][10] = 9'b100001000;
assign F[30][11] = 9'b100001000;
assign F[30][12] = 9'b100001000;
assign F[30][13] = 9'b100001000;
assign F[30][14] = 9'b100010001;
assign F[30][15] = 9'b100001000;
assign F[30][16] = 9'b100001000;
assign F[30][17] = 9'b100000000;
assign F[30][18] = 9'b100000000;
assign F[30][19] = 9'b100100100;
assign F[30][20] = 9'b100100100;
assign F[30][21] = 9'b100000000;
assign F[30][22] = 9'b100000000;
assign F[30][23] = 9'b100001000;
assign F[30][24] = 9'b100001000;
assign F[30][25] = 9'b100010001;
assign F[30][26] = 9'b100001000;
assign F[30][27] = 9'b100000100;
assign F[30][28] = 9'b100001000;
assign F[30][29] = 9'b100001000;
assign F[30][30] = 9'b100001000;
assign F[30][31] = 9'b100001000;
assign F[30][32] = 9'b100000000;
assign F[30][33] = 9'b100100100;
assign F[30][34] = 9'b100000000;
assign F[30][35] = 9'b100000000;
assign F[31][4] = 9'b100000000;
assign F[31][5] = 9'b100000000;
assign F[31][6] = 9'b100100100;
assign F[31][7] = 9'b100000000;
assign F[31][8] = 9'b100001000;
assign F[31][9] = 9'b100001000;
assign F[31][10] = 9'b100001000;
assign F[31][11] = 9'b100001000;
assign F[31][12] = 9'b100001000;
assign F[31][13] = 9'b100001101;
assign F[31][14] = 9'b100010001;
assign F[31][15] = 9'b100001000;
assign F[31][16] = 9'b100001000;
assign F[31][17] = 9'b100000000;
assign F[31][18] = 9'b100000000;
assign F[31][19] = 9'b100100100;
assign F[31][20] = 9'b100100100;
assign F[31][21] = 9'b100000000;
assign F[31][22] = 9'b100000000;
assign F[31][23] = 9'b100001000;
assign F[31][24] = 9'b100001000;
assign F[31][25] = 9'b100010001;
assign F[31][26] = 9'b100001101;
assign F[31][27] = 9'b100001000;
assign F[31][28] = 9'b100001000;
assign F[31][29] = 9'b100001000;
assign F[31][30] = 9'b100001000;
assign F[31][31] = 9'b100001000;
assign F[31][32] = 9'b100000000;
assign F[31][33] = 9'b100100100;
assign F[31][34] = 9'b100000000;
assign F[31][35] = 9'b100000000;
assign F[32][4] = 9'b100000000;
assign F[32][5] = 9'b100000000;
assign F[32][6] = 9'b100100000;
assign F[32][7] = 9'b100000000;
assign F[32][8] = 9'b100001000;
assign F[32][9] = 9'b100001101;
assign F[32][10] = 9'b100001000;
assign F[32][11] = 9'b100001000;
assign F[32][12] = 9'b100000100;
assign F[32][13] = 9'b100000100;
assign F[32][14] = 9'b100001101;
assign F[32][15] = 9'b100001000;
assign F[32][16] = 9'b100000000;
assign F[32][17] = 9'b100000000;
assign F[32][18] = 9'b100100100;
assign F[32][19] = 9'b100100100;
assign F[32][20] = 9'b100100100;
assign F[32][21] = 9'b100100100;
assign F[32][22] = 9'b100000000;
assign F[32][23] = 9'b100000000;
assign F[32][24] = 9'b100001000;
assign F[32][25] = 9'b100001101;
assign F[32][26] = 9'b100000100;
assign F[32][27] = 9'b100000100;
assign F[32][28] = 9'b100001000;
assign F[32][29] = 9'b100001000;
assign F[32][30] = 9'b100001000;
assign F[32][31] = 9'b100001000;
assign F[32][32] = 9'b100000000;
assign F[32][33] = 9'b100100000;
assign F[32][34] = 9'b100000000;
assign F[32][35] = 9'b100000000;
assign F[33][4] = 9'b100000000;
assign F[33][5] = 9'b100000100;
assign F[33][6] = 9'b100000000;
assign F[33][7] = 9'b100000000;
assign F[33][8] = 9'b100000000;
assign F[33][9] = 9'b100000100;
assign F[33][10] = 9'b100000100;
assign F[33][11] = 9'b100000100;
assign F[33][12] = 9'b100000000;
assign F[33][13] = 9'b100000000;
assign F[33][14] = 9'b100001000;
assign F[33][15] = 9'b100000000;
assign F[33][16] = 9'b100000100;
assign F[33][17] = 9'b100000000;
assign F[33][18] = 9'b100000000;
assign F[33][19] = 9'b100100100;
assign F[33][20] = 9'b100100100;
assign F[33][21] = 9'b100000000;
assign F[33][22] = 9'b100000000;
assign F[33][23] = 9'b100000100;
assign F[33][24] = 9'b100000000;
assign F[33][25] = 9'b100001000;
assign F[33][26] = 9'b100000000;
assign F[33][27] = 9'b100000000;
assign F[33][28] = 9'b100000100;
assign F[33][29] = 9'b100000100;
assign F[33][30] = 9'b100000000;
assign F[33][31] = 9'b100000000;
assign F[33][32] = 9'b100000000;
assign F[33][33] = 9'b100000000;
assign F[33][34] = 9'b100000100;
assign F[33][35] = 9'b100000100;
assign F[34][3] = 9'b100000000;
assign F[34][4] = 9'b100000100;
assign F[34][5] = 9'b100001000;
assign F[34][6] = 9'b100001000;
assign F[34][7] = 9'b100001000;
assign F[34][8] = 9'b100001000;
assign F[34][9] = 9'b100001000;
assign F[34][10] = 9'b100000100;
assign F[34][11] = 9'b100000100;
assign F[34][12] = 9'b100000000;
assign F[34][13] = 9'b100000000;
assign F[34][14] = 9'b100001000;
assign F[34][15] = 9'b100000000;
assign F[34][16] = 9'b100000100;
assign F[34][17] = 9'b100000100;
assign F[34][18] = 9'b100000000;
assign F[34][19] = 9'b100000000;
assign F[34][20] = 9'b100000000;
assign F[34][21] = 9'b100000000;
assign F[34][22] = 9'b100000100;
assign F[34][23] = 9'b100000100;
assign F[34][24] = 9'b100000000;
assign F[34][25] = 9'b100001000;
assign F[34][26] = 9'b100000000;
assign F[34][27] = 9'b100000000;
assign F[34][28] = 9'b100000100;
assign F[34][29] = 9'b100000100;
assign F[34][30] = 9'b100001000;
assign F[34][31] = 9'b100001000;
assign F[34][32] = 9'b100001000;
assign F[34][33] = 9'b100001101;
assign F[34][34] = 9'b100010001;
assign F[34][35] = 9'b100000100;
assign F[34][36] = 9'b100000000;
assign F[35][4] = 9'b100000000;
assign F[35][5] = 9'b100000000;
assign F[35][6] = 9'b100000000;
assign F[35][7] = 9'b100000100;
assign F[35][8] = 9'b100000100;
assign F[35][9] = 9'b100000100;
assign F[35][10] = 9'b100000100;
assign F[35][11] = 9'b100001000;
assign F[35][12] = 9'b100000100;
assign F[35][13] = 9'b100000100;
assign F[35][14] = 9'b100000100;
assign F[35][15] = 9'b100000000;
assign F[35][16] = 9'b100000000;
assign F[35][17] = 9'b100000100;
assign F[35][18] = 9'b100001000;
assign F[35][19] = 9'b100000100;
assign F[35][20] = 9'b100000100;
assign F[35][21] = 9'b100001000;
assign F[35][22] = 9'b100000100;
assign F[35][23] = 9'b100000000;
assign F[35][24] = 9'b100000000;
assign F[35][25] = 9'b100000100;
assign F[35][26] = 9'b100000100;
assign F[35][27] = 9'b100000100;
assign F[35][28] = 9'b100001000;
assign F[35][29] = 9'b100000100;
assign F[35][30] = 9'b100001000;
assign F[35][31] = 9'b100001000;
assign F[35][32] = 9'b100001000;
assign F[35][33] = 9'b100000100;
assign F[35][34] = 9'b100000000;
assign F[35][35] = 9'b100000000;
assign F[36][4] = 9'b100000000;
assign F[36][5] = 9'b100000000;
assign F[36][6] = 9'b100100100;
assign F[36][7] = 9'b100000000;
assign F[36][8] = 9'b100000000;
assign F[36][9] = 9'b100000100;
assign F[36][10] = 9'b100000100;
assign F[36][11] = 9'b100000100;
assign F[36][12] = 9'b100000100;
assign F[36][13] = 9'b100000000;
assign F[36][14] = 9'b100000000;
assign F[36][15] = 9'b100000000;
assign F[36][16] = 9'b100100100;
assign F[36][17] = 9'b100000000;
assign F[36][18] = 9'b100000000;
assign F[36][19] = 9'b100101100;
assign F[36][20] = 9'b100101100;
assign F[36][21] = 9'b100000000;
assign F[36][22] = 9'b100000000;
assign F[36][23] = 9'b100100100;
assign F[36][24] = 9'b100000000;
assign F[36][25] = 9'b100000000;
assign F[36][26] = 9'b100000000;
assign F[36][27] = 9'b100000100;
assign F[36][28] = 9'b100000100;
assign F[36][29] = 9'b100000100;
assign F[36][30] = 9'b100001000;
assign F[36][31] = 9'b100000000;
assign F[36][32] = 9'b100000000;
assign F[36][33] = 9'b100100100;
assign F[36][34] = 9'b100000000;
assign F[36][35] = 9'b100000000;
assign F[37][4] = 9'b100000000;
assign F[37][5] = 9'b100000000;
assign F[37][6] = 9'b100100100;
assign F[37][7] = 9'b100100100;
assign F[37][8] = 9'b100000000;
assign F[37][9] = 9'b100001000;
assign F[37][10] = 9'b100001000;
assign F[37][11] = 9'b100000100;
assign F[37][12] = 9'b100000100;
assign F[37][13] = 9'b100000000;
assign F[37][14] = 9'b100000000;
assign F[37][15] = 9'b100000000;
assign F[37][16] = 9'b100100000;
assign F[37][17] = 9'b100100100;
assign F[37][18] = 9'b100000000;
assign F[37][19] = 9'b100001000;
assign F[37][20] = 9'b100001000;
assign F[37][21] = 9'b100000000;
assign F[37][22] = 9'b100100100;
assign F[37][23] = 9'b100100000;
assign F[37][24] = 9'b100000000;
assign F[37][25] = 9'b100000000;
assign F[37][26] = 9'b100000000;
assign F[37][27] = 9'b100000100;
assign F[37][28] = 9'b100000100;
assign F[37][29] = 9'b100001101;
assign F[37][30] = 9'b100001100;
assign F[37][31] = 9'b100000000;
assign F[37][32] = 9'b100100100;
assign F[37][33] = 9'b100100100;
assign F[37][34] = 9'b100000000;
assign F[37][35] = 9'b100000000;
assign F[38][5] = 9'b100000000;
assign F[38][6] = 9'b100100100;
assign F[38][7] = 9'b100100100;
assign F[38][8] = 9'b100100100;
assign F[38][9] = 9'b100000000;
assign F[38][10] = 9'b100000000;
assign F[38][11] = 9'b100000000;
assign F[38][12] = 9'b100000000;
assign F[38][13] = 9'b100000000;
assign F[38][14] = 9'b100000000;
assign F[38][15] = 9'b100001000;
assign F[38][16] = 9'b100000100;
assign F[38][17] = 9'b100000000;
assign F[38][18] = 9'b100000000;
assign F[38][19] = 9'b100000100;
assign F[38][20] = 9'b100000100;
assign F[38][21] = 9'b100000000;
assign F[38][22] = 9'b100000000;
assign F[38][23] = 9'b100000100;
assign F[38][24] = 9'b100010001;
assign F[38][25] = 9'b100000000;
assign F[38][26] = 9'b100000000;
assign F[38][27] = 9'b100000000;
assign F[38][28] = 9'b100000000;
assign F[38][29] = 9'b100000000;
assign F[38][30] = 9'b100000000;
assign F[38][31] = 9'b100100100;
assign F[38][32] = 9'b100100100;
assign F[38][33] = 9'b100100100;
assign F[38][34] = 9'b100000000;
assign F[39][6] = 9'b100000000;
assign F[39][7] = 9'b100000000;
assign F[39][8] = 9'b100000000;
assign F[39][9] = 9'b100000000;
assign F[39][10] = 9'b100000000;
assign F[39][11] = 9'b100000000;
assign F[39][12] = 9'b100000000;
assign F[39][13] = 9'b100000000;
assign F[39][14] = 9'b100000000;
assign F[39][15] = 9'b100001000;
assign F[39][16] = 9'b100001000;
assign F[39][17] = 9'b100000100;
assign F[39][18] = 9'b100000000;
assign F[39][19] = 9'b100000000;
assign F[39][20] = 9'b100000000;
assign F[39][21] = 9'b100000000;
assign F[39][22] = 9'b100000100;
assign F[39][23] = 9'b100001000;
assign F[39][24] = 9'b100010001;
assign F[39][25] = 9'b100000000;
assign F[39][26] = 9'b100000000;
assign F[39][27] = 9'b100000000;
assign F[39][28] = 9'b100000000;
assign F[39][29] = 9'b100000000;
assign F[39][30] = 9'b100000000;
assign F[39][31] = 9'b100000000;
assign F[39][32] = 9'b100000000;
assign F[39][33] = 9'b100000000;
assign F[40][13] = 9'b100000000;
assign F[40][14] = 9'b100000000;
assign F[40][15] = 9'b100001000;
assign F[40][16] = 9'b100001000;
assign F[40][17] = 9'b100001000;
assign F[40][18] = 9'b100000100;
assign F[40][19] = 9'b100000100;
assign F[40][20] = 9'b100000100;
assign F[40][21] = 9'b100000100;
assign F[40][22] = 9'b100001000;
assign F[40][23] = 9'b110001000;
assign F[40][24] = 9'b100010001;
assign F[40][25] = 9'b100000000;
assign F[40][26] = 9'b100000000;
assign F[41][14] = 9'b100000000;
assign F[41][15] = 9'b100000100;
assign F[41][16] = 9'b100001000;
assign F[41][17] = 9'b100001000;
assign F[41][18] = 9'b101010001;
assign F[41][19] = 9'b110010110;
assign F[41][20] = 9'b110010110;
assign F[41][21] = 9'b101010001;
assign F[41][22] = 9'b100001000;
assign F[41][23] = 9'b100010001;
assign F[41][24] = 9'b100001000;
assign F[41][25] = 9'b100000000;
assign F[42][15] = 9'b100000000;
assign F[42][16] = 9'b100001000;
assign F[42][17] = 9'b100001000;
assign F[42][18] = 9'b100101001;
assign F[42][19] = 9'b100101101;
assign F[42][20] = 9'b100101101;
assign F[42][21] = 9'b100101001;
assign F[42][22] = 9'b100001000;
assign F[42][23] = 9'b100001101;
assign F[42][24] = 9'b100000000;
assign F[43][1] = 9'b100000000;
assign F[43][2] = 9'b100000000;
assign F[43][3] = 9'b100000000;
assign F[43][4] = 9'b100000000;
assign F[43][5] = 9'b100000000;
assign F[43][6] = 9'b100000000;
assign F[43][7] = 9'b100000000;
assign F[43][12] = 9'b100000000;
assign F[43][13] = 9'b100000000;
assign F[43][14] = 9'b100000000;
assign F[43][15] = 9'b100000000;
assign F[43][16] = 9'b100001000;
assign F[43][17] = 9'b100001000;
assign F[43][18] = 9'b100000100;
assign F[43][19] = 9'b100000100;
assign F[43][20] = 9'b100000100;
assign F[43][21] = 9'b100000100;
assign F[43][22] = 9'b100001000;
assign F[43][23] = 9'b100001101;
assign F[43][24] = 9'b100000000;
assign F[43][25] = 9'b100000000;
assign F[43][26] = 9'b100000000;
assign F[43][27] = 9'b100000000;
assign F[43][32] = 9'b100000000;
assign F[43][33] = 9'b100000000;
assign F[43][34] = 9'b100000000;
assign F[43][35] = 9'b100000000;
assign F[43][36] = 9'b100000000;
assign F[43][37] = 9'b100000000;
assign F[43][38] = 9'b100000000;
assign F[44][0] = 9'b100000000;
assign F[44][1] = 9'b100000000;
assign F[44][2] = 9'b100100100;
assign F[44][3] = 9'b100100100;
assign F[44][4] = 9'b100100100;
assign F[44][5] = 9'b100100100;
assign F[44][6] = 9'b100100100;
assign F[44][7] = 9'b100000000;
assign F[44][8] = 9'b100000000;
assign F[44][10] = 9'b100000000;
assign F[44][11] = 9'b100000000;
assign F[44][12] = 9'b100100100;
assign F[44][13] = 9'b100000000;
assign F[44][14] = 9'b100000000;
assign F[44][15] = 9'b100000000;
assign F[44][16] = 9'b100001000;
assign F[44][17] = 9'b100001000;
assign F[44][18] = 9'b110010110;
assign F[44][19] = 9'b101001101;
assign F[44][20] = 9'b101001101;
assign F[44][21] = 9'b110010110;
assign F[44][22] = 9'b100001000;
assign F[44][23] = 9'b100001101;
assign F[44][24] = 9'b100000000;
assign F[44][25] = 9'b100000000;
assign F[44][26] = 9'b100000000;
assign F[44][27] = 9'b100100100;
assign F[44][28] = 9'b100000000;
assign F[44][29] = 9'b100000000;
assign F[44][31] = 9'b100000000;
assign F[44][32] = 9'b100000000;
assign F[44][33] = 9'b100100100;
assign F[44][34] = 9'b100100100;
assign F[44][35] = 9'b100100100;
assign F[44][36] = 9'b100100100;
assign F[44][37] = 9'b100100100;
assign F[44][38] = 9'b100000000;
assign F[44][39] = 9'b100000000;
assign F[45][0] = 9'b100000000;
assign F[45][1] = 9'b100000000;
assign F[45][2] = 9'b100100100;
assign F[45][3] = 9'b100000000;
assign F[45][4] = 9'b100000000;
assign F[45][5] = 9'b100000000;
assign F[45][6] = 9'b100100100;
assign F[45][7] = 9'b100000000;
assign F[45][8] = 9'b100000000;
assign F[45][9] = 9'b100000000;
assign F[45][10] = 9'b100000000;
assign F[45][11] = 9'b100100100;
assign F[45][12] = 9'b100000000;
assign F[45][13] = 9'b100000000;
assign F[45][14] = 9'b100000000;
assign F[45][15] = 9'b100000000;
assign F[45][16] = 9'b100001000;
assign F[45][17] = 9'b100001000;
assign F[45][18] = 9'b101110001;
assign F[45][19] = 9'b100101101;
assign F[45][20] = 9'b100101101;
assign F[45][21] = 9'b110010010;
assign F[45][22] = 9'b100001000;
assign F[45][23] = 9'b100001101;
assign F[45][24] = 9'b100000000;
assign F[45][25] = 9'b100000000;
assign F[45][26] = 9'b100000000;
assign F[45][27] = 9'b100000000;
assign F[45][28] = 9'b100100100;
assign F[45][29] = 9'b100000000;
assign F[45][30] = 9'b100000000;
assign F[45][31] = 9'b100000000;
assign F[45][32] = 9'b100000000;
assign F[45][33] = 9'b100100100;
assign F[45][34] = 9'b100000000;
assign F[45][35] = 9'b100000000;
assign F[45][36] = 9'b100000000;
assign F[45][37] = 9'b100100100;
assign F[45][38] = 9'b100000000;
assign F[45][39] = 9'b100000000;
assign F[46][0] = 9'b100000000;
assign F[46][1] = 9'b100000000;
assign F[46][2] = 9'b100100100;
assign F[46][3] = 9'b100000000;
assign F[46][4] = 9'b100000000;
assign F[46][5] = 9'b100000000;
assign F[46][6] = 9'b100100100;
assign F[46][7] = 9'b100000000;
assign F[46][8] = 9'b100000000;
assign F[46][9] = 9'b100000000;
assign F[46][10] = 9'b100000000;
assign F[46][11] = 9'b100000000;
assign F[46][12] = 9'b100000000;
assign F[46][13] = 9'b100000000;
assign F[46][14] = 9'b100000000;
assign F[46][15] = 9'b100000000;
assign F[46][16] = 9'b100001000;
assign F[46][17] = 9'b100001000;
assign F[46][18] = 9'b101001101;
assign F[46][19] = 9'b101110001;
assign F[46][20] = 9'b101001101;
assign F[46][21] = 9'b100000100;
assign F[46][22] = 9'b100001101;
assign F[46][23] = 9'b100001101;
assign F[46][24] = 9'b100000000;
assign F[46][25] = 9'b100000000;
assign F[46][26] = 9'b100000000;
assign F[46][27] = 9'b100000000;
assign F[46][28] = 9'b100000000;
assign F[46][29] = 9'b100000000;
assign F[46][30] = 9'b100000000;
assign F[46][31] = 9'b100000000;
assign F[46][32] = 9'b100000000;
assign F[46][33] = 9'b100100100;
assign F[46][34] = 9'b100000000;
assign F[46][35] = 9'b100000000;
assign F[46][36] = 9'b100000000;
assign F[46][37] = 9'b100100100;
assign F[46][38] = 9'b100000000;
assign F[46][39] = 9'b100000000;
assign F[47][0] = 9'b100000000;
assign F[47][1] = 9'b100000000;
assign F[47][2] = 9'b100100100;
assign F[47][3] = 9'b100000000;
assign F[47][4] = 9'b100000000;
assign F[47][5] = 9'b100000000;
assign F[47][6] = 9'b100100100;
assign F[47][7] = 9'b100000000;
assign F[47][8] = 9'b100000000;
assign F[47][9] = 9'b100000000;
assign F[47][10] = 9'b100000000;
assign F[47][11] = 9'b100000000;
assign F[47][12] = 9'b100000000;
assign F[47][13] = 9'b100000000;
assign F[47][14] = 9'b100000000;
assign F[47][15] = 9'b100000000;
assign F[47][16] = 9'b100000000;
assign F[47][17] = 9'b100001000;
assign F[47][18] = 9'b101010001;
assign F[47][19] = 9'b101001101;
assign F[47][20] = 9'b100101101;
assign F[47][21] = 9'b100101101;
assign F[47][22] = 9'b100001101;
assign F[47][23] = 9'b100000000;
assign F[47][24] = 9'b100000000;
assign F[47][25] = 9'b100000000;
assign F[47][26] = 9'b100000000;
assign F[47][27] = 9'b100000000;
assign F[47][28] = 9'b100000000;
assign F[47][29] = 9'b100000000;
assign F[47][30] = 9'b100000000;
assign F[47][31] = 9'b100000000;
assign F[47][32] = 9'b100000000;
assign F[47][33] = 9'b100100100;
assign F[47][34] = 9'b100000000;
assign F[47][35] = 9'b100000000;
assign F[47][36] = 9'b100000000;
assign F[47][37] = 9'b100100100;
assign F[47][38] = 9'b100000000;
assign F[47][39] = 9'b100000000;
assign F[48][0] = 9'b100000000;
assign F[48][1] = 9'b100000000;
assign F[48][2] = 9'b100100100;
assign F[48][3] = 9'b100100100;
assign F[48][4] = 9'b100100100;
assign F[48][5] = 9'b100100100;
assign F[48][6] = 9'b100100100;
assign F[48][7] = 9'b100000000;
assign F[48][8] = 9'b100000000;
assign F[48][9] = 9'b100000000;
assign F[48][10] = 9'b100000000;
assign F[48][14] = 9'b100000000;
assign F[48][15] = 9'b100000000;
assign F[48][16] = 9'b100000000;
assign F[48][17] = 9'b100001000;
assign F[48][18] = 9'b101010001;
assign F[48][19] = 9'b100101001;
assign F[48][20] = 9'b100101001;
assign F[48][21] = 9'b101110101;
assign F[48][22] = 9'b100001101;
assign F[48][23] = 9'b100000000;
assign F[48][24] = 9'b100000000;
assign F[48][25] = 9'b100000000;
assign F[48][29] = 9'b100000000;
assign F[48][30] = 9'b100000000;
assign F[48][31] = 9'b100000000;
assign F[48][32] = 9'b100000000;
assign F[48][33] = 9'b100100100;
assign F[48][34] = 9'b100100100;
assign F[48][35] = 9'b100100100;
assign F[48][36] = 9'b100100100;
assign F[48][37] = 9'b100100100;
assign F[48][38] = 9'b100000000;
assign F[48][39] = 9'b100000000;
assign F[49][1] = 9'b100000000;
assign F[49][2] = 9'b100000000;
assign F[49][3] = 9'b100000000;
assign F[49][4] = 9'b100000000;
assign F[49][5] = 9'b100000000;
assign F[49][6] = 9'b100000000;
assign F[49][7] = 9'b100000000;
assign F[49][8] = 9'b100000000;
assign F[49][15] = 9'b100000000;
assign F[49][16] = 9'b100000000;
assign F[49][17] = 9'b100001000;
assign F[49][18] = 9'b101010001;
assign F[49][19] = 9'b110010001;
assign F[49][20] = 9'b110010010;
assign F[49][21] = 9'b101010001;
assign F[49][22] = 9'b100001101;
assign F[49][23] = 9'b100000000;
assign F[49][24] = 9'b100000000;
assign F[49][31] = 9'b100000000;
assign F[49][32] = 9'b100000000;
assign F[49][33] = 9'b100000000;
assign F[49][34] = 9'b100000000;
assign F[49][35] = 9'b100000000;
assign F[49][36] = 9'b100000000;
assign F[49][37] = 9'b100000000;
assign F[49][38] = 9'b100000000;
assign F[50][2] = 9'b100000000;
assign F[50][3] = 9'b100000000;
assign F[50][4] = 9'b100000000;
assign F[50][5] = 9'b100000000;
assign F[50][6] = 9'b100000000;
assign F[50][16] = 9'b100000000;
assign F[50][17] = 9'b100001000;
assign F[50][18] = 9'b100101101;
assign F[50][19] = 9'b100101101;
assign F[50][20] = 9'b100101101;
assign F[50][21] = 9'b100010001;
assign F[50][22] = 9'b100001101;
assign F[50][23] = 9'b100000000;
assign F[50][33] = 9'b100000000;
assign F[50][34] = 9'b100000000;
assign F[50][35] = 9'b100000000;
assign F[50][36] = 9'b100000000;
assign F[50][37] = 9'b100000000;
assign F[51][16] = 9'b100000000;
assign F[51][17] = 9'b100001000;
assign F[51][18] = 9'b100001111;
assign F[51][19] = 9'b100110111;
assign F[51][20] = 9'b100011100;
assign F[51][21] = 9'b100011100;
assign F[51][22] = 9'b100001101;
assign F[51][23] = 9'b100000000;
assign F[52][16] = 9'b100000000;
assign F[52][17] = 9'b100000100;
assign F[52][18] = 9'b100101101;
assign F[52][19] = 9'b100101101;
assign F[52][20] = 9'b100110001;
assign F[52][21] = 9'b100110001;
assign F[52][22] = 9'b100001000;
assign F[52][23] = 9'b100000000;
assign F[53][1] = 9'b100000000;
assign F[53][2] = 9'b100000000;
assign F[53][3] = 9'b100000000;
assign F[53][4] = 9'b100000000;
assign F[53][5] = 9'b100000000;
assign F[53][6] = 9'b100000000;
assign F[53][7] = 9'b100000000;
assign F[53][8] = 9'b100000000;
assign F[53][17] = 9'b100000000;
assign F[53][18] = 9'b100101001;
assign F[53][19] = 9'b101001101;
assign F[53][20] = 9'b101010001;
assign F[53][21] = 9'b101001101;
assign F[53][22] = 9'b100000000;
assign F[53][30] = 9'b100000000;
assign F[53][31] = 9'b100000000;
assign F[53][32] = 9'b100000000;
assign F[53][33] = 9'b100000000;
assign F[53][34] = 9'b100000000;
assign F[53][35] = 9'b100000000;
assign F[53][36] = 9'b100000000;
assign F[53][37] = 9'b100000000;
assign F[54][1] = 9'b100000000;
assign F[54][2] = 9'b100000100;
assign F[54][3] = 9'b100000100;
assign F[54][4] = 9'b101001001;
assign F[54][5] = 9'b110010001;
assign F[54][6] = 9'b110001101;
assign F[54][7] = 9'b100000000;
assign F[54][8] = 9'b100100100;
assign F[54][9] = 9'b100000000;
assign F[54][10] = 9'b100000000;
assign F[54][11] = 9'b100000000;
assign F[54][12] = 9'b100000000;
assign F[54][17] = 9'b100000000;
assign F[54][18] = 9'b100001000;
assign F[54][19] = 9'b101001000;
assign F[54][20] = 9'b101001000;
assign F[54][21] = 9'b100001101;
assign F[54][22] = 9'b100000000;
assign F[54][25] = 9'b100000000;
assign F[54][26] = 9'b100000000;
assign F[54][27] = 9'b100100100;
assign F[54][28] = 9'b100000000;
assign F[54][29] = 9'b100000000;
assign F[54][30] = 9'b100000000;
assign F[54][31] = 9'b100000000;
assign F[54][32] = 9'b100000000;
assign F[54][33] = 9'b110010001;
assign F[54][34] = 9'b101001001;
assign F[54][35] = 9'b100001000;
assign F[54][36] = 9'b100001000;
assign F[54][37] = 9'b100000000;
assign F[55][1] = 9'b100000000;
assign F[55][2] = 9'b100000100;
assign F[55][3] = 9'b100001000;
assign F[55][4] = 9'b100000100;
assign F[55][5] = 9'b100101001;
assign F[55][6] = 9'b100101000;
assign F[55][7] = 9'b100100100;
assign F[55][8] = 9'b110010010;
assign F[55][9] = 9'b100100100;
assign F[55][10] = 9'b110001101;
assign F[55][11] = 9'b101001001;
assign F[55][12] = 9'b100100100;
assign F[55][13] = 9'b101001000;
assign F[55][14] = 9'b100000000;
assign F[55][15] = 9'b100000000;
assign F[55][16] = 9'b100000000;
assign F[55][17] = 9'b100000000;
assign F[55][18] = 9'b100000100;
assign F[55][19] = 9'b100000100;
assign F[55][20] = 9'b100001000;
assign F[55][21] = 9'b100001000;
assign F[55][22] = 9'b100000000;
assign F[55][23] = 9'b100000000;
assign F[55][24] = 9'b100000000;
assign F[55][25] = 9'b100000000;
assign F[55][26] = 9'b101101101;
assign F[55][27] = 9'b110010010;
assign F[55][28] = 9'b101101101;
assign F[55][29] = 9'b100000000;
assign F[55][30] = 9'b100000000;
assign F[55][31] = 9'b100000100;
assign F[55][32] = 9'b100000100;
assign F[55][33] = 9'b100101001;
assign F[55][34] = 9'b100000100;
assign F[55][35] = 9'b100001101;
assign F[55][36] = 9'b100001000;
assign F[55][37] = 9'b100000000;
assign F[56][1] = 9'b100000000;
assign F[56][2] = 9'b100101100;
assign F[56][3] = 9'b101010100;
assign F[56][4] = 9'b100110000;
assign F[56][5] = 9'b100110000;
assign F[56][6] = 9'b100110000;
assign F[56][7] = 9'b100001000;
assign F[56][8] = 9'b100001000;
assign F[56][9] = 9'b100001000;
assign F[56][10] = 9'b100001000;
assign F[56][11] = 9'b100000100;
assign F[56][12] = 9'b101001001;
assign F[56][13] = 9'b101101101;
assign F[56][14] = 9'b100100100;
assign F[56][15] = 9'b100100100;
assign F[56][16] = 9'b100100000;
assign F[56][17] = 9'b100000000;
assign F[56][18] = 9'b100000000;
assign F[56][19] = 9'b100000000;
assign F[56][20] = 9'b100000000;
assign F[56][21] = 9'b100000000;
assign F[56][22] = 9'b100000000;
assign F[56][23] = 9'b100100000;
assign F[56][24] = 9'b100100100;
assign F[56][25] = 9'b100100100;
assign F[56][26] = 9'b100100100;
assign F[56][27] = 9'b100000100;
assign F[56][28] = 9'b100000100;
assign F[56][29] = 9'b101001001;
assign F[56][30] = 9'b110010101;
assign F[56][31] = 9'b100110100;
assign F[56][32] = 9'b100110100;
assign F[56][33] = 9'b100110000;
assign F[56][34] = 9'b100110000;
assign F[56][35] = 9'b100001100;
assign F[56][36] = 9'b100000100;
assign F[56][37] = 9'b100000000;
assign F[57][2] = 9'b100000100;
assign F[57][3] = 9'b100100100;
assign F[57][4] = 9'b100000100;
assign F[57][5] = 9'b100100100;
assign F[57][6] = 9'b100101000;
assign F[57][7] = 9'b101010000;
assign F[57][8] = 9'b110010001;
assign F[57][9] = 9'b100001000;
assign F[57][10] = 9'b101110001;
assign F[57][11] = 9'b101001101;
assign F[57][12] = 9'b100000100;
assign F[57][13] = 9'b100000100;
assign F[57][14] = 9'b100001000;
assign F[57][15] = 9'b100001000;
assign F[57][16] = 9'b100100100;
assign F[57][17] = 9'b100100100;
assign F[57][18] = 9'b100001000;
assign F[57][19] = 9'b100000100;
assign F[57][20] = 9'b100000100;
assign F[57][21] = 9'b100001000;
assign F[57][22] = 9'b100101000;
assign F[57][23] = 9'b100101000;
assign F[57][24] = 9'b100001000;
assign F[57][25] = 9'b100001101;
assign F[57][26] = 9'b100001000;
assign F[57][27] = 9'b101110001;
assign F[57][28] = 9'b101010001;
assign F[57][29] = 9'b100010000;
assign F[57][30] = 9'b101111100;
assign F[57][31] = 9'b100000100;
assign F[57][32] = 9'b100000100;
assign F[57][33] = 9'b100000100;
assign F[57][34] = 9'b100100100;
assign F[57][35] = 9'b100000100;
assign F[58][7] = 9'b100000000;
assign F[58][8] = 9'b100000000;
assign F[58][9] = 9'b100000000;
assign F[58][10] = 9'b100000000;
assign F[58][11] = 9'b100000000;
assign F[58][12] = 9'b100000000;
assign F[58][13] = 9'b100000000;
assign F[58][14] = 9'b100000000;
assign F[58][15] = 9'b100000100;
assign F[58][16] = 9'b100000100;
assign F[58][17] = 9'b100000100;
assign F[58][18] = 9'b100001000;
assign F[58][19] = 9'b100001000;
assign F[58][20] = 9'b100001000;
assign F[58][21] = 9'b100001101;
assign F[58][22] = 9'b100001000;
assign F[58][23] = 9'b100001000;
assign F[58][24] = 9'b100001000;
assign F[58][25] = 9'b100000000;
assign F[58][26] = 9'b100000000;
assign F[58][27] = 9'b100000000;
assign F[58][28] = 9'b100000000;
assign F[58][29] = 9'b100000000;
assign F[58][30] = 9'b100000000;
assign F[59][18] = 9'b100000000;
assign F[59][19] = 9'b100000000;
assign F[59][20] = 9'b100000000;
assign F[59][21] = 9'b100000000;
//Total de Lineas = 1727
endmodule

