`timescale 1ns / 1ps
module carroazul (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (F[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= F[vcount- posy][hcount- posx][7:5];
				green <= F[vcount- posy][hcount- posx][4:2];
            blue 	<= F[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 25;
parameter RESOLUCION_Y = 70;
wire [8:0] F[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign F[6][10] = 9'b101100100;
assign F[6][11] = 9'b100000000;
assign F[6][12] = 9'b100000000;
assign F[6][13] = 9'b100000000;
assign F[6][14] = 9'b100000000;
assign F[6][15] = 9'b101000100;
assign F[6][16] = 9'b111100100;
assign F[7][6] = 9'b110000100;
assign F[7][7] = 9'b110100100;
assign F[7][8] = 9'b110100100;
assign F[7][9] = 9'b111100100;
assign F[7][10] = 9'b100100100;
assign F[7][11] = 9'b100000000;
assign F[7][12] = 9'b100000100;
assign F[7][13] = 9'b100000100;
assign F[7][14] = 9'b100000100;
assign F[7][15] = 9'b100000100;
assign F[7][16] = 9'b110100100;
assign F[7][17] = 9'b110100100;
assign F[7][18] = 9'b110100100;
assign F[7][19] = 9'b110000100;
assign F[8][5] = 9'b100000100;
assign F[8][6] = 9'b101100100;
assign F[8][7] = 9'b111100100;
assign F[8][8] = 9'b110100100;
assign F[8][9] = 9'b101100100;
assign F[8][10] = 9'b100000000;
assign F[8][11] = 9'b100000100;
assign F[8][12] = 9'b100000100;
assign F[8][13] = 9'b100000100;
assign F[8][14] = 9'b100000100;
assign F[8][15] = 9'b100000000;
assign F[8][16] = 9'b101000100;
assign F[8][17] = 9'b110100100;
assign F[8][18] = 9'b110100100;
assign F[8][19] = 9'b110000100;
assign F[8][20] = 9'b100100100;
assign F[9][5] = 9'b100000100;
assign F[9][6] = 9'b101100100;
assign F[9][7] = 9'b110100100;
assign F[9][8] = 9'b110000100;
assign F[9][9] = 9'b100000000;
assign F[9][10] = 9'b100000000;
assign F[9][11] = 9'b100000100;
assign F[9][12] = 9'b101101100;
assign F[9][13] = 9'b110010000;
assign F[9][14] = 9'b100000100;
assign F[9][15] = 9'b100000000;
assign F[9][16] = 9'b100000000;
assign F[9][17] = 9'b110000100;
assign F[9][18] = 9'b110100100;
assign F[9][19] = 9'b110000100;
assign F[9][20] = 9'b100100100;
assign F[10][5] = 9'b100000100;
assign F[10][6] = 9'b101100100;
assign F[10][7] = 9'b111100100;
assign F[10][8] = 9'b101100100;
assign F[10][9] = 9'b100000000;
assign F[10][10] = 9'b100000000;
assign F[10][11] = 9'b100000100;
assign F[10][12] = 9'b100000100;
assign F[10][13] = 9'b100101000;
assign F[10][14] = 9'b100000100;
assign F[10][15] = 9'b100000000;
assign F[10][16] = 9'b100000000;
assign F[10][17] = 9'b101000100;
assign F[10][18] = 9'b111100100;
assign F[10][19] = 9'b110000100;
assign F[10][20] = 9'b100100100;
assign F[11][5] = 9'b100000100;
assign F[11][6] = 9'b101100100;
assign F[11][7] = 9'b111100100;
assign F[11][8] = 9'b101000100;
assign F[11][9] = 9'b100000100;
assign F[11][10] = 9'b100000000;
assign F[11][11] = 9'b100000000;
assign F[11][12] = 9'b100101001;
assign F[11][13] = 9'b101001001;
assign F[11][14] = 9'b100000100;
assign F[11][15] = 9'b100000000;
assign F[11][16] = 9'b100000100;
assign F[11][17] = 9'b100100100;
assign F[11][18] = 9'b110100100;
assign F[11][19] = 9'b110000100;
assign F[11][20] = 9'b100100100;
assign F[12][5] = 9'b100000100;
assign F[12][6] = 9'b101100100;
assign F[12][7] = 9'b111100100;
assign F[12][8] = 9'b100100100;
assign F[12][9] = 9'b100000000;
assign F[12][10] = 9'b100000000;
assign F[12][11] = 9'b100000000;
assign F[12][12] = 9'b100101001;
assign F[12][13] = 9'b101001101;
assign F[12][14] = 9'b100000100;
assign F[12][15] = 9'b100000000;
assign F[12][16] = 9'b100000000;
assign F[12][17] = 9'b100000000;
assign F[12][18] = 9'b110100100;
assign F[12][19] = 9'b110000100;
assign F[12][20] = 9'b100100100;
assign F[13][5] = 9'b100000100;
assign F[13][6] = 9'b101100100;
assign F[13][7] = 9'b111100100;
assign F[13][11] = 9'b100000100;
assign F[13][12] = 9'b100101001;
assign F[13][13] = 9'b101001101;
assign F[13][14] = 9'b100000100;
assign F[13][19] = 9'b110000100;
assign F[13][20] = 9'b100100100;
assign F[14][4] = 9'b100000000;
assign F[14][5] = 9'b100000000;
assign F[14][6] = 9'b100000000;
assign F[14][7] = 9'b100000000;
assign F[14][11] = 9'b100000100;
assign F[14][12] = 9'b100000101;
assign F[14][13] = 9'b100000101;
assign F[14][14] = 9'b100000100;
assign F[14][19] = 9'b100000000;
assign F[14][20] = 9'b100000000;
assign F[14][21] = 9'b100000000;
assign F[14][22] = 9'b100000000;
assign F[15][3] = 9'b100000000;
assign F[15][4] = 9'b100000000;
assign F[15][5] = 9'b100000000;
assign F[15][6] = 9'b100000000;
assign F[15][7] = 9'b100000000;
assign F[15][11] = 9'b100000100;
assign F[15][12] = 9'b100000101;
assign F[15][13] = 9'b100000101;
assign F[15][14] = 9'b100000100;
assign F[15][18] = 9'b100000000;
assign F[15][19] = 9'b100000000;
assign F[15][20] = 9'b100000000;
assign F[15][21] = 9'b100000000;
assign F[15][22] = 9'b100000000;
assign F[16][3] = 9'b100000000;
assign F[16][4] = 9'b100000000;
assign F[16][5] = 9'b100000000;
assign F[16][6] = 9'b100000000;
assign F[16][7] = 9'b100000000;
assign F[16][11] = 9'b100000100;
assign F[16][12] = 9'b110110101;
assign F[16][13] = 9'b111111101;
assign F[16][14] = 9'b100101000;
assign F[16][18] = 9'b100000000;
assign F[16][19] = 9'b100000000;
assign F[16][20] = 9'b100000000;
assign F[16][21] = 9'b100000000;
assign F[16][22] = 9'b100000000;
assign F[17][3] = 9'b100000000;
assign F[17][4] = 9'b100000000;
assign F[17][5] = 9'b100000000;
assign F[17][6] = 9'b100000000;
assign F[17][7] = 9'b100000000;
assign F[17][11] = 9'b100000100;
assign F[17][12] = 9'b101101101;
assign F[17][13] = 9'b110010001;
assign F[17][14] = 9'b100000100;
assign F[17][18] = 9'b100000000;
assign F[17][19] = 9'b100000000;
assign F[17][20] = 9'b100000000;
assign F[17][21] = 9'b100000000;
assign F[17][22] = 9'b100000000;
assign F[18][3] = 9'b100000000;
assign F[18][4] = 9'b100000000;
assign F[18][5] = 9'b100000000;
assign F[18][6] = 9'b100000000;
assign F[18][7] = 9'b100000000;
assign F[18][8] = 9'b100100100;
assign F[18][9] = 9'b100100100;
assign F[18][10] = 9'b100100100;
assign F[18][11] = 9'b100000100;
assign F[18][12] = 9'b101001101;
assign F[18][13] = 9'b101101101;
assign F[18][14] = 9'b100000100;
assign F[18][15] = 9'b100000100;
assign F[18][16] = 9'b100100100;
assign F[18][17] = 9'b100100100;
assign F[18][18] = 9'b100000000;
assign F[18][19] = 9'b100000000;
assign F[18][20] = 9'b100000000;
assign F[18][21] = 9'b100000000;
assign F[18][22] = 9'b100000000;
assign F[19][3] = 9'b100000000;
assign F[19][4] = 9'b100000000;
assign F[19][5] = 9'b100000000;
assign F[19][6] = 9'b100000000;
assign F[19][7] = 9'b100000000;
assign F[19][8] = 9'b100100100;
assign F[19][9] = 9'b100100100;
assign F[19][11] = 9'b100000100;
assign F[19][12] = 9'b101001101;
assign F[19][13] = 9'b101101101;
assign F[19][14] = 9'b100000100;
assign F[19][15] = 9'b100000000;
assign F[19][16] = 9'b100100100;
assign F[19][17] = 9'b100100100;
assign F[19][18] = 9'b100000000;
assign F[19][19] = 9'b100000000;
assign F[19][20] = 9'b100000000;
assign F[19][21] = 9'b100000000;
assign F[19][22] = 9'b100000000;
assign F[20][3] = 9'b100000000;
assign F[20][4] = 9'b100000000;
assign F[20][5] = 9'b100000000;
assign F[20][6] = 9'b100000000;
assign F[20][7] = 9'b100000000;
assign F[20][9] = 9'b100100100;
assign F[20][10] = 9'b100100100;
assign F[20][11] = 9'b100000100;
assign F[20][12] = 9'b100000101;
assign F[20][13] = 9'b100000101;
assign F[20][14] = 9'b100000100;
assign F[20][15] = 9'b100000100;
assign F[20][16] = 9'b100100100;
assign F[20][17] = 9'b100100100;
assign F[20][18] = 9'b100000000;
assign F[20][19] = 9'b100000000;
assign F[20][20] = 9'b100000000;
assign F[20][21] = 9'b100000000;
assign F[20][22] = 9'b100000000;
assign F[21][3] = 9'b100000000;
assign F[21][4] = 9'b100000000;
assign F[21][5] = 9'b100000000;
assign F[21][6] = 9'b100000000;
assign F[21][7] = 9'b100000000;
assign F[21][10] = 9'b100000100;
assign F[21][11] = 9'b100000100;
assign F[21][12] = 9'b100101001;
assign F[21][13] = 9'b101001001;
assign F[21][14] = 9'b100000100;
assign F[21][15] = 9'b100000100;
assign F[21][18] = 9'b100000000;
assign F[21][19] = 9'b100000000;
assign F[21][20] = 9'b100000000;
assign F[21][21] = 9'b100000000;
assign F[21][22] = 9'b100000000;
assign F[22][3] = 9'b100000000;
assign F[22][4] = 9'b100000000;
assign F[22][5] = 9'b100000000;
assign F[22][6] = 9'b100000000;
assign F[22][7] = 9'b100000000;
assign F[22][11] = 9'b100000000;
assign F[22][12] = 9'b101110010;
assign F[22][13] = 9'b111111111;
assign F[22][14] = 9'b100000100;
assign F[22][18] = 9'b100000000;
assign F[22][19] = 9'b100000000;
assign F[22][20] = 9'b100000000;
assign F[22][21] = 9'b100000000;
assign F[22][22] = 9'b100000000;
assign F[23][3] = 9'b100000000;
assign F[23][4] = 9'b100000000;
assign F[23][5] = 9'b100000000;
assign F[23][6] = 9'b100000000;
assign F[23][7] = 9'b100000000;
assign F[23][11] = 9'b100000000;
assign F[23][12] = 9'b101110010;
assign F[23][13] = 9'b111111111;
assign F[23][14] = 9'b100000100;
assign F[23][15] = 9'b100000100;
assign F[23][18] = 9'b100000000;
assign F[23][19] = 9'b100000000;
assign F[23][20] = 9'b100000000;
assign F[23][21] = 9'b100000000;
assign F[23][22] = 9'b100000000;
assign F[24][11] = 9'b100000000;
assign F[24][12] = 9'b101110010;
assign F[24][13] = 9'b111111111;
assign F[24][14] = 9'b100000100;
assign F[24][15] = 9'b100000100;
assign F[25][11] = 9'b100000000;
assign F[25][12] = 9'b110010010;
assign F[25][13] = 9'b111111111;
assign F[25][14] = 9'b100000100;
assign F[25][15] = 9'b100000100;
assign F[26][10] = 9'b100000100;
assign F[26][11] = 9'b100000100;
assign F[26][12] = 9'b101001101;
assign F[26][13] = 9'b101110001;
assign F[26][14] = 9'b100000100;
assign F[26][15] = 9'b100000100;
assign F[27][10] = 9'b100000100;
assign F[27][11] = 9'b100000100;
assign F[27][12] = 9'b100000100;
assign F[27][13] = 9'b100000100;
assign F[27][14] = 9'b100000100;
assign F[27][15] = 9'b100000100;
assign F[28][10] = 9'b100000100;
assign F[28][11] = 9'b100000100;
assign F[28][12] = 9'b100000100;
assign F[28][13] = 9'b100000100;
assign F[28][14] = 9'b100000100;
assign F[28][15] = 9'b100000100;
assign F[29][6] = 9'b100000000;
assign F[29][7] = 9'b100000000;
assign F[29][8] = 9'b100000000;
assign F[29][9] = 9'b100100000;
assign F[29][10] = 9'b100100100;
assign F[29][11] = 9'b100000100;
assign F[29][12] = 9'b100000100;
assign F[29][13] = 9'b100000100;
assign F[29][14] = 9'b100000100;
assign F[29][15] = 9'b100000100;
assign F[29][16] = 9'b101000000;
assign F[29][17] = 9'b100000000;
assign F[29][18] = 9'b100000000;
assign F[29][19] = 9'b100000000;
assign F[30][6] = 9'b100000000;
assign F[30][7] = 9'b100000100;
assign F[30][8] = 9'b100000100;
assign F[30][9] = 9'b101100100;
assign F[30][10] = 9'b101100100;
assign F[30][11] = 9'b100000000;
assign F[30][12] = 9'b100000000;
assign F[30][13] = 9'b100000000;
assign F[30][14] = 9'b100000000;
assign F[30][15] = 9'b100100100;
assign F[30][16] = 9'b110000100;
assign F[30][17] = 9'b100000100;
assign F[30][18] = 9'b100000100;
assign F[30][19] = 9'b100000000;
assign F[31][6] = 9'b100000100;
assign F[31][7] = 9'b100000101;
assign F[31][8] = 9'b100000100;
assign F[31][9] = 9'b101100100;
assign F[31][10] = 9'b101100100;
assign F[31][11] = 9'b100000000;
assign F[31][12] = 9'b100000000;
assign F[31][13] = 9'b100000000;
assign F[31][14] = 9'b100000000;
assign F[31][15] = 9'b100100100;
assign F[31][16] = 9'b110000100;
assign F[31][17] = 9'b100000100;
assign F[31][18] = 9'b100000101;
assign F[31][19] = 9'b100000100;
assign F[32][6] = 9'b100000100;
assign F[32][7] = 9'b100000101;
assign F[32][8] = 9'b100000101;
assign F[32][9] = 9'b101100100;
assign F[32][10] = 9'b101100100;
assign F[32][11] = 9'b100000000;
assign F[32][12] = 9'b100000000;
assign F[32][13] = 9'b100000000;
assign F[32][14] = 9'b100000000;
assign F[32][15] = 9'b100100100;
assign F[32][16] = 9'b110000100;
assign F[32][17] = 9'b100000100;
assign F[32][18] = 9'b100000101;
assign F[32][19] = 9'b100000100;
assign F[33][6] = 9'b100000100;
assign F[33][7] = 9'b100000101;
assign F[33][8] = 9'b100000101;
assign F[33][9] = 9'b101100100;
assign F[33][10] = 9'b101100100;
assign F[33][11] = 9'b100000000;
assign F[33][12] = 9'b100000000;
assign F[33][13] = 9'b100000000;
assign F[33][14] = 9'b100000000;
assign F[33][15] = 9'b100100100;
assign F[33][16] = 9'b110000100;
assign F[33][17] = 9'b100000100;
assign F[33][18] = 9'b100000101;
assign F[33][19] = 9'b100000100;
assign F[34][6] = 9'b100000100;
assign F[34][7] = 9'b100000101;
assign F[34][8] = 9'b100000101;
assign F[34][9] = 9'b101000100;
assign F[34][10] = 9'b101100100;
assign F[34][11] = 9'b100000100;
assign F[34][12] = 9'b100000000;
assign F[34][13] = 9'b100000000;
assign F[34][14] = 9'b100000000;
assign F[34][15] = 9'b101000100;
assign F[34][16] = 9'b110000100;
assign F[34][17] = 9'b100000100;
assign F[34][18] = 9'b100000101;
assign F[34][19] = 9'b100000100;
assign F[35][6] = 9'b100000100;
assign F[35][7] = 9'b100000101;
assign F[35][8] = 9'b100000101;
assign F[35][9] = 9'b101000000;
assign F[35][10] = 9'b110001000;
assign F[35][11] = 9'b110001100;
assign F[35][12] = 9'b100000000;
assign F[35][13] = 9'b100000000;
assign F[35][14] = 9'b101101100;
assign F[35][15] = 9'b101101000;
assign F[35][16] = 9'b110000000;
assign F[35][17] = 9'b100000100;
assign F[35][18] = 9'b100000101;
assign F[35][19] = 9'b100000100;
assign F[36][6] = 9'b100000100;
assign F[36][7] = 9'b100000101;
assign F[36][8] = 9'b100000101;
assign F[36][9] = 9'b101000100;
assign F[36][10] = 9'b101100100;
assign F[36][11] = 9'b111111100;
assign F[36][12] = 9'b101101100;
assign F[36][13] = 9'b101001000;
assign F[36][14] = 9'b111111100;
assign F[36][15] = 9'b101101000;
assign F[36][16] = 9'b110000000;
assign F[36][17] = 9'b100000100;
assign F[36][18] = 9'b100000101;
assign F[36][19] = 9'b100000100;
assign F[37][6] = 9'b100000100;
assign F[37][7] = 9'b100000101;
assign F[37][8] = 9'b100000101;
assign F[37][9] = 9'b101000100;
assign F[37][10] = 9'b101100100;
assign F[37][11] = 9'b110010000;
assign F[37][12] = 9'b100100100;
assign F[37][13] = 9'b100000000;
assign F[37][14] = 9'b110001100;
assign F[37][15] = 9'b101101000;
assign F[37][16] = 9'b110000000;
assign F[37][17] = 9'b100000100;
assign F[37][18] = 9'b100000101;
assign F[37][19] = 9'b100000100;
assign F[38][6] = 9'b100000100;
assign F[38][7] = 9'b100000100;
assign F[38][8] = 9'b100000100;
assign F[38][9] = 9'b101100100;
assign F[38][10] = 9'b101100100;
assign F[38][11] = 9'b110010000;
assign F[38][12] = 9'b110001100;
assign F[38][13] = 9'b101001000;
assign F[38][14] = 9'b111111100;
assign F[38][15] = 9'b101000100;
assign F[38][16] = 9'b110000100;
assign F[38][17] = 9'b100000100;
assign F[38][18] = 9'b100000100;
assign F[38][19] = 9'b100000100;
assign F[39][6] = 9'b100000000;
assign F[39][7] = 9'b100000100;
assign F[39][8] = 9'b100000100;
assign F[39][9] = 9'b101100100;
assign F[39][10] = 9'b101000000;
assign F[39][11] = 9'b110010000;
assign F[39][12] = 9'b110110000;
assign F[39][13] = 9'b101101100;
assign F[39][14] = 9'b111111100;
assign F[39][15] = 9'b100100100;
assign F[39][16] = 9'b110000100;
assign F[39][17] = 9'b100000100;
assign F[39][18] = 9'b100000100;
assign F[39][19] = 9'b100000000;
assign F[40][6] = 9'b100000000;
assign F[40][7] = 9'b100000100;
assign F[40][8] = 9'b100000100;
assign F[40][9] = 9'b101100100;
assign F[40][10] = 9'b101000000;
assign F[40][11] = 9'b101101100;
assign F[40][12] = 9'b110110000;
assign F[40][13] = 9'b101101100;
assign F[40][14] = 9'b110110100;
assign F[40][15] = 9'b100100100;
assign F[40][16] = 9'b110000100;
assign F[40][17] = 9'b100000100;
assign F[40][18] = 9'b100000100;
assign F[40][19] = 9'b100000000;
assign F[41][6] = 9'b100000000;
assign F[41][7] = 9'b100000000;
assign F[41][8] = 9'b100000100;
assign F[41][9] = 9'b101100100;
assign F[41][10] = 9'b101000000;
assign F[41][11] = 9'b101001100;
assign F[41][12] = 9'b110110000;
assign F[41][13] = 9'b101101100;
assign F[41][14] = 9'b110010000;
assign F[41][15] = 9'b100000000;
assign F[41][16] = 9'b110000100;
assign F[41][17] = 9'b100000100;
assign F[41][18] = 9'b100000100;
assign F[41][19] = 9'b100000000;
assign F[42][6] = 9'b100000000;
assign F[42][7] = 9'b100000000;
assign F[42][8] = 9'b100000100;
assign F[42][9] = 9'b101100100;
assign F[42][10] = 9'b101000000;
assign F[42][11] = 9'b100101000;
assign F[42][12] = 9'b110010000;
assign F[42][13] = 9'b101101100;
assign F[42][14] = 9'b101101100;
assign F[42][15] = 9'b100000000;
assign F[42][16] = 9'b110000100;
assign F[42][17] = 9'b100000100;
assign F[42][18] = 9'b100000000;
assign F[42][19] = 9'b100000000;
assign F[43][6] = 9'b100000000;
assign F[43][7] = 9'b100000000;
assign F[43][8] = 9'b100000100;
assign F[43][9] = 9'b101100100;
assign F[43][10] = 9'b101100000;
assign F[43][11] = 9'b100101000;
assign F[43][12] = 9'b110010000;
assign F[43][13] = 9'b101101100;
assign F[43][14] = 9'b101001100;
assign F[43][15] = 9'b100000000;
assign F[43][16] = 9'b110000100;
assign F[43][17] = 9'b100000100;
assign F[43][18] = 9'b100000000;
assign F[43][19] = 9'b100000000;
assign F[44][6] = 9'b100000000;
assign F[44][7] = 9'b100000000;
assign F[44][8] = 9'b100000000;
assign F[44][9] = 9'b101100100;
assign F[44][10] = 9'b101100100;
assign F[44][11] = 9'b100000100;
assign F[44][12] = 9'b110001100;
assign F[44][13] = 9'b101101100;
assign F[44][14] = 9'b101001000;
assign F[44][15] = 9'b100100000;
assign F[44][16] = 9'b110000100;
assign F[44][17] = 9'b100000000;
assign F[44][18] = 9'b100000000;
assign F[44][19] = 9'b100000000;
assign F[45][6] = 9'b100000000;
assign F[45][7] = 9'b100000000;
assign F[45][8] = 9'b100000000;
assign F[45][9] = 9'b101100100;
assign F[45][10] = 9'b101100100;
assign F[45][11] = 9'b100000100;
assign F[45][12] = 9'b101101100;
assign F[45][13] = 9'b101101100;
assign F[45][14] = 9'b100101000;
assign F[45][15] = 9'b100100100;
assign F[45][16] = 9'b110000100;
assign F[45][17] = 9'b100000000;
assign F[45][18] = 9'b100000000;
assign F[45][19] = 9'b100000000;
assign F[46][6] = 9'b100000000;
assign F[46][7] = 9'b100000000;
assign F[46][8] = 9'b100000000;
assign F[46][9] = 9'b101000000;
assign F[46][10] = 9'b101100100;
assign F[46][11] = 9'b100000100;
assign F[46][12] = 9'b101001100;
assign F[46][13] = 9'b101101100;
assign F[46][14] = 9'b100000100;
assign F[46][15] = 9'b100100100;
assign F[46][16] = 9'b101100100;
assign F[46][17] = 9'b100000000;
assign F[46][18] = 9'b100000000;
assign F[46][19] = 9'b100000000;
assign F[47][6] = 9'b100000000;
assign F[47][7] = 9'b100000000;
assign F[47][8] = 9'b100000000;
assign F[47][9] = 9'b100100000;
assign F[47][10] = 9'b101000100;
assign F[47][11] = 9'b100000100;
assign F[47][12] = 9'b100101000;
assign F[47][13] = 9'b101001000;
assign F[47][14] = 9'b100000100;
assign F[47][15] = 9'b100100100;
assign F[47][16] = 9'b101000000;
assign F[47][17] = 9'b100000000;
assign F[47][18] = 9'b100000000;
assign F[47][19] = 9'b100000000;
assign F[48][6] = 9'b100000000;
assign F[48][7] = 9'b100000000;
assign F[48][8] = 9'b100000000;
assign F[48][9] = 9'b100100000;
assign F[48][10] = 9'b101000100;
assign F[48][11] = 9'b100000100;
assign F[48][12] = 9'b100101000;
assign F[48][13] = 9'b100101000;
assign F[48][14] = 9'b100000100;
assign F[48][15] = 9'b100100100;
assign F[48][16] = 9'b100100000;
assign F[48][17] = 9'b100000000;
assign F[48][18] = 9'b100000000;
assign F[48][19] = 9'b100000000;
assign F[49][6] = 9'b100000000;
assign F[49][7] = 9'b100000000;
assign F[49][8] = 9'b100000000;
assign F[49][9] = 9'b100000000;
assign F[49][10] = 9'b100100100;
assign F[49][11] = 9'b100000100;
assign F[49][12] = 9'b100000100;
assign F[49][13] = 9'b100000100;
assign F[49][14] = 9'b100000100;
assign F[49][15] = 9'b100000100;
assign F[49][16] = 9'b100000000;
assign F[49][17] = 9'b100000000;
assign F[49][18] = 9'b100000000;
assign F[49][19] = 9'b100000000;
assign F[50][5] = 9'b100000000;
assign F[50][6] = 9'b100000000;
assign F[50][7] = 9'b100000000;
assign F[50][8] = 9'b100000000;
assign F[50][9] = 9'b100000000;
assign F[50][10] = 9'b100000100;
assign F[50][11] = 9'b100000100;
assign F[50][12] = 9'b100000100;
assign F[50][13] = 9'b100000100;
assign F[50][14] = 9'b100000100;
assign F[50][15] = 9'b100000100;
assign F[50][16] = 9'b100000000;
assign F[50][18] = 9'b100000000;
assign F[50][19] = 9'b100000000;
assign F[50][20] = 9'b100000000;
assign F[50][21] = 9'b100000000;
assign F[51][3] = 9'b100000000;
assign F[51][4] = 9'b100000000;
assign F[51][5] = 9'b100000000;
assign F[51][6] = 9'b100000000;
assign F[51][7] = 9'b100000000;
assign F[51][8] = 9'b100000000;
assign F[51][10] = 9'b100000000;
assign F[51][11] = 9'b100000100;
assign F[51][12] = 9'b100000100;
assign F[51][13] = 9'b100000100;
assign F[51][14] = 9'b100000100;
assign F[51][15] = 9'b100000100;
assign F[51][16] = 9'b100000000;
assign F[51][17] = 9'b100000000;
assign F[51][18] = 9'b100000000;
assign F[51][19] = 9'b100000000;
assign F[51][20] = 9'b100000000;
assign F[51][21] = 9'b100000000;
assign F[51][22] = 9'b100000000;
assign F[52][3] = 9'b100000000;
assign F[52][4] = 9'b100000000;
assign F[52][5] = 9'b100000000;
assign F[52][6] = 9'b100000000;
assign F[52][7] = 9'b100000000;
assign F[52][8] = 9'b100000000;
assign F[52][9] = 9'b100000000;
assign F[52][10] = 9'b100000000;
assign F[52][11] = 9'b100000100;
assign F[52][12] = 9'b100000100;
assign F[52][13] = 9'b100000100;
assign F[52][14] = 9'b100000100;
assign F[52][15] = 9'b100000100;
assign F[52][16] = 9'b100000000;
assign F[52][17] = 9'b100000000;
assign F[52][18] = 9'b100000000;
assign F[52][19] = 9'b100000000;
assign F[52][20] = 9'b100000000;
assign F[52][21] = 9'b100000000;
assign F[52][22] = 9'b100000000;
assign F[53][3] = 9'b100000000;
assign F[53][4] = 9'b100000000;
assign F[53][5] = 9'b100000000;
assign F[53][6] = 9'b100000000;
assign F[53][7] = 9'b100000000;
assign F[53][8] = 9'b100000000;
assign F[53][10] = 9'b100000000;
assign F[53][11] = 9'b100000100;
assign F[53][12] = 9'b100000100;
assign F[53][13] = 9'b100000100;
assign F[53][14] = 9'b100000100;
assign F[53][15] = 9'b100000000;
assign F[53][16] = 9'b100000000;
assign F[53][17] = 9'b100000000;
assign F[53][18] = 9'b100000000;
assign F[53][19] = 9'b100000000;
assign F[53][20] = 9'b100000000;
assign F[53][21] = 9'b100000000;
assign F[53][22] = 9'b100000000;
assign F[54][3] = 9'b100000000;
assign F[54][4] = 9'b100000000;
assign F[54][5] = 9'b100000000;
assign F[54][6] = 9'b100000000;
assign F[54][7] = 9'b100000000;
assign F[54][8] = 9'b100000000;
assign F[54][9] = 9'b100100100;
assign F[54][10] = 9'b100100000;
assign F[54][11] = 9'b100000100;
assign F[54][12] = 9'b100000100;
assign F[54][13] = 9'b100000100;
assign F[54][14] = 9'b100000100;
assign F[54][15] = 9'b100100100;
assign F[54][16] = 9'b100100100;
assign F[54][17] = 9'b100000000;
assign F[54][18] = 9'b100000000;
assign F[54][19] = 9'b100000000;
assign F[54][20] = 9'b100000000;
assign F[54][21] = 9'b100000000;
assign F[54][22] = 9'b100000000;
assign F[55][3] = 9'b100000000;
assign F[55][4] = 9'b100000000;
assign F[55][5] = 9'b100000000;
assign F[55][6] = 9'b100000000;
assign F[55][7] = 9'b100000000;
assign F[55][8] = 9'b100000000;
assign F[55][9] = 9'b100100100;
assign F[55][10] = 9'b100100100;
assign F[55][11] = 9'b100000100;
assign F[55][12] = 9'b100000100;
assign F[55][13] = 9'b100000100;
assign F[55][14] = 9'b100000100;
assign F[55][15] = 9'b100100100;
assign F[55][16] = 9'b100100100;
assign F[55][17] = 9'b100000000;
assign F[55][18] = 9'b100000000;
assign F[55][19] = 9'b100000000;
assign F[55][20] = 9'b100000000;
assign F[55][21] = 9'b100000000;
assign F[55][22] = 9'b100000000;
assign F[56][3] = 9'b100000000;
assign F[56][4] = 9'b100000000;
assign F[56][5] = 9'b100000000;
assign F[56][6] = 9'b100000000;
assign F[56][7] = 9'b100000000;
assign F[56][8] = 9'b100000000;
assign F[56][9] = 9'b100100100;
assign F[56][10] = 9'b100100000;
assign F[56][11] = 9'b100000000;
assign F[56][12] = 9'b100000100;
assign F[56][13] = 9'b100000100;
assign F[56][14] = 9'b100000100;
assign F[56][15] = 9'b100000000;
assign F[56][16] = 9'b100100100;
assign F[56][17] = 9'b100000000;
assign F[56][18] = 9'b100000000;
assign F[56][19] = 9'b100000000;
assign F[56][20] = 9'b100000000;
assign F[56][21] = 9'b100000000;
assign F[56][22] = 9'b100000000;
assign F[57][3] = 9'b100000000;
assign F[57][4] = 9'b100000000;
assign F[57][5] = 9'b100000000;
assign F[57][6] = 9'b100000000;
assign F[57][7] = 9'b100000000;
assign F[57][8] = 9'b100000000;
assign F[57][9] = 9'b100000000;
assign F[57][10] = 9'b100100100;
assign F[57][11] = 9'b100000100;
assign F[57][12] = 9'b100000100;
assign F[57][13] = 9'b100000100;
assign F[57][14] = 9'b100000100;
assign F[57][15] = 9'b100100100;
assign F[57][16] = 9'b100100100;
assign F[57][17] = 9'b100000000;
assign F[57][18] = 9'b100000000;
assign F[57][19] = 9'b100000000;
assign F[57][20] = 9'b100000000;
assign F[57][21] = 9'b100000000;
assign F[57][22] = 9'b100000000;
assign F[58][3] = 9'b100000000;
assign F[58][4] = 9'b100000000;
assign F[58][5] = 9'b100000000;
assign F[58][6] = 9'b100000000;
assign F[58][7] = 9'b100000000;
assign F[58][8] = 9'b100000000;
assign F[58][10] = 9'b100000000;
assign F[58][11] = 9'b100000100;
assign F[58][12] = 9'b100000100;
assign F[58][13] = 9'b100000100;
assign F[58][14] = 9'b100000100;
assign F[58][15] = 9'b100100000;
assign F[58][16] = 9'b100000000;
assign F[58][17] = 9'b100000000;
assign F[58][18] = 9'b100000000;
assign F[58][19] = 9'b100000000;
assign F[58][20] = 9'b100000000;
assign F[58][21] = 9'b100000000;
assign F[58][22] = 9'b100000000;
assign F[59][3] = 9'b100000000;
assign F[59][4] = 9'b100000000;
assign F[59][5] = 9'b100000000;
assign F[59][6] = 9'b100000000;
assign F[59][7] = 9'b100000000;
assign F[59][8] = 9'b100000000;
assign F[59][9] = 9'b100000000;
assign F[59][10] = 9'b100000000;
assign F[59][15] = 9'b100000000;
assign F[59][16] = 9'b100000000;
assign F[59][17] = 9'b100000000;
assign F[59][18] = 9'b100000000;
assign F[59][19] = 9'b100000000;
assign F[59][20] = 9'b100000000;
assign F[59][21] = 9'b100000000;
assign F[59][22] = 9'b100000000;
assign F[60][4] = 9'b100000000;
assign F[60][5] = 9'b100000000;
assign F[60][6] = 9'b100100000;
assign F[60][7] = 9'b100000100;
assign F[60][8] = 9'b100000100;
assign F[60][9] = 9'b100000100;
assign F[60][10] = 9'b100000100;
assign F[60][11] = 9'b100000100;
assign F[60][12] = 9'b100000100;
assign F[60][13] = 9'b100000100;
assign F[60][14] = 9'b100000100;
assign F[60][15] = 9'b100000100;
assign F[60][16] = 9'b100000100;
assign F[60][17] = 9'b100000100;
assign F[60][18] = 9'b100000100;
assign F[60][19] = 9'b100100100;
assign F[60][20] = 9'b100000000;
assign F[60][21] = 9'b100000000;
assign F[60][22] = 9'b100000000;
assign F[61][6] = 9'b100100100;
assign F[61][7] = 9'b100000100;
assign F[61][8] = 9'b100000100;
assign F[61][9] = 9'b100000100;
assign F[61][10] = 9'b100000100;
assign F[61][11] = 9'b100000100;
assign F[61][12] = 9'b100000100;
assign F[61][13] = 9'b100000100;
assign F[61][14] = 9'b100000100;
assign F[61][15] = 9'b100000100;
assign F[61][16] = 9'b100000100;
assign F[61][17] = 9'b100000100;
assign F[61][18] = 9'b100000100;
assign F[61][19] = 9'b100100100;
assign F[62][6] = 9'b100100100;
assign F[62][7] = 9'b100100100;
assign F[62][8] = 9'b100000100;
assign F[62][9] = 9'b100000000;
assign F[62][10] = 9'b100000000;
assign F[62][11] = 9'b100000000;
assign F[62][12] = 9'b100000000;
assign F[62][13] = 9'b100000000;
assign F[62][14] = 9'b100000000;
assign F[62][15] = 9'b100000000;
assign F[62][16] = 9'b100000000;
assign F[62][17] = 9'b100000100;
assign F[62][18] = 9'b100000100;
assign F[62][19] = 9'b100100100;
assign F[63][6] = 9'b100100100;
assign F[63][7] = 9'b100000100;
assign F[63][8] = 9'b100101001;
assign F[63][9] = 9'b101101101;
assign F[63][10] = 9'b101101101;
assign F[63][11] = 9'b101101101;
assign F[63][12] = 9'b101101101;
assign F[63][13] = 9'b101101101;
assign F[63][14] = 9'b101101101;
assign F[63][15] = 9'b101101101;
assign F[63][16] = 9'b101101101;
assign F[63][17] = 9'b100101001;
assign F[63][18] = 9'b100000100;
assign F[63][19] = 9'b100100100;
assign F[64][6] = 9'b100100100;
assign F[64][7] = 9'b100000000;
assign F[64][8] = 9'b110010110;
assign F[64][9] = 9'b111111111;
assign F[64][10] = 9'b111111111;
assign F[64][11] = 9'b111111111;
assign F[64][12] = 9'b111111111;
assign F[64][13] = 9'b111111111;
assign F[64][14] = 9'b111111111;
assign F[64][15] = 9'b111111111;
assign F[64][16] = 9'b111111111;
assign F[64][17] = 9'b110010111;
assign F[64][18] = 9'b100000000;
assign F[64][19] = 9'b100100100;
assign F[65][6] = 9'b100100100;
assign F[65][7] = 9'b100000100;
assign F[65][8] = 9'b100101001;
assign F[65][9] = 9'b101001101;
assign F[65][10] = 9'b101001101;
assign F[65][11] = 9'b101001101;
assign F[65][12] = 9'b101001101;
assign F[65][13] = 9'b101001101;
assign F[65][14] = 9'b101001101;
assign F[65][15] = 9'b101001101;
assign F[65][16] = 9'b101001101;
assign F[65][17] = 9'b100101001;
assign F[65][18] = 9'b100000100;
assign F[65][19] = 9'b100100100;
//Total de Lineas = 867
endmodule


