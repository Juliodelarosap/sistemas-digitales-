`timescale 1ns / 1ps
module pantalla_de_inicio (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (F[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= F[vcount- posy][hcount- posx][7:5];
				green <= F[vcount- posy][hcount- posx][4:2];
            blue 	<= F[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 200;
parameter RESOLUCION_Y = 300;
wire [8:0] F[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign F[118][37] = 9'b111111100;
assign F[118][38] = 9'b110111100;
assign F[118][39] = 9'b110011100;
assign F[118][40] = 9'b110011100;
assign F[118][41] = 9'b110111100;
assign F[118][42] = 9'b110111100;
assign F[118][43] = 9'b110111100;
assign F[118][44] = 9'b110111100;
assign F[118][45] = 9'b110111100;
assign F[118][46] = 9'b110111100;
assign F[118][47] = 9'b110111100;
assign F[118][48] = 9'b110111100;
assign F[118][49] = 9'b110111100;
assign F[118][50] = 9'b110111100;
assign F[118][51] = 9'b110111100;
assign F[118][53] = 9'b101010001;
assign F[118][54] = 9'b100110100;
assign F[118][55] = 9'b100110101;
assign F[118][56] = 9'b100110001;
assign F[118][57] = 9'b100110001;
assign F[118][58] = 9'b100110001;
assign F[118][59] = 9'b100110001;
assign F[118][60] = 9'b100110101;
assign F[118][61] = 9'b100110101;
assign F[118][65] = 9'b100110001;
assign F[118][66] = 9'b100110101;
assign F[118][67] = 9'b100110001;
assign F[118][68] = 9'b100110001;
assign F[118][69] = 9'b100110001;
assign F[118][70] = 9'b100110000;
assign F[118][71] = 9'b100110001;
assign F[118][72] = 9'b110111111;
assign F[118][73] = 9'b111111100;
assign F[118][74] = 9'b110111100;
assign F[118][75] = 9'b110011100;
assign F[118][76] = 9'b110111100;
assign F[118][77] = 9'b110111100;
assign F[118][78] = 9'b110111100;
assign F[118][79] = 9'b110111100;
assign F[118][80] = 9'b110111100;
assign F[118][81] = 9'b110111100;
assign F[118][82] = 9'b110111100;
assign F[118][83] = 9'b110111100;
assign F[118][84] = 9'b110111100;
assign F[118][85] = 9'b110111100;
assign F[118][86] = 9'b110111101;
assign F[118][93] = 9'b101010101;
assign F[118][94] = 9'b100110101;
assign F[118][95] = 9'b100110101;
assign F[118][96] = 9'b100010000;
assign F[118][97] = 9'b100010000;
assign F[118][98] = 9'b100010000;
assign F[118][99] = 9'b100010000;
assign F[118][100] = 9'b100110001;
assign F[118][101] = 9'b100110001;
assign F[118][102] = 9'b100110101;
assign F[118][103] = 9'b100110001;
assign F[118][104] = 9'b101010101;
assign F[118][110] = 9'b110111100;
assign F[118][111] = 9'b110111100;
assign F[118][112] = 9'b110111100;
assign F[118][113] = 9'b110111100;
assign F[118][114] = 9'b110111100;
assign F[118][115] = 9'b110111100;
assign F[118][116] = 9'b110111100;
assign F[118][117] = 9'b110111100;
assign F[118][127] = 9'b101110101;
assign F[118][128] = 9'b100110000;
assign F[118][129] = 9'b100110001;
assign F[118][130] = 9'b100110001;
assign F[118][131] = 9'b100110001;
assign F[118][132] = 9'b100110001;
assign F[118][133] = 9'b100110100;
assign F[118][134] = 9'b100110001;
assign F[118][139] = 9'b111111101;
assign F[118][140] = 9'b110111100;
assign F[118][141] = 9'b110111100;
assign F[118][142] = 9'b110111100;
assign F[118][143] = 9'b110111100;
assign F[118][144] = 9'b110111100;
assign F[118][145] = 9'b110111100;
assign F[118][146] = 9'b110111101;
assign F[118][150] = 9'b111111100;
assign F[118][151] = 9'b110111100;
assign F[118][152] = 9'b110111100;
assign F[118][153] = 9'b110111100;
assign F[118][154] = 9'b110111101;
assign F[119][37] = 9'b111111100;
assign F[119][38] = 9'b110111100;
assign F[119][39] = 9'b110111100;
assign F[119][40] = 9'b110111100;
assign F[119][41] = 9'b110111100;
assign F[119][42] = 9'b110111100;
assign F[119][43] = 9'b110111100;
assign F[119][44] = 9'b110111100;
assign F[119][45] = 9'b110111100;
assign F[119][46] = 9'b110111100;
assign F[119][47] = 9'b110111100;
assign F[119][48] = 9'b110111100;
assign F[119][49] = 9'b110111100;
assign F[119][50] = 9'b111111100;
assign F[119][51] = 9'b110111100;
assign F[119][53] = 9'b101010000;
assign F[119][54] = 9'b100110100;
assign F[119][55] = 9'b100010100;
assign F[119][56] = 9'b100010100;
assign F[119][57] = 9'b100010100;
assign F[119][58] = 9'b100010100;
assign F[119][59] = 9'b100010100;
assign F[119][60] = 9'b100010100;
assign F[119][61] = 9'b100010101;
assign F[119][65] = 9'b100010100;
assign F[119][66] = 9'b100010100;
assign F[119][67] = 9'b100010100;
assign F[119][68] = 9'b100010100;
assign F[119][69] = 9'b100010100;
assign F[119][70] = 9'b100010100;
assign F[119][71] = 9'b100110101;
assign F[119][72] = 9'b111111111;
assign F[119][73] = 9'b111111100;
assign F[119][74] = 9'b110111100;
assign F[119][75] = 9'b110111100;
assign F[119][76] = 9'b110111100;
assign F[119][77] = 9'b110111100;
assign F[119][78] = 9'b110111100;
assign F[119][79] = 9'b110111100;
assign F[119][80] = 9'b110111100;
assign F[119][81] = 9'b110111100;
assign F[119][82] = 9'b110111100;
assign F[119][83] = 9'b110111100;
assign F[119][84] = 9'b110111100;
assign F[119][85] = 9'b110111100;
assign F[119][86] = 9'b110111101;
assign F[119][93] = 9'b100110100;
assign F[119][94] = 9'b100010100;
assign F[119][95] = 9'b100010000;
assign F[119][96] = 9'b100010000;
assign F[119][97] = 9'b100010000;
assign F[119][98] = 9'b100010000;
assign F[119][99] = 9'b100010000;
assign F[119][100] = 9'b100010000;
assign F[119][101] = 9'b100010000;
assign F[119][102] = 9'b100010100;
assign F[119][103] = 9'b100010100;
assign F[119][104] = 9'b100010100;
assign F[119][105] = 9'b100110001;
assign F[119][106] = 9'b101010101;
assign F[119][110] = 9'b111111100;
assign F[119][111] = 9'b111111100;
assign F[119][112] = 9'b110111100;
assign F[119][113] = 9'b110111100;
assign F[119][114] = 9'b110111100;
assign F[119][115] = 9'b110111100;
assign F[119][116] = 9'b110111100;
assign F[119][117] = 9'b110111100;
assign F[119][118] = 9'b110011101;
assign F[119][127] = 9'b101010000;
assign F[119][128] = 9'b100010100;
assign F[119][129] = 9'b100110100;
assign F[119][130] = 9'b100010100;
assign F[119][131] = 9'b100010100;
assign F[119][132] = 9'b100010100;
assign F[119][133] = 9'b100010100;
assign F[119][134] = 9'b100110101;
assign F[119][135] = 9'b101011110;
assign F[119][139] = 9'b111111101;
assign F[119][140] = 9'b111111100;
assign F[119][141] = 9'b110111100;
assign F[119][142] = 9'b110111100;
assign F[119][143] = 9'b110111100;
assign F[119][144] = 9'b110111100;
assign F[119][145] = 9'b110111100;
assign F[119][146] = 9'b110011100;
assign F[119][147] = 9'b110111101;
assign F[119][150] = 9'b111111100;
assign F[119][151] = 9'b111111100;
assign F[119][152] = 9'b110111100;
assign F[119][153] = 9'b110111100;
assign F[119][154] = 9'b110011100;
assign F[120][37] = 9'b111111100;
assign F[120][38] = 9'b110011100;
assign F[120][39] = 9'b110111100;
assign F[120][40] = 9'b110011100;
assign F[120][41] = 9'b110011100;
assign F[120][42] = 9'b110011100;
assign F[120][43] = 9'b110011100;
assign F[120][44] = 9'b110011100;
assign F[120][45] = 9'b110011100;
assign F[120][46] = 9'b110011100;
assign F[120][47] = 9'b110011100;
assign F[120][48] = 9'b110011100;
assign F[120][49] = 9'b110011100;
assign F[120][50] = 9'b110111100;
assign F[120][51] = 9'b110111100;
assign F[120][53] = 9'b101010000;
assign F[120][54] = 9'b100110100;
assign F[120][55] = 9'b100010000;
assign F[120][56] = 9'b100010000;
assign F[120][57] = 9'b100010000;
assign F[120][58] = 9'b100010000;
assign F[120][59] = 9'b100010000;
assign F[120][60] = 9'b100010100;
assign F[120][61] = 9'b100110101;
assign F[120][65] = 9'b100110000;
assign F[120][66] = 9'b100010000;
assign F[120][67] = 9'b100010000;
assign F[120][68] = 9'b100010000;
assign F[120][69] = 9'b100010000;
assign F[120][70] = 9'b100010000;
assign F[120][71] = 9'b100110001;
assign F[120][72] = 9'b111111111;
assign F[120][73] = 9'b111111100;
assign F[120][74] = 9'b110111100;
assign F[120][75] = 9'b110011100;
assign F[120][76] = 9'b110011100;
assign F[120][77] = 9'b110011100;
assign F[120][78] = 9'b110011100;
assign F[120][79] = 9'b110011100;
assign F[120][80] = 9'b110011100;
assign F[120][81] = 9'b110011100;
assign F[120][82] = 9'b110011100;
assign F[120][83] = 9'b110011100;
assign F[120][84] = 9'b110011100;
assign F[120][85] = 9'b110111100;
assign F[120][86] = 9'b110111101;
assign F[120][93] = 9'b101010000;
assign F[120][94] = 9'b100010000;
assign F[120][95] = 9'b100010000;
assign F[120][96] = 9'b100010000;
assign F[120][97] = 9'b100010000;
assign F[120][98] = 9'b100010000;
assign F[120][99] = 9'b100010000;
assign F[120][100] = 9'b100010000;
assign F[120][101] = 9'b100010000;
assign F[120][102] = 9'b100010000;
assign F[120][103] = 9'b100010000;
assign F[120][104] = 9'b100010000;
assign F[120][105] = 9'b100110000;
assign F[120][106] = 9'b100010001;
assign F[120][107] = 9'b100110001;
assign F[120][110] = 9'b111111100;
assign F[120][111] = 9'b110111100;
assign F[120][112] = 9'b110011100;
assign F[120][113] = 9'b110111100;
assign F[120][114] = 9'b110011100;
assign F[120][115] = 9'b110011100;
assign F[120][116] = 9'b110111100;
assign F[120][117] = 9'b110111100;
assign F[120][118] = 9'b110111101;
assign F[120][127] = 9'b100110000;
assign F[120][128] = 9'b100010100;
assign F[120][129] = 9'b100110000;
assign F[120][130] = 9'b100010000;
assign F[120][131] = 9'b100010000;
assign F[120][132] = 9'b100010000;
assign F[120][133] = 9'b100010000;
assign F[120][134] = 9'b100010100;
assign F[120][135] = 9'b100111110;
assign F[120][139] = 9'b111111101;
assign F[120][140] = 9'b111111100;
assign F[120][141] = 9'b110011100;
assign F[120][142] = 9'b110011100;
assign F[120][143] = 9'b110011100;
assign F[120][144] = 9'b110011100;
assign F[120][145] = 9'b110111100;
assign F[120][146] = 9'b110111100;
assign F[120][147] = 9'b110011100;
assign F[120][148] = 9'b110111101;
assign F[120][150] = 9'b111111100;
assign F[120][151] = 9'b110111100;
assign F[120][152] = 9'b110011100;
assign F[120][153] = 9'b110111100;
assign F[120][154] = 9'b110111101;
assign F[121][37] = 9'b111111100;
assign F[121][38] = 9'b110011100;
assign F[121][39] = 9'b110111100;
assign F[121][40] = 9'b110011100;
assign F[121][41] = 9'b110011100;
assign F[121][42] = 9'b110011100;
assign F[121][43] = 9'b110011100;
assign F[121][44] = 9'b110011100;
assign F[121][45] = 9'b110011100;
assign F[121][46] = 9'b110011100;
assign F[121][47] = 9'b110011100;
assign F[121][48] = 9'b110011100;
assign F[121][49] = 9'b110011100;
assign F[121][50] = 9'b110111100;
assign F[121][51] = 9'b110111100;
assign F[121][53] = 9'b101010100;
assign F[121][54] = 9'b100110100;
assign F[121][55] = 9'b100010000;
assign F[121][56] = 9'b100010000;
assign F[121][57] = 9'b100010000;
assign F[121][58] = 9'b100010000;
assign F[121][59] = 9'b100010000;
assign F[121][60] = 9'b100010101;
assign F[121][61] = 9'b100110101;
assign F[121][65] = 9'b100110000;
assign F[121][66] = 9'b100010000;
assign F[121][67] = 9'b100010000;
assign F[121][68] = 9'b100010000;
assign F[121][69] = 9'b100010000;
assign F[121][70] = 9'b100010000;
assign F[121][71] = 9'b100110101;
assign F[121][72] = 9'b111111111;
assign F[121][73] = 9'b111111101;
assign F[121][74] = 9'b110111100;
assign F[121][75] = 9'b110011100;
assign F[121][76] = 9'b110011100;
assign F[121][77] = 9'b110011100;
assign F[121][78] = 9'b110011100;
assign F[121][79] = 9'b110011100;
assign F[121][80] = 9'b110011100;
assign F[121][81] = 9'b110011100;
assign F[121][82] = 9'b110011100;
assign F[121][83] = 9'b110011100;
assign F[121][84] = 9'b110011100;
assign F[121][85] = 9'b110111100;
assign F[121][86] = 9'b110111101;
assign F[121][93] = 9'b101010101;
assign F[121][94] = 9'b100010000;
assign F[121][95] = 9'b100010000;
assign F[121][96] = 9'b100010000;
assign F[121][97] = 9'b100010000;
assign F[121][98] = 9'b100010000;
assign F[121][99] = 9'b100010000;
assign F[121][100] = 9'b100010000;
assign F[121][101] = 9'b100010000;
assign F[121][102] = 9'b100010000;
assign F[121][103] = 9'b100010000;
assign F[121][104] = 9'b100010000;
assign F[121][105] = 9'b100110000;
assign F[121][106] = 9'b100010100;
assign F[121][107] = 9'b100010001;
assign F[121][108] = 9'b101010110;
assign F[121][110] = 9'b111111100;
assign F[121][111] = 9'b110111100;
assign F[121][112] = 9'b110011100;
assign F[121][113] = 9'b110111100;
assign F[121][114] = 9'b110011100;
assign F[121][115] = 9'b110011100;
assign F[121][116] = 9'b110111100;
assign F[121][117] = 9'b110111100;
assign F[121][118] = 9'b110111101;
assign F[121][126] = 9'b110011101;
assign F[121][127] = 9'b100110000;
assign F[121][128] = 9'b100010000;
assign F[121][129] = 9'b100010000;
assign F[121][130] = 9'b100110000;
assign F[121][131] = 9'b100010000;
assign F[121][132] = 9'b100010000;
assign F[121][133] = 9'b100010000;
assign F[121][134] = 9'b100010100;
assign F[121][135] = 9'b100110101;
assign F[121][139] = 9'b111111101;
assign F[121][140] = 9'b111111100;
assign F[121][141] = 9'b110111100;
assign F[121][142] = 9'b110011100;
assign F[121][143] = 9'b110011100;
assign F[121][144] = 9'b110111100;
assign F[121][145] = 9'b110111100;
assign F[121][146] = 9'b110011100;
assign F[121][147] = 9'b110011100;
assign F[121][148] = 9'b110011100;
assign F[121][149] = 9'b110111101;
assign F[121][150] = 9'b111111100;
assign F[121][151] = 9'b110111100;
assign F[121][152] = 9'b110011100;
assign F[121][153] = 9'b110111100;
assign F[121][154] = 9'b110111101;
assign F[122][37] = 9'b111111100;
assign F[122][38] = 9'b110111100;
assign F[122][39] = 9'b110111100;
assign F[122][40] = 9'b110011100;
assign F[122][41] = 9'b110011100;
assign F[122][42] = 9'b110011100;
assign F[122][43] = 9'b110011100;
assign F[122][44] = 9'b110011100;
assign F[122][45] = 9'b110011100;
assign F[122][46] = 9'b110011100;
assign F[122][47] = 9'b110011100;
assign F[122][48] = 9'b110111100;
assign F[122][49] = 9'b110111100;
assign F[122][50] = 9'b110111100;
assign F[122][51] = 9'b110011100;
assign F[122][53] = 9'b101110100;
assign F[122][54] = 9'b100110100;
assign F[122][55] = 9'b100010000;
assign F[122][56] = 9'b100010000;
assign F[122][57] = 9'b100010000;
assign F[122][58] = 9'b100010000;
assign F[122][59] = 9'b100010000;
assign F[122][60] = 9'b100110101;
assign F[122][61] = 9'b100110101;
assign F[122][65] = 9'b100110000;
assign F[122][66] = 9'b100010000;
assign F[122][67] = 9'b100010000;
assign F[122][68] = 9'b100010000;
assign F[122][69] = 9'b100010000;
assign F[122][70] = 9'b100010000;
assign F[122][71] = 9'b100110101;
assign F[122][72] = 9'b111111111;
assign F[122][73] = 9'b111111101;
assign F[122][74] = 9'b110111100;
assign F[122][75] = 9'b110011100;
assign F[122][76] = 9'b110011100;
assign F[122][77] = 9'b110011100;
assign F[122][78] = 9'b110011100;
assign F[122][79] = 9'b110011100;
assign F[122][80] = 9'b110011100;
assign F[122][81] = 9'b110011100;
assign F[122][82] = 9'b110111100;
assign F[122][83] = 9'b110111100;
assign F[122][84] = 9'b110011100;
assign F[122][85] = 9'b110011100;
assign F[122][86] = 9'b110111101;
assign F[122][93] = 9'b101010100;
assign F[122][94] = 9'b100010100;
assign F[122][95] = 9'b100010000;
assign F[122][96] = 9'b100010000;
assign F[122][97] = 9'b100010000;
assign F[122][98] = 9'b100010000;
assign F[122][99] = 9'b100010000;
assign F[122][100] = 9'b100010000;
assign F[122][101] = 9'b100010000;
assign F[122][102] = 9'b100010000;
assign F[122][103] = 9'b100010000;
assign F[122][104] = 9'b100010000;
assign F[122][105] = 9'b100010001;
assign F[122][106] = 9'b100010000;
assign F[122][107] = 9'b100010100;
assign F[122][108] = 9'b100110101;
assign F[122][110] = 9'b111111100;
assign F[122][111] = 9'b110111100;
assign F[122][112] = 9'b110011100;
assign F[122][113] = 9'b110011100;
assign F[122][114] = 9'b110011100;
assign F[122][115] = 9'b110011100;
assign F[122][116] = 9'b110011100;
assign F[122][117] = 9'b110111100;
assign F[122][118] = 9'b110111101;
assign F[122][126] = 9'b101110101;
assign F[122][127] = 9'b100110100;
assign F[122][128] = 9'b100010000;
assign F[122][129] = 9'b100110000;
assign F[122][130] = 9'b100010000;
assign F[122][131] = 9'b100010000;
assign F[122][132] = 9'b100010000;
assign F[122][133] = 9'b100010000;
assign F[122][134] = 9'b100010000;
assign F[122][135] = 9'b100110101;
assign F[122][140] = 9'b111111100;
assign F[122][141] = 9'b110111100;
assign F[122][142] = 9'b110011100;
assign F[122][143] = 9'b110011100;
assign F[122][144] = 9'b110111100;
assign F[122][145] = 9'b110011100;
assign F[122][146] = 9'b110011100;
assign F[122][147] = 9'b110011100;
assign F[122][148] = 9'b110111100;
assign F[122][149] = 9'b110111100;
assign F[122][150] = 9'b110111100;
assign F[122][151] = 9'b110011100;
assign F[122][152] = 9'b110011100;
assign F[122][153] = 9'b110111100;
assign F[122][154] = 9'b110111101;
assign F[123][37] = 9'b111111100;
assign F[123][38] = 9'b110111100;
assign F[123][39] = 9'b110011100;
assign F[123][40] = 9'b110111100;
assign F[123][41] = 9'b110011100;
assign F[123][42] = 9'b110011100;
assign F[123][43] = 9'b110011100;
assign F[123][44] = 9'b110011100;
assign F[123][45] = 9'b110011100;
assign F[123][46] = 9'b110011100;
assign F[123][47] = 9'b110011100;
assign F[123][48] = 9'b110011100;
assign F[123][49] = 9'b110011100;
assign F[123][50] = 9'b110111100;
assign F[123][51] = 9'b110111100;
assign F[123][53] = 9'b101110101;
assign F[123][54] = 9'b100110100;
assign F[123][55] = 9'b100010000;
assign F[123][56] = 9'b100010000;
assign F[123][57] = 9'b100010000;
assign F[123][58] = 9'b100010000;
assign F[123][59] = 9'b100010000;
assign F[123][60] = 9'b100010101;
assign F[123][61] = 9'b100110101;
assign F[123][65] = 9'b100110000;
assign F[123][66] = 9'b100010000;
assign F[123][67] = 9'b100010000;
assign F[123][68] = 9'b100010000;
assign F[123][69] = 9'b100010000;
assign F[123][70] = 9'b100010000;
assign F[123][71] = 9'b100110101;
assign F[123][72] = 9'b111111111;
assign F[123][73] = 9'b111111101;
assign F[123][74] = 9'b110111100;
assign F[123][75] = 9'b110011100;
assign F[123][76] = 9'b110011100;
assign F[123][77] = 9'b110011100;
assign F[123][78] = 9'b110011100;
assign F[123][79] = 9'b110011100;
assign F[123][80] = 9'b110011100;
assign F[123][81] = 9'b110011100;
assign F[123][82] = 9'b110011100;
assign F[123][83] = 9'b110111100;
assign F[123][84] = 9'b110111100;
assign F[123][85] = 9'b110011100;
assign F[123][93] = 9'b100110000;
assign F[123][94] = 9'b100010100;
assign F[123][95] = 9'b100110000;
assign F[123][96] = 9'b100010000;
assign F[123][97] = 9'b100010000;
assign F[123][98] = 9'b100010000;
assign F[123][99] = 9'b100010000;
assign F[123][100] = 9'b100010001;
assign F[123][101] = 9'b101010101;
assign F[123][102] = 9'b101010101;
assign F[123][103] = 9'b100110000;
assign F[123][104] = 9'b100010000;
assign F[123][105] = 9'b100010000;
assign F[123][106] = 9'b100010000;
assign F[123][107] = 9'b100010000;
assign F[123][108] = 9'b100110001;
assign F[123][110] = 9'b111111100;
assign F[123][111] = 9'b110111100;
assign F[123][112] = 9'b110011100;
assign F[123][113] = 9'b110011100;
assign F[123][114] = 9'b110011100;
assign F[123][115] = 9'b110111100;
assign F[123][116] = 9'b110011100;
assign F[123][117] = 9'b110111100;
assign F[123][118] = 9'b110111110;
assign F[123][126] = 9'b101010000;
assign F[123][127] = 9'b100110100;
assign F[123][128] = 9'b100010000;
assign F[123][129] = 9'b100110000;
assign F[123][130] = 9'b100010000;
assign F[123][131] = 9'b100010000;
assign F[123][132] = 9'b100010000;
assign F[123][133] = 9'b100010000;
assign F[123][134] = 9'b100010000;
assign F[123][135] = 9'b100110101;
assign F[123][136] = 9'b101011111;
assign F[123][140] = 9'b111111100;
assign F[123][141] = 9'b110111100;
assign F[123][142] = 9'b110011100;
assign F[123][143] = 9'b110011100;
assign F[123][144] = 9'b110011100;
assign F[123][145] = 9'b110011100;
assign F[123][146] = 9'b110011100;
assign F[123][147] = 9'b110011100;
assign F[123][148] = 9'b110011100;
assign F[123][149] = 9'b110011100;
assign F[123][150] = 9'b110011100;
assign F[123][151] = 9'b110011100;
assign F[123][152] = 9'b110011100;
assign F[123][153] = 9'b110111100;
assign F[123][154] = 9'b110111101;
assign F[124][41] = 9'b110111100;
assign F[124][42] = 9'b110111100;
assign F[124][43] = 9'b110011100;
assign F[124][44] = 9'b110011100;
assign F[124][45] = 9'b110111100;
assign F[124][46] = 9'b110111100;
assign F[124][47] = 9'b110011100;
assign F[124][53] = 9'b110011101;
assign F[124][54] = 9'b100110100;
assign F[124][55] = 9'b100010000;
assign F[124][56] = 9'b100010000;
assign F[124][57] = 9'b100010000;
assign F[124][58] = 9'b100010000;
assign F[124][59] = 9'b100010000;
assign F[124][60] = 9'b100010101;
assign F[124][61] = 9'b100111110;
assign F[124][65] = 9'b100110000;
assign F[124][66] = 9'b100010000;
assign F[124][67] = 9'b100010000;
assign F[124][68] = 9'b100010000;
assign F[124][69] = 9'b100010000;
assign F[124][70] = 9'b100010000;
assign F[124][71] = 9'b101011101;
assign F[124][72] = 9'b111111111;
assign F[124][73] = 9'b111111101;
assign F[124][74] = 9'b110111100;
assign F[124][75] = 9'b110011100;
assign F[124][76] = 9'b110011100;
assign F[124][77] = 9'b110011100;
assign F[124][78] = 9'b110011100;
assign F[124][79] = 9'b110011100;
assign F[124][80] = 9'b110111100;
assign F[124][81] = 9'b110111101;
assign F[124][93] = 9'b100110000;
assign F[124][94] = 9'b100010100;
assign F[124][95] = 9'b100010000;
assign F[124][96] = 9'b100010000;
assign F[124][97] = 9'b100010000;
assign F[124][98] = 9'b100010000;
assign F[124][99] = 9'b100010000;
assign F[124][100] = 9'b100110110;
assign F[124][101] = 9'b111111111;
assign F[124][102] = 9'b111111111;
assign F[124][103] = 9'b111111110;
assign F[124][104] = 9'b101010001;
assign F[124][105] = 9'b100010000;
assign F[124][106] = 9'b100010000;
assign F[124][107] = 9'b100010000;
assign F[124][108] = 9'b100110101;
assign F[124][110] = 9'b111111101;
assign F[124][111] = 9'b110111100;
assign F[124][112] = 9'b110011100;
assign F[124][113] = 9'b110011100;
assign F[124][114] = 9'b110011100;
assign F[124][115] = 9'b110111100;
assign F[124][116] = 9'b110011100;
assign F[124][117] = 9'b110111100;
assign F[124][118] = 9'b110111110;
assign F[124][126] = 9'b101010000;
assign F[124][127] = 9'b100010000;
assign F[124][128] = 9'b100010000;
assign F[124][129] = 9'b100010000;
assign F[124][130] = 9'b100010000;
assign F[124][131] = 9'b100010000;
assign F[124][132] = 9'b100010000;
assign F[124][133] = 9'b100010000;
assign F[124][134] = 9'b100010000;
assign F[124][135] = 9'b100010100;
assign F[124][136] = 9'b100110001;
assign F[124][140] = 9'b111111100;
assign F[124][141] = 9'b110111100;
assign F[124][142] = 9'b110011100;
assign F[124][143] = 9'b110011100;
assign F[124][144] = 9'b110011100;
assign F[124][145] = 9'b110011100;
assign F[124][146] = 9'b110011100;
assign F[124][147] = 9'b110011100;
assign F[124][148] = 9'b110011100;
assign F[124][149] = 9'b110011100;
assign F[124][150] = 9'b110011100;
assign F[124][151] = 9'b110011100;
assign F[124][152] = 9'b110011100;
assign F[124][153] = 9'b110111100;
assign F[124][154] = 9'b110111101;
assign F[125][41] = 9'b111111100;
assign F[125][42] = 9'b110111100;
assign F[125][43] = 9'b110011100;
assign F[125][44] = 9'b110011100;
assign F[125][45] = 9'b110011100;
assign F[125][46] = 9'b110011100;
assign F[125][47] = 9'b110011101;
assign F[125][53] = 9'b110011101;
assign F[125][54] = 9'b100110100;
assign F[125][55] = 9'b100010000;
assign F[125][56] = 9'b100010000;
assign F[125][57] = 9'b100010000;
assign F[125][58] = 9'b100010000;
assign F[125][59] = 9'b100010000;
assign F[125][60] = 9'b100110101;
assign F[125][61] = 9'b100111111;
assign F[125][65] = 9'b100110000;
assign F[125][66] = 9'b100010000;
assign F[125][67] = 9'b100010000;
assign F[125][68] = 9'b100010000;
assign F[125][69] = 9'b100010000;
assign F[125][70] = 9'b100010000;
assign F[125][71] = 9'b101011101;
assign F[125][72] = 9'b111111111;
assign F[125][73] = 9'b111111101;
assign F[125][74] = 9'b110111100;
assign F[125][75] = 9'b110011100;
assign F[125][76] = 9'b110011100;
assign F[125][77] = 9'b110011100;
assign F[125][78] = 9'b110011100;
assign F[125][79] = 9'b110011100;
assign F[125][80] = 9'b110011100;
assign F[125][81] = 9'b110111100;
assign F[125][82] = 9'b110111100;
assign F[125][83] = 9'b110111100;
assign F[125][84] = 9'b110111100;
assign F[125][85] = 9'b110111101;
assign F[125][93] = 9'b100110001;
assign F[125][94] = 9'b100010100;
assign F[125][95] = 9'b100010000;
assign F[125][96] = 9'b100010000;
assign F[125][97] = 9'b100010000;
assign F[125][98] = 9'b100010000;
assign F[125][99] = 9'b100010000;
assign F[125][100] = 9'b100111110;
assign F[125][101] = 9'b111111111;
assign F[125][102] = 9'b111111111;
assign F[125][103] = 9'b111111110;
assign F[125][104] = 9'b101010100;
assign F[125][105] = 9'b100010000;
assign F[125][106] = 9'b100010000;
assign F[125][107] = 9'b100010000;
assign F[125][108] = 9'b100110101;
assign F[125][110] = 9'b111111101;
assign F[125][111] = 9'b110111100;
assign F[125][112] = 9'b110011100;
assign F[125][113] = 9'b110011100;
assign F[125][114] = 9'b110011100;
assign F[125][115] = 9'b110111100;
assign F[125][116] = 9'b110111100;
assign F[125][117] = 9'b110011100;
assign F[125][125] = 9'b110010101;
assign F[125][126] = 9'b100110000;
assign F[125][127] = 9'b100010000;
assign F[125][128] = 9'b100010000;
assign F[125][129] = 9'b100010000;
assign F[125][130] = 9'b100010000;
assign F[125][131] = 9'b100010000;
assign F[125][132] = 9'b100010000;
assign F[125][133] = 9'b100010000;
assign F[125][134] = 9'b100010000;
assign F[125][135] = 9'b100010100;
assign F[125][136] = 9'b100110001;
assign F[125][140] = 9'b111111100;
assign F[125][141] = 9'b110111100;
assign F[125][142] = 9'b110011100;
assign F[125][143] = 9'b110011100;
assign F[125][144] = 9'b110011100;
assign F[125][145] = 9'b110011100;
assign F[125][146] = 9'b110011100;
assign F[125][147] = 9'b110011100;
assign F[125][148] = 9'b110011100;
assign F[125][149] = 9'b110011100;
assign F[125][150] = 9'b110011100;
assign F[125][151] = 9'b110011100;
assign F[125][152] = 9'b110011100;
assign F[125][153] = 9'b110111100;
assign F[125][154] = 9'b110111101;
assign F[126][41] = 9'b111111100;
assign F[126][42] = 9'b110111100;
assign F[126][43] = 9'b110011100;
assign F[126][44] = 9'b110011100;
assign F[126][45] = 9'b110011100;
assign F[126][46] = 9'b110111100;
assign F[126][47] = 9'b110111101;
assign F[126][53] = 9'b111111101;
assign F[126][54] = 9'b100110100;
assign F[126][55] = 9'b100010000;
assign F[126][56] = 9'b100010000;
assign F[126][57] = 9'b100010000;
assign F[126][58] = 9'b100010000;
assign F[126][59] = 9'b100010000;
assign F[126][60] = 9'b100010101;
assign F[126][61] = 9'b100111110;
assign F[126][62] = 9'b101111110;
assign F[126][63] = 9'b110010101;
assign F[126][64] = 9'b101110101;
assign F[126][65] = 9'b100110000;
assign F[126][66] = 9'b100010000;
assign F[126][67] = 9'b100010000;
assign F[126][68] = 9'b100010000;
assign F[126][69] = 9'b100010000;
assign F[126][70] = 9'b100010000;
assign F[126][71] = 9'b101011110;
assign F[126][72] = 9'b111111111;
assign F[126][73] = 9'b111111101;
assign F[126][74] = 9'b110111100;
assign F[126][75] = 9'b110011100;
assign F[126][76] = 9'b110011100;
assign F[126][77] = 9'b110011100;
assign F[126][78] = 9'b110011100;
assign F[126][79] = 9'b110011100;
assign F[126][80] = 9'b110011100;
assign F[126][81] = 9'b110011100;
assign F[126][82] = 9'b110111100;
assign F[126][83] = 9'b110011100;
assign F[126][84] = 9'b110111100;
assign F[126][85] = 9'b110111101;
assign F[126][93] = 9'b100110100;
assign F[126][94] = 9'b100010101;
assign F[126][95] = 9'b100110000;
assign F[126][96] = 9'b100010000;
assign F[126][97] = 9'b100010000;
assign F[126][98] = 9'b100010000;
assign F[126][99] = 9'b100010000;
assign F[126][100] = 9'b100110101;
assign F[126][101] = 9'b110011111;
assign F[126][102] = 9'b110011101;
assign F[126][103] = 9'b101010101;
assign F[126][104] = 9'b100110000;
assign F[126][105] = 9'b100110000;
assign F[126][106] = 9'b100010100;
assign F[126][107] = 9'b100110101;
assign F[126][110] = 9'b111111101;
assign F[126][111] = 9'b111111100;
assign F[126][112] = 9'b110011100;
assign F[126][113] = 9'b110011100;
assign F[126][114] = 9'b110011100;
assign F[126][115] = 9'b110111100;
assign F[126][116] = 9'b110111100;
assign F[126][117] = 9'b110011100;
assign F[126][124] = 9'b111111101;
assign F[126][125] = 9'b110011101;
assign F[126][126] = 9'b100010000;
assign F[126][127] = 9'b100110000;
assign F[126][128] = 9'b100010001;
assign F[126][129] = 9'b101111101;
assign F[126][130] = 9'b101010100;
assign F[126][131] = 9'b100010000;
assign F[126][132] = 9'b100010000;
assign F[126][133] = 9'b100010000;
assign F[126][134] = 9'b100010000;
assign F[126][135] = 9'b100010000;
assign F[126][136] = 9'b100010001;
assign F[126][137] = 9'b101010110;
assign F[126][140] = 9'b111111101;
assign F[126][141] = 9'b110111100;
assign F[126][142] = 9'b110011100;
assign F[126][143] = 9'b110011100;
assign F[126][144] = 9'b110111100;
assign F[126][145] = 9'b110011100;
assign F[126][146] = 9'b110011100;
assign F[126][147] = 9'b110011100;
assign F[126][148] = 9'b110011100;
assign F[126][149] = 9'b110011100;
assign F[126][150] = 9'b110011100;
assign F[126][151] = 9'b110011100;
assign F[126][152] = 9'b110011100;
assign F[126][153] = 9'b110111100;
assign F[126][154] = 9'b111111110;
assign F[127][37] = 9'b110111100;
assign F[127][38] = 9'b110111100;
assign F[127][39] = 9'b110111100;
assign F[127][40] = 9'b110111100;
assign F[127][41] = 9'b110111100;
assign F[127][42] = 9'b110011100;
assign F[127][43] = 9'b110011100;
assign F[127][44] = 9'b110011100;
assign F[127][45] = 9'b110111100;
assign F[127][46] = 9'b110111100;
assign F[127][47] = 9'b110011100;
assign F[127][48] = 9'b110111100;
assign F[127][49] = 9'b110111100;
assign F[127][50] = 9'b110111100;
assign F[127][51] = 9'b110111100;
assign F[127][52] = 9'b101111100;
assign F[127][53] = 9'b101010000;
assign F[127][54] = 9'b100110100;
assign F[127][55] = 9'b100010000;
assign F[127][56] = 9'b100010000;
assign F[127][57] = 9'b100010000;
assign F[127][58] = 9'b100010000;
assign F[127][59] = 9'b100010000;
assign F[127][60] = 9'b100010000;
assign F[127][61] = 9'b100010000;
assign F[127][62] = 9'b100110101;
assign F[127][63] = 9'b100110001;
assign F[127][64] = 9'b100110101;
assign F[127][65] = 9'b100010000;
assign F[127][66] = 9'b100010000;
assign F[127][67] = 9'b100010000;
assign F[127][68] = 9'b100010000;
assign F[127][69] = 9'b100010000;
assign F[127][70] = 9'b100010000;
assign F[127][71] = 9'b100110101;
assign F[127][72] = 9'b110011101;
assign F[127][73] = 9'b111111101;
assign F[127][74] = 9'b110111100;
assign F[127][75] = 9'b110011100;
assign F[127][76] = 9'b110011100;
assign F[127][77] = 9'b110011100;
assign F[127][78] = 9'b110011100;
assign F[127][79] = 9'b110011100;
assign F[127][80] = 9'b110011100;
assign F[127][81] = 9'b110111100;
assign F[127][82] = 9'b110111100;
assign F[127][83] = 9'b110111100;
assign F[127][84] = 9'b110111100;
assign F[127][85] = 9'b110111101;
assign F[127][86] = 9'b110111100;
assign F[127][87] = 9'b110111100;
assign F[127][88] = 9'b110111100;
assign F[127][89] = 9'b110111100;
assign F[127][90] = 9'b110111100;
assign F[127][91] = 9'b110111100;
assign F[127][92] = 9'b101010100;
assign F[127][93] = 9'b100110000;
assign F[127][94] = 9'b100010000;
assign F[127][95] = 9'b100010000;
assign F[127][96] = 9'b100010000;
assign F[127][97] = 9'b100010000;
assign F[127][98] = 9'b100010000;
assign F[127][99] = 9'b100010000;
assign F[127][100] = 9'b100010000;
assign F[127][101] = 9'b100010000;
assign F[127][102] = 9'b100010000;
assign F[127][103] = 9'b100010000;
assign F[127][104] = 9'b100010000;
assign F[127][105] = 9'b100010100;
assign F[127][106] = 9'b100010100;
assign F[127][107] = 9'b100110101;
assign F[127][108] = 9'b100110101;
assign F[127][109] = 9'b110011100;
assign F[127][110] = 9'b111111100;
assign F[127][111] = 9'b110111100;
assign F[127][112] = 9'b110011100;
assign F[127][113] = 9'b110011100;
assign F[127][114] = 9'b110011100;
assign F[127][115] = 9'b110011100;
assign F[127][116] = 9'b110111100;
assign F[127][117] = 9'b110011100;
assign F[127][118] = 9'b110011100;
assign F[127][119] = 9'b110111100;
assign F[127][120] = 9'b110111100;
assign F[127][121] = 9'b110011100;
assign F[127][122] = 9'b110011100;
assign F[127][123] = 9'b101010100;
assign F[127][124] = 9'b100110101;
assign F[127][125] = 9'b101010100;
assign F[127][126] = 9'b100010000;
assign F[127][127] = 9'b100010000;
assign F[127][128] = 9'b100010001;
assign F[127][129] = 9'b101011101;
assign F[127][130] = 9'b100110000;
assign F[127][131] = 9'b100010000;
assign F[127][132] = 9'b100010000;
assign F[127][133] = 9'b100010000;
assign F[127][134] = 9'b100010000;
assign F[127][135] = 9'b100010000;
assign F[127][136] = 9'b100010000;
assign F[127][137] = 9'b100110101;
assign F[127][138] = 9'b100110001;
assign F[127][139] = 9'b110011100;
assign F[127][140] = 9'b111111100;
assign F[127][141] = 9'b110111100;
assign F[127][142] = 9'b110011100;
assign F[127][143] = 9'b110111100;
assign F[127][144] = 9'b110111100;
assign F[127][145] = 9'b110111100;
assign F[127][146] = 9'b110111100;
assign F[127][147] = 9'b110111100;
assign F[127][148] = 9'b110011100;
assign F[127][149] = 9'b110011100;
assign F[127][150] = 9'b110011100;
assign F[127][151] = 9'b110011100;
assign F[127][152] = 9'b110011100;
assign F[127][153] = 9'b110111100;
assign F[127][154] = 9'b110111101;
assign F[128][37] = 9'b110011100;
assign F[128][38] = 9'b110011100;
assign F[128][39] = 9'b110011100;
assign F[128][40] = 9'b110111100;
assign F[128][41] = 9'b110111100;
assign F[128][42] = 9'b110111100;
assign F[128][43] = 9'b110111100;
assign F[128][44] = 9'b110011100;
assign F[128][45] = 9'b110011100;
assign F[128][46] = 9'b110011100;
assign F[128][47] = 9'b110011100;
assign F[128][48] = 9'b110111100;
assign F[128][49] = 9'b110111100;
assign F[128][50] = 9'b110011100;
assign F[128][51] = 9'b110111100;
assign F[128][52] = 9'b101111100;
assign F[128][53] = 9'b101010001;
assign F[128][54] = 9'b100110000;
assign F[128][55] = 9'b100110000;
assign F[128][56] = 9'b100010000;
assign F[128][57] = 9'b100010000;
assign F[128][58] = 9'b100010000;
assign F[128][59] = 9'b100010000;
assign F[128][60] = 9'b100110101;
assign F[128][61] = 9'b100110101;
assign F[128][62] = 9'b100110000;
assign F[128][63] = 9'b100010100;
assign F[128][64] = 9'b100010100;
assign F[128][65] = 9'b100110000;
assign F[128][66] = 9'b100010000;
assign F[128][67] = 9'b100010000;
assign F[128][68] = 9'b100010000;
assign F[128][69] = 9'b100010000;
assign F[128][70] = 9'b100010001;
assign F[128][71] = 9'b100110101;
assign F[128][72] = 9'b101110101;
assign F[128][73] = 9'b110111100;
assign F[128][74] = 9'b110111100;
assign F[128][75] = 9'b110011100;
assign F[128][76] = 9'b110011100;
assign F[128][77] = 9'b110011100;
assign F[128][78] = 9'b110011100;
assign F[128][79] = 9'b110111100;
assign F[128][80] = 9'b110011100;
assign F[128][81] = 9'b110111101;
assign F[128][82] = 9'b111111101;
assign F[128][83] = 9'b111111101;
assign F[128][84] = 9'b111111101;
assign F[128][85] = 9'b110111101;
assign F[128][86] = 9'b111111101;
assign F[128][87] = 9'b111111101;
assign F[128][88] = 9'b110111101;
assign F[128][89] = 9'b110111101;
assign F[128][90] = 9'b110111101;
assign F[128][91] = 9'b111111101;
assign F[128][92] = 9'b101110101;
assign F[128][93] = 9'b100110001;
assign F[128][94] = 9'b100010000;
assign F[128][95] = 9'b100110000;
assign F[128][96] = 9'b100010000;
assign F[128][97] = 9'b100010000;
assign F[128][98] = 9'b100010000;
assign F[128][99] = 9'b100010000;
assign F[128][100] = 9'b100110100;
assign F[128][101] = 9'b100010100;
assign F[128][102] = 9'b100110101;
assign F[128][103] = 9'b100110101;
assign F[128][104] = 9'b100110001;
assign F[128][105] = 9'b101010101;
assign F[128][106] = 9'b101010101;
assign F[128][107] = 9'b101010101;
assign F[128][108] = 9'b101010101;
assign F[128][109] = 9'b110011101;
assign F[128][110] = 9'b111111100;
assign F[128][111] = 9'b110111100;
assign F[128][112] = 9'b110011100;
assign F[128][113] = 9'b110111100;
assign F[128][114] = 9'b110011100;
assign F[128][115] = 9'b110011100;
assign F[128][116] = 9'b110011100;
assign F[128][117] = 9'b110111100;
assign F[128][118] = 9'b111111101;
assign F[128][119] = 9'b111111101;
assign F[128][120] = 9'b111111101;
assign F[128][121] = 9'b111111101;
assign F[128][122] = 9'b111111101;
assign F[128][123] = 9'b110111101;
assign F[128][124] = 9'b101010101;
assign F[128][125] = 9'b100010000;
assign F[128][126] = 9'b100010000;
assign F[128][127] = 9'b100010001;
assign F[128][128] = 9'b101010101;
assign F[128][129] = 9'b101111101;
assign F[128][130] = 9'b110011101;
assign F[128][131] = 9'b101010101;
assign F[128][132] = 9'b100010000;
assign F[128][133] = 9'b100010000;
assign F[128][134] = 9'b100110000;
assign F[128][135] = 9'b100110000;
assign F[128][136] = 9'b100010000;
assign F[128][137] = 9'b100010101;
assign F[128][138] = 9'b101010101;
assign F[128][139] = 9'b110011101;
assign F[128][140] = 9'b111111100;
assign F[128][141] = 9'b110011100;
assign F[128][142] = 9'b110011100;
assign F[128][143] = 9'b110111100;
assign F[128][144] = 9'b110011100;
assign F[128][145] = 9'b110111100;
assign F[128][146] = 9'b110111100;
assign F[128][147] = 9'b111111100;
assign F[128][148] = 9'b110111100;
assign F[128][149] = 9'b110111100;
assign F[128][150] = 9'b110011100;
assign F[128][151] = 9'b110011100;
assign F[128][152] = 9'b110011100;
assign F[128][153] = 9'b110011100;
assign F[128][154] = 9'b110011100;
assign F[129][41] = 9'b111111100;
assign F[129][42] = 9'b110111100;
assign F[129][43] = 9'b110011100;
assign F[129][44] = 9'b110011100;
assign F[129][45] = 9'b110111100;
assign F[129][46] = 9'b110111100;
assign F[129][47] = 9'b110011101;
assign F[129][54] = 9'b100110000;
assign F[129][55] = 9'b100010100;
assign F[129][56] = 9'b100010000;
assign F[129][57] = 9'b100010000;
assign F[129][58] = 9'b100010000;
assign F[129][59] = 9'b100010000;
assign F[129][60] = 9'b100110101;
assign F[129][61] = 9'b101111111;
assign F[129][62] = 9'b101110101;
assign F[129][63] = 9'b100110101;
assign F[129][64] = 9'b101010101;
assign F[129][65] = 9'b100110000;
assign F[129][66] = 9'b100010000;
assign F[129][67] = 9'b100010000;
assign F[129][68] = 9'b100010000;
assign F[129][69] = 9'b100010000;
assign F[129][70] = 9'b100010101;
assign F[129][71] = 9'b101011110;
assign F[129][74] = 9'b110111100;
assign F[129][75] = 9'b110111100;
assign F[129][76] = 9'b110011100;
assign F[129][77] = 9'b110011100;
assign F[129][78] = 9'b110011100;
assign F[129][79] = 9'b110111100;
assign F[129][80] = 9'b110011100;
assign F[129][93] = 9'b101110101;
assign F[129][94] = 9'b100110101;
assign F[129][95] = 9'b100010000;
assign F[129][96] = 9'b100010000;
assign F[129][97] = 9'b100010000;
assign F[129][98] = 9'b100010000;
assign F[129][99] = 9'b100010000;
assign F[129][100] = 9'b100110001;
assign F[129][101] = 9'b100110001;
assign F[129][102] = 9'b101011101;
assign F[129][103] = 9'b101111110;
assign F[129][111] = 9'b110111100;
assign F[129][112] = 9'b110111100;
assign F[129][113] = 9'b110111100;
assign F[129][114] = 9'b110011100;
assign F[129][115] = 9'b110011100;
assign F[129][116] = 9'b110011100;
assign F[129][117] = 9'b110111100;
assign F[129][118] = 9'b111111111;
assign F[129][119] = 9'b111111111;
assign F[129][120] = 9'b111111111;
assign F[129][121] = 9'b111111111;
assign F[129][122] = 9'b111111110;
assign F[129][123] = 9'b111111111;
assign F[129][124] = 9'b101110101;
assign F[129][125] = 9'b100010000;
assign F[129][126] = 9'b100010000;
assign F[129][127] = 9'b100110101;
assign F[129][128] = 9'b110011111;
assign F[129][129] = 9'b111111111;
assign F[129][130] = 9'b111111110;
assign F[129][131] = 9'b101111101;
assign F[129][132] = 9'b100010000;
assign F[129][133] = 9'b100010000;
assign F[129][134] = 9'b100010000;
assign F[129][135] = 9'b100010000;
assign F[129][136] = 9'b100010000;
assign F[129][137] = 9'b100010101;
assign F[129][138] = 9'b101111111;
assign F[129][141] = 9'b110111100;
assign F[129][142] = 9'b110011100;
assign F[129][143] = 9'b110111100;
assign F[129][144] = 9'b110011100;
assign F[129][148] = 9'b111111101;
assign F[129][149] = 9'b111111100;
assign F[129][150] = 9'b110111100;
assign F[129][151] = 9'b110111100;
assign F[129][152] = 9'b110111100;
assign F[129][153] = 9'b110011100;
assign F[130][41] = 9'b111111100;
assign F[130][42] = 9'b110111100;
assign F[130][43] = 9'b110011100;
assign F[130][44] = 9'b110011100;
assign F[130][45] = 9'b110111100;
assign F[130][46] = 9'b110111100;
assign F[130][47] = 9'b110011101;
assign F[130][54] = 9'b100110000;
assign F[130][55] = 9'b100010100;
assign F[130][56] = 9'b100010000;
assign F[130][57] = 9'b100010000;
assign F[130][58] = 9'b100010000;
assign F[130][59] = 9'b100010000;
assign F[130][60] = 9'b100111101;
assign F[130][61] = 9'b101111111;
assign F[130][65] = 9'b100110000;
assign F[130][66] = 9'b100010000;
assign F[130][67] = 9'b100010000;
assign F[130][68] = 9'b100010000;
assign F[130][69] = 9'b100010000;
assign F[130][70] = 9'b100110101;
assign F[130][71] = 9'b101011110;
assign F[130][74] = 9'b111111100;
assign F[130][75] = 9'b110111100;
assign F[130][76] = 9'b110011100;
assign F[130][77] = 9'b110011100;
assign F[130][78] = 9'b110011100;
assign F[130][79] = 9'b110011100;
assign F[130][80] = 9'b110011100;
assign F[130][81] = 9'b110111100;
assign F[130][82] = 9'b110111100;
assign F[130][83] = 9'b110111100;
assign F[130][84] = 9'b110111100;
assign F[130][85] = 9'b110011100;
assign F[130][93] = 9'b101110101;
assign F[130][94] = 9'b100110101;
assign F[130][95] = 9'b100010000;
assign F[130][96] = 9'b100010000;
assign F[130][97] = 9'b100010000;
assign F[130][98] = 9'b100010000;
assign F[130][99] = 9'b100110101;
assign F[130][111] = 9'b110111100;
assign F[130][112] = 9'b110111100;
assign F[130][113] = 9'b110111100;
assign F[130][114] = 9'b110011100;
assign F[130][115] = 9'b110111100;
assign F[130][116] = 9'b110011100;
assign F[130][117] = 9'b110011100;
assign F[130][118] = 9'b110111100;
assign F[130][119] = 9'b110111100;
assign F[130][120] = 9'b110111100;
assign F[130][121] = 9'b110111100;
assign F[130][122] = 9'b110111100;
assign F[130][123] = 9'b111111101;
assign F[130][124] = 9'b101010100;
assign F[130][125] = 9'b100010000;
assign F[130][126] = 9'b100010000;
assign F[130][127] = 9'b100110101;
assign F[130][128] = 9'b100110101;
assign F[130][129] = 9'b100110101;
assign F[130][130] = 9'b100110100;
assign F[130][131] = 9'b100010100;
assign F[130][132] = 9'b100010000;
assign F[130][133] = 9'b100010000;
assign F[130][134] = 9'b100010000;
assign F[130][135] = 9'b100010000;
assign F[130][136] = 9'b100110000;
assign F[130][137] = 9'b100010101;
assign F[130][138] = 9'b100110001;
assign F[130][141] = 9'b110111100;
assign F[130][142] = 9'b110011100;
assign F[130][143] = 9'b110111100;
assign F[130][144] = 9'b110011100;
assign F[130][150] = 9'b111111101;
assign F[130][151] = 9'b110111100;
assign F[130][152] = 9'b111111100;
assign F[130][153] = 9'b110011100;
assign F[131][41] = 9'b111111100;
assign F[131][42] = 9'b111111100;
assign F[131][43] = 9'b110111100;
assign F[131][44] = 9'b110111100;
assign F[131][45] = 9'b110111100;
assign F[131][46] = 9'b110111100;
assign F[131][47] = 9'b110011101;
assign F[131][54] = 9'b100110000;
assign F[131][55] = 9'b100110101;
assign F[131][56] = 9'b100110100;
assign F[131][57] = 9'b100110100;
assign F[131][58] = 9'b100110100;
assign F[131][59] = 9'b100010100;
assign F[131][60] = 9'b100111101;
assign F[131][61] = 9'b101111111;
assign F[131][65] = 9'b101010101;
assign F[131][66] = 9'b100010100;
assign F[131][67] = 9'b100110100;
assign F[131][68] = 9'b100110100;
assign F[131][69] = 9'b100010100;
assign F[131][70] = 9'b100110101;
assign F[131][71] = 9'b101011110;
assign F[131][74] = 9'b111111100;
assign F[131][75] = 9'b111111100;
assign F[131][76] = 9'b110111100;
assign F[131][77] = 9'b110111100;
assign F[131][78] = 9'b110111100;
assign F[131][79] = 9'b110111100;
assign F[131][80] = 9'b110111100;
assign F[131][81] = 9'b110111100;
assign F[131][82] = 9'b110111100;
assign F[131][83] = 9'b110111100;
assign F[131][84] = 9'b110111100;
assign F[131][85] = 9'b110011100;
assign F[131][93] = 9'b101110101;
assign F[131][94] = 9'b100111101;
assign F[131][95] = 9'b100010100;
assign F[131][96] = 9'b100110101;
assign F[131][97] = 9'b100110100;
assign F[131][98] = 9'b100110100;
assign F[131][99] = 9'b100110101;
assign F[131][100] = 9'b100110101;
assign F[131][111] = 9'b111111100;
assign F[131][112] = 9'b110111100;
assign F[131][113] = 9'b110111100;
assign F[131][114] = 9'b110111100;
assign F[131][115] = 9'b110111100;
assign F[131][116] = 9'b110111100;
assign F[131][117] = 9'b110111100;
assign F[131][118] = 9'b110111100;
assign F[131][119] = 9'b110111100;
assign F[131][120] = 9'b110111100;
assign F[131][121] = 9'b110111100;
assign F[131][122] = 9'b110111101;
assign F[131][123] = 9'b110010101;
assign F[131][124] = 9'b100111100;
assign F[131][125] = 9'b100010100;
assign F[131][126] = 9'b100110101;
assign F[131][127] = 9'b101111101;
assign F[131][128] = 9'b101010000;
assign F[131][129] = 9'b100010000;
assign F[131][130] = 9'b100110101;
assign F[131][131] = 9'b101111101;
assign F[131][132] = 9'b101010101;
assign F[131][133] = 9'b100010100;
assign F[131][134] = 9'b100010100;
assign F[131][135] = 9'b100010100;
assign F[131][136] = 9'b100110100;
assign F[131][137] = 9'b100110100;
assign F[131][138] = 9'b100110101;
assign F[131][141] = 9'b111111100;
assign F[131][142] = 9'b110111100;
assign F[131][143] = 9'b111111100;
assign F[131][144] = 9'b110011100;
assign F[131][152] = 9'b111111100;
assign F[131][153] = 9'b110111100;
assign F[132][41] = 9'b111111101;
assign F[132][42] = 9'b110111100;
assign F[132][43] = 9'b110011100;
assign F[132][44] = 9'b110011100;
assign F[132][45] = 9'b110111100;
assign F[132][46] = 9'b110111100;
assign F[132][54] = 9'b101010000;
assign F[132][55] = 9'b100110000;
assign F[132][56] = 9'b100110000;
assign F[132][57] = 9'b100110000;
assign F[132][58] = 9'b100110000;
assign F[132][59] = 9'b100010000;
assign F[132][60] = 9'b100110101;
assign F[132][61] = 9'b101111111;
assign F[132][65] = 9'b101010001;
assign F[132][66] = 9'b100010000;
assign F[132][67] = 9'b100110000;
assign F[132][68] = 9'b100110000;
assign F[132][69] = 9'b100110000;
assign F[132][70] = 9'b100110001;
assign F[132][74] = 9'b111111100;
assign F[132][75] = 9'b110111100;
assign F[132][76] = 9'b110011100;
assign F[132][77] = 9'b110011100;
assign F[132][78] = 9'b110011100;
assign F[132][79] = 9'b110011100;
assign F[132][80] = 9'b110111100;
assign F[132][81] = 9'b110111100;
assign F[132][82] = 9'b110011100;
assign F[132][83] = 9'b110111100;
assign F[132][84] = 9'b110011100;
assign F[132][94] = 9'b100110001;
assign F[132][95] = 9'b100110000;
assign F[132][96] = 9'b100110000;
assign F[132][97] = 9'b100110000;
assign F[132][98] = 9'b100110000;
assign F[132][99] = 9'b100110001;
assign F[132][111] = 9'b110111100;
assign F[132][112] = 9'b110111100;
assign F[132][113] = 9'b110111100;
assign F[132][114] = 9'b110011100;
assign F[132][115] = 9'b110011100;
assign F[132][116] = 9'b110011100;
assign F[132][117] = 9'b110011100;
assign F[132][118] = 9'b110011100;
assign F[132][119] = 9'b110011100;
assign F[132][120] = 9'b110011100;
assign F[132][121] = 9'b110111100;
assign F[132][122] = 9'b110111101;
assign F[132][124] = 9'b100110000;
assign F[132][125] = 9'b100010000;
assign F[132][126] = 9'b100110001;
assign F[132][129] = 9'b101010001;
assign F[132][133] = 9'b100110000;
assign F[132][134] = 9'b100110001;
assign F[132][135] = 9'b100110000;
assign F[132][136] = 9'b100110000;
assign F[132][137] = 9'b100110000;
assign F[132][138] = 9'b100110001;
assign F[132][141] = 9'b110111100;
assign F[132][142] = 9'b110011100;
assign F[132][143] = 9'b110111100;
assign F[141][69] = 9'b100110000;
assign F[141][70] = 9'b100110000;
assign F[141][71] = 9'b100110000;
assign F[141][72] = 9'b100110000;
assign F[141][73] = 9'b100110000;
assign F[141][74] = 9'b100110000;
assign F[141][75] = 9'b100010001;
assign F[141][84] = 9'b110111100;
assign F[141][85] = 9'b110011100;
assign F[141][86] = 9'b110011100;
assign F[141][87] = 9'b110011100;
assign F[141][88] = 9'b110111100;
assign F[141][89] = 9'b110011100;
assign F[141][96] = 9'b100110000;
assign F[141][97] = 9'b100010001;
assign F[141][98] = 9'b100110001;
assign F[141][99] = 9'b100110000;
assign F[141][100] = 9'b100110000;
assign F[141][101] = 9'b100110001;
assign F[141][110] = 9'b100110000;
assign F[141][111] = 9'b100010000;
assign F[141][112] = 9'b100010000;
assign F[141][113] = 9'b100110001;
assign F[141][114] = 9'b100110001;
assign F[141][118] = 9'b110111100;
assign F[141][119] = 9'b110011100;
assign F[141][120] = 9'b110111100;
assign F[141][121] = 9'b110111100;
assign F[141][122] = 9'b110111100;
assign F[141][123] = 9'b110111100;
assign F[141][124] = 9'b110111100;
assign F[141][125] = 9'b110011100;
assign F[141][126] = 9'b110011100;
assign F[141][127] = 9'b110011100;
assign F[141][128] = 9'b110011100;
assign F[141][129] = 9'b110111100;
assign F[142][65] = 9'b101110101;
assign F[142][66] = 9'b100110001;
assign F[142][67] = 9'b100110000;
assign F[142][68] = 9'b100010100;
assign F[142][69] = 9'b100110100;
assign F[142][70] = 9'b100110100;
assign F[142][71] = 9'b100110100;
assign F[142][72] = 9'b100110100;
assign F[142][73] = 9'b100110100;
assign F[142][74] = 9'b100110100;
assign F[142][75] = 9'b100010101;
assign F[142][76] = 9'b100110101;
assign F[142][82] = 9'b111111100;
assign F[142][83] = 9'b110111100;
assign F[142][84] = 9'b110111100;
assign F[142][85] = 9'b110111100;
assign F[142][86] = 9'b110111100;
assign F[142][87] = 9'b110111100;
assign F[142][88] = 9'b110111100;
assign F[142][89] = 9'b110111100;
assign F[142][90] = 9'b110111101;
assign F[142][96] = 9'b100110000;
assign F[142][97] = 9'b100010100;
assign F[142][98] = 9'b100110101;
assign F[142][99] = 9'b100010100;
assign F[142][100] = 9'b100110100;
assign F[142][101] = 9'b100010101;
assign F[142][102] = 9'b100110001;
assign F[142][103] = 9'b101111111;
assign F[142][108] = 9'b110011101;
assign F[142][109] = 9'b100110000;
assign F[142][110] = 9'b100010100;
assign F[142][111] = 9'b100010100;
assign F[142][112] = 9'b100110100;
assign F[142][113] = 9'b100010100;
assign F[142][114] = 9'b100010101;
assign F[142][117] = 9'b111111100;
assign F[142][118] = 9'b111111100;
assign F[142][119] = 9'b110111100;
assign F[142][120] = 9'b110111100;
assign F[142][121] = 9'b110111100;
assign F[142][122] = 9'b110111100;
assign F[142][123] = 9'b110111100;
assign F[142][124] = 9'b110111100;
assign F[142][125] = 9'b110111100;
assign F[142][126] = 9'b110111100;
assign F[142][127] = 9'b110111100;
assign F[142][128] = 9'b110111100;
assign F[142][129] = 9'b110011100;
assign F[143][64] = 9'b110010101;
assign F[143][65] = 9'b100110001;
assign F[143][66] = 9'b100110100;
assign F[143][67] = 9'b100010100;
assign F[143][68] = 9'b100010000;
assign F[143][69] = 9'b100010000;
assign F[143][70] = 9'b100010000;
assign F[143][71] = 9'b100010000;
assign F[143][72] = 9'b100010000;
assign F[143][73] = 9'b100010000;
assign F[143][74] = 9'b100010000;
assign F[143][75] = 9'b100010000;
assign F[143][76] = 9'b100110101;
assign F[143][77] = 9'b110011111;
assign F[143][82] = 9'b111111100;
assign F[143][83] = 9'b110111100;
assign F[143][84] = 9'b110011100;
assign F[143][85] = 9'b110011100;
assign F[143][86] = 9'b110011100;
assign F[143][87] = 9'b110011100;
assign F[143][88] = 9'b110011100;
assign F[143][89] = 9'b110111100;
assign F[143][90] = 9'b110011101;
assign F[143][96] = 9'b100110000;
assign F[143][97] = 9'b100010000;
assign F[143][98] = 9'b100010000;
assign F[143][99] = 9'b100010000;
assign F[143][100] = 9'b100110000;
assign F[143][101] = 9'b100010000;
assign F[143][102] = 9'b100010101;
assign F[143][103] = 9'b100110101;
assign F[143][108] = 9'b101010000;
assign F[143][109] = 9'b100010100;
assign F[143][110] = 9'b100010000;
assign F[143][111] = 9'b100010000;
assign F[143][112] = 9'b100010000;
assign F[143][113] = 9'b100010000;
assign F[143][114] = 9'b100010001;
assign F[143][117] = 9'b111111100;
assign F[143][118] = 9'b110111100;
assign F[143][119] = 9'b110011100;
assign F[143][120] = 9'b110111100;
assign F[143][121] = 9'b110011100;
assign F[143][122] = 9'b110011100;
assign F[143][123] = 9'b110011100;
assign F[143][124] = 9'b110011100;
assign F[143][125] = 9'b110011100;
assign F[143][126] = 9'b110011100;
assign F[143][127] = 9'b110011100;
assign F[143][128] = 9'b110111100;
assign F[143][129] = 9'b110011100;
assign F[144][63] = 9'b101110101;
assign F[144][64] = 9'b100110100;
assign F[144][65] = 9'b100010001;
assign F[144][66] = 9'b100010000;
assign F[144][67] = 9'b100010000;
assign F[144][68] = 9'b100010000;
assign F[144][69] = 9'b100010000;
assign F[144][70] = 9'b100010000;
assign F[144][71] = 9'b100010000;
assign F[144][72] = 9'b100010000;
assign F[144][73] = 9'b100010000;
assign F[144][74] = 9'b100010000;
assign F[144][75] = 9'b100010000;
assign F[144][76] = 9'b100110101;
assign F[144][82] = 9'b111111100;
assign F[144][83] = 9'b110111100;
assign F[144][84] = 9'b110011100;
assign F[144][85] = 9'b110011100;
assign F[144][86] = 9'b110011100;
assign F[144][87] = 9'b110011100;
assign F[144][88] = 9'b110011100;
assign F[144][89] = 9'b110111100;
assign F[144][90] = 9'b110011100;
assign F[144][96] = 9'b100110000;
assign F[144][97] = 9'b100010000;
assign F[144][98] = 9'b100010000;
assign F[144][99] = 9'b100010000;
assign F[144][100] = 9'b100010000;
assign F[144][101] = 9'b100010000;
assign F[144][102] = 9'b100110000;
assign F[144][103] = 9'b100010101;
assign F[144][104] = 9'b100110101;
assign F[144][107] = 9'b101110101;
assign F[144][108] = 9'b100010000;
assign F[144][109] = 9'b100110000;
assign F[144][110] = 9'b100010000;
assign F[144][111] = 9'b100010000;
assign F[144][112] = 9'b100010000;
assign F[144][113] = 9'b100010000;
assign F[144][114] = 9'b100010001;
assign F[144][117] = 9'b111111100;
assign F[144][118] = 9'b110111100;
assign F[144][119] = 9'b110011100;
assign F[144][120] = 9'b110111100;
assign F[144][121] = 9'b110011100;
assign F[144][122] = 9'b110011100;
assign F[144][123] = 9'b110011100;
assign F[144][124] = 9'b110011100;
assign F[144][125] = 9'b110011100;
assign F[144][126] = 9'b110011100;
assign F[144][127] = 9'b110011100;
assign F[144][128] = 9'b110111100;
assign F[144][129] = 9'b110011100;
assign F[145][62] = 9'b111111101;
assign F[145][63] = 9'b100110100;
assign F[145][64] = 9'b100010000;
assign F[145][65] = 9'b100110000;
assign F[145][66] = 9'b100010000;
assign F[145][67] = 9'b100010000;
assign F[145][68] = 9'b100010000;
assign F[145][69] = 9'b100010000;
assign F[145][70] = 9'b100110000;
assign F[145][71] = 9'b100010000;
assign F[145][72] = 9'b100010000;
assign F[145][73] = 9'b100010000;
assign F[145][74] = 9'b100010000;
assign F[145][75] = 9'b100010000;
assign F[145][76] = 9'b100110101;
assign F[145][77] = 9'b101111111;
assign F[145][81] = 9'b111111101;
assign F[145][82] = 9'b111111100;
assign F[145][83] = 9'b110011100;
assign F[145][84] = 9'b110011100;
assign F[145][85] = 9'b110011100;
assign F[145][86] = 9'b110011100;
assign F[145][87] = 9'b110011100;
assign F[145][88] = 9'b110011100;
assign F[145][89] = 9'b110111100;
assign F[145][90] = 9'b110011100;
assign F[145][96] = 9'b100110000;
assign F[145][97] = 9'b100010000;
assign F[145][98] = 9'b100010000;
assign F[145][99] = 9'b100010000;
assign F[145][100] = 9'b100110000;
assign F[145][101] = 9'b100010000;
assign F[145][102] = 9'b100010000;
assign F[145][103] = 9'b100010000;
assign F[145][104] = 9'b100110001;
assign F[145][106] = 9'b101110101;
assign F[145][107] = 9'b100110100;
assign F[145][108] = 9'b100010000;
assign F[145][109] = 9'b100010000;
assign F[145][110] = 9'b100010000;
assign F[145][111] = 9'b100010000;
assign F[145][112] = 9'b100010000;
assign F[145][113] = 9'b100010000;
assign F[145][114] = 9'b100010001;
assign F[145][117] = 9'b111111100;
assign F[145][118] = 9'b110111100;
assign F[145][119] = 9'b110011100;
assign F[145][120] = 9'b110011100;
assign F[145][121] = 9'b110011100;
assign F[145][122] = 9'b110011100;
assign F[145][123] = 9'b110011100;
assign F[145][124] = 9'b110011100;
assign F[145][125] = 9'b110011100;
assign F[145][126] = 9'b110011100;
assign F[145][127] = 9'b110111100;
assign F[145][128] = 9'b110111100;
assign F[145][129] = 9'b110011100;
assign F[146][62] = 9'b110010101;
assign F[146][63] = 9'b100110100;
assign F[146][64] = 9'b100010000;
assign F[146][65] = 9'b100010000;
assign F[146][66] = 9'b100010000;
assign F[146][67] = 9'b100010000;
assign F[146][68] = 9'b100010000;
assign F[146][69] = 9'b100010000;
assign F[146][70] = 9'b100110000;
assign F[146][71] = 9'b100010000;
assign F[146][72] = 9'b100010100;
assign F[146][73] = 9'b100110101;
assign F[146][74] = 9'b100110101;
assign F[146][75] = 9'b100110100;
assign F[146][76] = 9'b100110001;
assign F[146][81] = 9'b111111100;
assign F[146][82] = 9'b110111100;
assign F[146][83] = 9'b110011100;
assign F[146][84] = 9'b110011100;
assign F[146][85] = 9'b110011100;
assign F[146][86] = 9'b110011100;
assign F[146][87] = 9'b110011100;
assign F[146][88] = 9'b110011100;
assign F[146][89] = 9'b110111100;
assign F[146][90] = 9'b110011100;
assign F[146][91] = 9'b110011101;
assign F[146][96] = 9'b101010101;
assign F[146][97] = 9'b100010000;
assign F[146][98] = 9'b100110000;
assign F[146][99] = 9'b100010000;
assign F[146][100] = 9'b100010000;
assign F[146][101] = 9'b100010000;
assign F[146][102] = 9'b100010000;
assign F[146][103] = 9'b100010000;
assign F[146][104] = 9'b100010000;
assign F[146][105] = 9'b100110001;
assign F[146][106] = 9'b100110000;
assign F[146][107] = 9'b100010000;
assign F[146][108] = 9'b100010000;
assign F[146][109] = 9'b100010000;
assign F[146][110] = 9'b100110000;
assign F[146][111] = 9'b100010000;
assign F[146][112] = 9'b100010000;
assign F[146][113] = 9'b100110000;
assign F[146][114] = 9'b100010101;
assign F[146][117] = 9'b111111100;
assign F[146][118] = 9'b110111100;
assign F[146][119] = 9'b110011100;
assign F[146][120] = 9'b110011100;
assign F[146][121] = 9'b110011100;
assign F[146][122] = 9'b110011100;
assign F[146][123] = 9'b110011100;
assign F[146][124] = 9'b110011100;
assign F[146][125] = 9'b110011100;
assign F[146][126] = 9'b110111100;
assign F[146][127] = 9'b110111100;
assign F[146][128] = 9'b111111100;
assign F[146][129] = 9'b110011100;
assign F[147][62] = 9'b101010000;
assign F[147][63] = 9'b100010100;
assign F[147][64] = 9'b100010000;
assign F[147][65] = 9'b100010000;
assign F[147][66] = 9'b100010000;
assign F[147][67] = 9'b100010000;
assign F[147][68] = 9'b100010000;
assign F[147][69] = 9'b100010000;
assign F[147][70] = 9'b100010100;
assign F[147][71] = 9'b100110101;
assign F[147][72] = 9'b101010101;
assign F[147][73] = 9'b101010101;
assign F[147][74] = 9'b101110101;
assign F[147][75] = 9'b101110101;
assign F[147][81] = 9'b111111100;
assign F[147][82] = 9'b110111100;
assign F[147][83] = 9'b110011100;
assign F[147][84] = 9'b110011100;
assign F[147][85] = 9'b110011100;
assign F[147][86] = 9'b110011100;
assign F[147][87] = 9'b110011100;
assign F[147][88] = 9'b110011100;
assign F[147][89] = 9'b110011100;
assign F[147][90] = 9'b110111100;
assign F[147][91] = 9'b110011100;
assign F[147][96] = 9'b101010101;
assign F[147][97] = 9'b100010000;
assign F[147][98] = 9'b100010000;
assign F[147][99] = 9'b100010000;
assign F[147][100] = 9'b100010000;
assign F[147][101] = 9'b100010000;
assign F[147][102] = 9'b100010000;
assign F[147][103] = 9'b100010000;
assign F[147][104] = 9'b100010000;
assign F[147][105] = 9'b100010000;
assign F[147][106] = 9'b100010000;
assign F[147][107] = 9'b100010000;
assign F[147][108] = 9'b100010000;
assign F[147][109] = 9'b100010000;
assign F[147][110] = 9'b100110000;
assign F[147][111] = 9'b100010000;
assign F[147][112] = 9'b100010000;
assign F[147][113] = 9'b100110000;
assign F[147][114] = 9'b100010101;
assign F[147][117] = 9'b111111100;
assign F[147][118] = 9'b110111100;
assign F[147][119] = 9'b110111100;
assign F[147][120] = 9'b110011100;
assign F[147][121] = 9'b110011100;
assign F[147][122] = 9'b110011100;
assign F[147][123] = 9'b110011100;
assign F[147][124] = 9'b110111100;
assign F[147][125] = 9'b111111101;
assign F[147][126] = 9'b111111101;
assign F[147][127] = 9'b111111101;
assign F[147][128] = 9'b110111100;
assign F[148][62] = 9'b100110001;
assign F[148][63] = 9'b100010101;
assign F[148][64] = 9'b100010000;
assign F[148][65] = 9'b100110000;
assign F[148][66] = 9'b100010000;
assign F[148][67] = 9'b100010000;
assign F[148][68] = 9'b100010000;
assign F[148][69] = 9'b100010001;
assign F[148][70] = 9'b100110001;
assign F[148][71] = 9'b110011111;
assign F[148][81] = 9'b111111100;
assign F[148][82] = 9'b110111100;
assign F[148][83] = 9'b110011100;
assign F[148][84] = 9'b110011100;
assign F[148][85] = 9'b110011100;
assign F[148][86] = 9'b110011100;
assign F[148][87] = 9'b110011100;
assign F[148][88] = 9'b110011100;
assign F[148][89] = 9'b110011100;
assign F[148][90] = 9'b110111100;
assign F[148][91] = 9'b110111100;
assign F[148][92] = 9'b110111101;
assign F[148][96] = 9'b101010101;
assign F[148][97] = 9'b100010000;
assign F[148][98] = 9'b100010000;
assign F[148][99] = 9'b100010000;
assign F[148][100] = 9'b100010000;
assign F[148][101] = 9'b100010000;
assign F[148][102] = 9'b100010000;
assign F[148][103] = 9'b100010000;
assign F[148][104] = 9'b100010000;
assign F[148][105] = 9'b100010000;
assign F[148][106] = 9'b100010000;
assign F[148][107] = 9'b100010000;
assign F[148][108] = 9'b100010000;
assign F[148][109] = 9'b100010000;
assign F[148][110] = 9'b100110000;
assign F[148][111] = 9'b100010000;
assign F[148][112] = 9'b100010000;
assign F[148][113] = 9'b100110000;
assign F[148][114] = 9'b100010101;
assign F[148][117] = 9'b111111100;
assign F[148][118] = 9'b110111100;
assign F[148][119] = 9'b110111100;
assign F[148][120] = 9'b110011100;
assign F[148][121] = 9'b110011100;
assign F[148][122] = 9'b110111100;
assign F[148][123] = 9'b110011100;
assign F[148][124] = 9'b110111101;
assign F[148][125] = 9'b111111111;
assign F[149][62] = 9'b100110101;
assign F[149][63] = 9'b100010100;
assign F[149][64] = 9'b100010000;
assign F[149][65] = 9'b100110000;
assign F[149][66] = 9'b100010000;
assign F[149][67] = 9'b100110000;
assign F[149][68] = 9'b100010101;
assign F[149][69] = 9'b100110101;
assign F[149][75] = 9'b100110000;
assign F[149][76] = 9'b100010000;
assign F[149][77] = 9'b100010001;
assign F[149][80] = 9'b111111101;
assign F[149][81] = 9'b111111100;
assign F[149][82] = 9'b110011100;
assign F[149][83] = 9'b110011100;
assign F[149][84] = 9'b110111101;
assign F[149][85] = 9'b111111100;
assign F[149][86] = 9'b110111100;
assign F[149][87] = 9'b110011100;
assign F[149][88] = 9'b110111100;
assign F[149][89] = 9'b110011100;
assign F[149][90] = 9'b110011100;
assign F[149][91] = 9'b110111100;
assign F[149][92] = 9'b110011100;
assign F[149][96] = 9'b101010001;
assign F[149][97] = 9'b100010000;
assign F[149][98] = 9'b100010000;
assign F[149][99] = 9'b100010000;
assign F[149][100] = 9'b100010000;
assign F[149][101] = 9'b100010000;
assign F[149][102] = 9'b100110000;
assign F[149][103] = 9'b100010000;
assign F[149][104] = 9'b100010000;
assign F[149][105] = 9'b100010000;
assign F[149][106] = 9'b100010000;
assign F[149][107] = 9'b100010000;
assign F[149][108] = 9'b100010000;
assign F[149][109] = 9'b100010000;
assign F[149][110] = 9'b100010000;
assign F[149][111] = 9'b100110001;
assign F[149][112] = 9'b100010000;
assign F[149][113] = 9'b100110000;
assign F[149][114] = 9'b100110101;
assign F[149][117] = 9'b111111101;
assign F[149][118] = 9'b110111100;
assign F[149][119] = 9'b110111100;
assign F[149][120] = 9'b110011100;
assign F[149][121] = 9'b110011100;
assign F[149][122] = 9'b110011100;
assign F[149][123] = 9'b110011100;
assign F[149][124] = 9'b110011100;
assign F[149][125] = 9'b110011100;
assign F[149][126] = 9'b110111100;
assign F[149][127] = 9'b110111100;
assign F[149][128] = 9'b111111100;
assign F[149][129] = 9'b111111101;
assign F[150][62] = 9'b100110000;
assign F[150][63] = 9'b100010100;
assign F[150][64] = 9'b100110000;
assign F[150][65] = 9'b100010000;
assign F[150][66] = 9'b100010000;
assign F[150][67] = 9'b100110000;
assign F[150][68] = 9'b100010100;
assign F[150][69] = 9'b100110101;
assign F[150][70] = 9'b100110000;
assign F[150][71] = 9'b100010000;
assign F[150][72] = 9'b100010000;
assign F[150][73] = 9'b100110000;
assign F[150][74] = 9'b100010000;
assign F[150][75] = 9'b100110101;
assign F[150][76] = 9'b100010100;
assign F[150][77] = 9'b100010101;
assign F[150][78] = 9'b100110101;
assign F[150][79] = 9'b110111100;
assign F[150][80] = 9'b110111100;
assign F[150][81] = 9'b110111100;
assign F[150][82] = 9'b110011100;
assign F[150][83] = 9'b110011100;
assign F[150][84] = 9'b110111100;
assign F[150][85] = 9'b111111100;
assign F[150][86] = 9'b110011100;
assign F[150][87] = 9'b110011100;
assign F[150][88] = 9'b110011100;
assign F[150][89] = 9'b110011100;
assign F[150][90] = 9'b110011100;
assign F[150][91] = 9'b110111100;
assign F[150][92] = 9'b110111100;
assign F[150][93] = 9'b110111100;
assign F[150][94] = 9'b110011100;
assign F[150][95] = 9'b101010101;
assign F[150][96] = 9'b100110001;
assign F[150][97] = 9'b100110000;
assign F[150][98] = 9'b100010000;
assign F[150][99] = 9'b100010000;
assign F[150][100] = 9'b100110000;
assign F[150][101] = 9'b100010000;
assign F[150][102] = 9'b100010000;
assign F[150][103] = 9'b100110000;
assign F[150][104] = 9'b100110000;
assign F[150][105] = 9'b100010000;
assign F[150][106] = 9'b100110000;
assign F[150][107] = 9'b100010000;
assign F[150][108] = 9'b100010000;
assign F[150][109] = 9'b100010000;
assign F[150][110] = 9'b100010000;
assign F[150][111] = 9'b100110000;
assign F[150][112] = 9'b100110000;
assign F[150][113] = 9'b100010000;
assign F[150][114] = 9'b100010001;
assign F[150][115] = 9'b100110101;
assign F[150][116] = 9'b101111100;
assign F[150][117] = 9'b111111100;
assign F[150][118] = 9'b110111100;
assign F[150][119] = 9'b110011100;
assign F[150][120] = 9'b110011100;
assign F[150][121] = 9'b110011100;
assign F[150][122] = 9'b110011100;
assign F[150][123] = 9'b110011100;
assign F[150][124] = 9'b110111100;
assign F[150][125] = 9'b110111100;
assign F[150][126] = 9'b110111100;
assign F[150][127] = 9'b110111100;
assign F[150][128] = 9'b110111100;
assign F[150][129] = 9'b110111100;
assign F[150][130] = 9'b110111100;
assign F[150][131] = 9'b111111101;
assign F[151][62] = 9'b100110001;
assign F[151][63] = 9'b100010100;
assign F[151][64] = 9'b100010000;
assign F[151][65] = 9'b100110000;
assign F[151][66] = 9'b100010000;
assign F[151][67] = 9'b100110000;
assign F[151][68] = 9'b100010000;
assign F[151][69] = 9'b100110001;
assign F[151][70] = 9'b100111101;
assign F[151][71] = 9'b101111101;
assign F[151][72] = 9'b101011101;
assign F[151][73] = 9'b101111101;
assign F[151][74] = 9'b100110100;
assign F[151][75] = 9'b100110000;
assign F[151][76] = 9'b100010000;
assign F[151][77] = 9'b100010001;
assign F[151][78] = 9'b101011101;
assign F[151][79] = 9'b111111101;
assign F[151][80] = 9'b110111100;
assign F[151][81] = 9'b110011100;
assign F[151][82] = 9'b110011100;
assign F[151][83] = 9'b110111100;
assign F[151][84] = 9'b111111101;
assign F[151][85] = 9'b111111101;
assign F[151][86] = 9'b111111100;
assign F[151][87] = 9'b110111100;
assign F[151][88] = 9'b110011100;
assign F[151][89] = 9'b110011100;
assign F[151][90] = 9'b110011100;
assign F[151][91] = 9'b110011100;
assign F[151][92] = 9'b110111100;
assign F[151][93] = 9'b110111100;
assign F[151][94] = 9'b110011100;
assign F[151][95] = 9'b100110000;
assign F[151][96] = 9'b100010000;
assign F[151][97] = 9'b100010100;
assign F[151][98] = 9'b100010000;
assign F[151][99] = 9'b100110000;
assign F[151][100] = 9'b100110001;
assign F[151][101] = 9'b100110101;
assign F[151][102] = 9'b100110000;
assign F[151][103] = 9'b100010000;
assign F[151][104] = 9'b100010000;
assign F[151][105] = 9'b100010000;
assign F[151][106] = 9'b100010000;
assign F[151][107] = 9'b100010000;
assign F[151][108] = 9'b100010000;
assign F[151][109] = 9'b100110101;
assign F[151][110] = 9'b101010101;
assign F[151][111] = 9'b100110000;
assign F[151][112] = 9'b100010000;
assign F[151][113] = 9'b100010000;
assign F[151][114] = 9'b100010001;
assign F[151][115] = 9'b100110101;
assign F[151][116] = 9'b101110100;
assign F[151][117] = 9'b110111100;
assign F[151][118] = 9'b110011100;
assign F[151][119] = 9'b110011100;
assign F[151][120] = 9'b110011100;
assign F[151][121] = 9'b110011100;
assign F[151][122] = 9'b110111100;
assign F[151][123] = 9'b110111100;
assign F[151][124] = 9'b110011100;
assign F[151][125] = 9'b110011100;
assign F[151][126] = 9'b110111100;
assign F[151][127] = 9'b110111100;
assign F[151][128] = 9'b110111100;
assign F[151][129] = 9'b110111100;
assign F[151][130] = 9'b110111100;
assign F[151][131] = 9'b111111101;
assign F[152][63] = 9'b101010001;
assign F[152][64] = 9'b100010100;
assign F[152][65] = 9'b100110000;
assign F[152][66] = 9'b100010000;
assign F[152][67] = 9'b100010000;
assign F[152][68] = 9'b100010000;
assign F[152][69] = 9'b100010000;
assign F[152][70] = 9'b100110101;
assign F[152][71] = 9'b110011111;
assign F[152][72] = 9'b111111111;
assign F[152][73] = 9'b111111111;
assign F[152][74] = 9'b101010101;
assign F[152][75] = 9'b100010000;
assign F[152][76] = 9'b100010000;
assign F[152][77] = 9'b100010000;
assign F[152][78] = 9'b101111111;
assign F[152][79] = 9'b111111111;
assign F[152][80] = 9'b110111100;
assign F[152][81] = 9'b110011100;
assign F[152][82] = 9'b110011100;
assign F[152][83] = 9'b111111101;
assign F[152][84] = 9'b111111111;
assign F[152][85] = 9'b111111111;
assign F[152][86] = 9'b111111101;
assign F[152][87] = 9'b110111100;
assign F[152][88] = 9'b110011100;
assign F[152][89] = 9'b110011100;
assign F[152][90] = 9'b110011100;
assign F[152][91] = 9'b110011100;
assign F[152][92] = 9'b110111100;
assign F[152][93] = 9'b110111100;
assign F[152][96] = 9'b101010000;
assign F[152][97] = 9'b100110100;
assign F[152][98] = 9'b100110000;
assign F[152][99] = 9'b100010000;
assign F[152][100] = 9'b100010101;
assign F[152][101] = 9'b110011111;
assign F[152][102] = 9'b101110101;
assign F[152][103] = 9'b100010000;
assign F[152][104] = 9'b100010000;
assign F[152][105] = 9'b100010000;
assign F[152][106] = 9'b100010000;
assign F[152][107] = 9'b100010000;
assign F[152][108] = 9'b100110001;
assign F[152][109] = 9'b101111111;
assign F[152][110] = 9'b110111101;
assign F[152][111] = 9'b100110000;
assign F[152][112] = 9'b100010001;
assign F[152][113] = 9'b100110000;
assign F[152][114] = 9'b100110101;
assign F[152][115] = 9'b110011111;
assign F[152][118] = 9'b110111100;
assign F[152][119] = 9'b110011100;
assign F[152][120] = 9'b110011100;
assign F[152][121] = 9'b110011100;
assign F[152][122] = 9'b110111100;
assign F[152][123] = 9'b110111100;
assign F[152][124] = 9'b110011100;
assign F[153][64] = 9'b101010100;
assign F[153][65] = 9'b100010100;
assign F[153][66] = 9'b100010100;
assign F[153][67] = 9'b100110000;
assign F[153][68] = 9'b100010000;
assign F[153][69] = 9'b100010000;
assign F[153][70] = 9'b100010000;
assign F[153][71] = 9'b100010001;
assign F[153][72] = 9'b100110101;
assign F[153][73] = 9'b101010101;
assign F[153][74] = 9'b100110000;
assign F[153][75] = 9'b100010000;
assign F[153][76] = 9'b100010000;
assign F[153][77] = 9'b100010001;
assign F[153][78] = 9'b110011111;
assign F[153][79] = 9'b111111101;
assign F[153][80] = 9'b110111100;
assign F[153][81] = 9'b110011100;
assign F[153][82] = 9'b110011100;
assign F[153][83] = 9'b110111100;
assign F[153][84] = 9'b110111100;
assign F[153][85] = 9'b110111100;
assign F[153][86] = 9'b110111100;
assign F[153][87] = 9'b110111100;
assign F[153][88] = 9'b110011100;
assign F[153][89] = 9'b110011100;
assign F[153][90] = 9'b110011100;
assign F[153][91] = 9'b110111100;
assign F[153][92] = 9'b110111100;
assign F[153][93] = 9'b110011100;
assign F[153][96] = 9'b101010000;
assign F[153][97] = 9'b100110100;
assign F[153][98] = 9'b100010000;
assign F[153][99] = 9'b100010000;
assign F[153][100] = 9'b100111110;
assign F[153][101] = 9'b110011111;
assign F[153][103] = 9'b101010100;
assign F[153][104] = 9'b100110000;
assign F[153][105] = 9'b100010000;
assign F[153][106] = 9'b100010000;
assign F[153][107] = 9'b100110001;
assign F[153][108] = 9'b101011110;
assign F[153][111] = 9'b100110000;
assign F[153][112] = 9'b100010000;
assign F[153][113] = 9'b100010000;
assign F[153][114] = 9'b100110101;
assign F[153][118] = 9'b110111100;
assign F[153][119] = 9'b110011100;
assign F[153][120] = 9'b110011100;
assign F[153][121] = 9'b110011100;
assign F[153][122] = 9'b110011100;
assign F[153][123] = 9'b110111100;
assign F[153][124] = 9'b110011100;
assign F[153][125] = 9'b110011100;
assign F[153][126] = 9'b110011100;
assign F[153][127] = 9'b110111100;
assign F[153][128] = 9'b110111100;
assign F[153][129] = 9'b110011100;
assign F[154][65] = 9'b101110101;
assign F[154][66] = 9'b100110000;
assign F[154][67] = 9'b100010100;
assign F[154][68] = 9'b100010100;
assign F[154][69] = 9'b100010100;
assign F[154][70] = 9'b100010000;
assign F[154][71] = 9'b100010000;
assign F[154][72] = 9'b100010000;
assign F[154][73] = 9'b100010000;
assign F[154][74] = 9'b100010000;
assign F[154][75] = 9'b100110000;
assign F[154][76] = 9'b100010000;
assign F[154][77] = 9'b100010001;
assign F[154][78] = 9'b110011110;
assign F[154][79] = 9'b111111100;
assign F[154][80] = 9'b110111100;
assign F[154][81] = 9'b110111100;
assign F[154][82] = 9'b110111101;
assign F[154][83] = 9'b111111100;
assign F[154][84] = 9'b110111100;
assign F[154][85] = 9'b110011100;
assign F[154][86] = 9'b110111101;
assign F[154][87] = 9'b111111100;
assign F[154][88] = 9'b110111100;
assign F[154][89] = 9'b110111100;
assign F[154][90] = 9'b110111100;
assign F[154][91] = 9'b110111100;
assign F[154][92] = 9'b110111100;
assign F[154][93] = 9'b110011100;
assign F[154][96] = 9'b101010000;
assign F[154][97] = 9'b100110100;
assign F[154][98] = 9'b100010100;
assign F[154][99] = 9'b100010100;
assign F[154][100] = 9'b100111110;
assign F[154][101] = 9'b110011111;
assign F[154][104] = 9'b101010101;
assign F[154][105] = 9'b100110100;
assign F[154][106] = 9'b100010101;
assign F[154][107] = 9'b101011110;
assign F[154][111] = 9'b100110000;
assign F[154][112] = 9'b100010100;
assign F[154][113] = 9'b100010100;
assign F[154][114] = 9'b100110101;
assign F[154][115] = 9'b101111111;
assign F[154][118] = 9'b111111100;
assign F[154][119] = 9'b110111100;
assign F[154][120] = 9'b110111100;
assign F[154][121] = 9'b110111100;
assign F[154][122] = 9'b110111100;
assign F[154][123] = 9'b110111100;
assign F[154][124] = 9'b110111100;
assign F[154][125] = 9'b111111100;
assign F[154][126] = 9'b111111100;
assign F[154][127] = 9'b111111100;
assign F[154][128] = 9'b111111100;
assign F[154][129] = 9'b110111101;
assign F[155][67] = 9'b101010101;
assign F[155][68] = 9'b100110100;
assign F[155][69] = 9'b100110001;
assign F[155][70] = 9'b100110001;
assign F[155][71] = 9'b100110000;
assign F[155][72] = 9'b100110100;
assign F[155][73] = 9'b100010100;
assign F[155][74] = 9'b100110100;
assign F[155][75] = 9'b100110100;
assign F[155][76] = 9'b100010001;
assign F[155][77] = 9'b100110001;
assign F[155][78] = 9'b110011101;
assign F[155][79] = 9'b111111100;
assign F[155][80] = 9'b110111100;
assign F[155][81] = 9'b110011100;
assign F[155][83] = 9'b111111101;
assign F[155][84] = 9'b110111100;
assign F[155][85] = 9'b110111101;
assign F[155][88] = 9'b110111100;
assign F[155][89] = 9'b110111100;
assign F[155][90] = 9'b110011100;
assign F[155][91] = 9'b110111100;
assign F[155][92] = 9'b110111100;
assign F[155][93] = 9'b110011100;
assign F[155][96] = 9'b101010101;
assign F[155][97] = 9'b100110101;
assign F[155][98] = 9'b100110000;
assign F[155][99] = 9'b100110000;
assign F[155][100] = 9'b100111110;
assign F[155][101] = 9'b110011111;
assign F[155][105] = 9'b100110101;
assign F[155][106] = 9'b101010101;
assign F[155][111] = 9'b100110001;
assign F[155][112] = 9'b100110100;
assign F[155][113] = 9'b100110000;
assign F[155][114] = 9'b100110101;
assign F[155][118] = 9'b110111100;
assign F[155][119] = 9'b110011100;
assign F[155][120] = 9'b110111100;
assign F[155][121] = 9'b110111100;
assign F[155][122] = 9'b110111100;
assign F[155][123] = 9'b110111100;
assign F[155][124] = 9'b110111100;
assign F[155][125] = 9'b110111100;
assign F[155][126] = 9'b110111100;
assign F[155][127] = 9'b110011100;
assign F[155][128] = 9'b110111100;
assign F[155][129] = 9'b111111101;
//Total de Lineas = 2184
endmodule

