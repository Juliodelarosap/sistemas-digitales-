`timescale 1ns / 1ps
module f1_principal (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (F[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= F[vcount- posy][hcount- posx][7:5];
				green <= F[vcount- posy][hcount- posx][4:2];
            blue 	<= F[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 30;
parameter RESOLUCION_Y = 75;
wire [8:0] F[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign F[1][6] = 9'b101110100;
assign F[1][7] = 9'b110010100;
assign F[1][8] = 9'b110010100;
assign F[1][9] = 9'b110010100;
assign F[1][10] = 9'b110010100;
assign F[1][11] = 9'b110010100;
assign F[1][12] = 9'b110010100;
assign F[1][13] = 9'b110010100;
assign F[1][14] = 9'b110010100;
assign F[1][15] = 9'b110010100;
assign F[1][16] = 9'b110010100;
assign F[1][17] = 9'b110010100;
assign F[1][18] = 9'b110010100;
assign F[1][19] = 9'b110010100;
assign F[1][20] = 9'b110010100;
assign F[1][21] = 9'b110010100;
assign F[1][22] = 9'b110010100;
assign F[2][2] = 9'b110001101;
assign F[2][3] = 9'b101110000;
assign F[2][4] = 9'b110010100;
assign F[2][5] = 9'b110011100;
assign F[2][6] = 9'b110011100;
assign F[2][7] = 9'b110011100;
assign F[2][8] = 9'b110011100;
assign F[2][9] = 9'b110011100;
assign F[2][10] = 9'b110011100;
assign F[2][11] = 9'b110011100;
assign F[2][12] = 9'b110011100;
assign F[2][13] = 9'b110011100;
assign F[2][14] = 9'b110011100;
assign F[2][15] = 9'b110011100;
assign F[2][16] = 9'b110011100;
assign F[2][17] = 9'b110011100;
assign F[2][18] = 9'b110011100;
assign F[2][19] = 9'b110011100;
assign F[2][20] = 9'b110011100;
assign F[2][21] = 9'b110011100;
assign F[2][22] = 9'b110011100;
assign F[2][23] = 9'b110011100;
assign F[2][24] = 9'b110010100;
assign F[2][25] = 9'b101110100;
assign F[2][26] = 9'b101101101;
assign F[2][27] = 9'b110010001;
assign F[3][2] = 9'b110001101;
assign F[3][3] = 9'b101110001;
assign F[3][4] = 9'b110011100;
assign F[3][5] = 9'b110010100;
assign F[3][6] = 9'b110010100;
assign F[3][7] = 9'b110010100;
assign F[3][8] = 9'b110010100;
assign F[3][9] = 9'b110010100;
assign F[3][10] = 9'b110010100;
assign F[3][11] = 9'b110010100;
assign F[3][12] = 9'b110010100;
assign F[3][13] = 9'b110010100;
assign F[3][14] = 9'b110010100;
assign F[3][15] = 9'b110010100;
assign F[3][16] = 9'b110010100;
assign F[3][17] = 9'b110010100;
assign F[3][18] = 9'b110010100;
assign F[3][19] = 9'b110010100;
assign F[3][20] = 9'b110010100;
assign F[3][21] = 9'b110010100;
assign F[3][22] = 9'b110010100;
assign F[3][23] = 9'b110010100;
assign F[3][24] = 9'b110011100;
assign F[3][25] = 9'b110011100;
assign F[3][26] = 9'b110010001;
assign F[3][27] = 9'b110010001;
assign F[4][2] = 9'b110010001;
assign F[4][3] = 9'b101101101;
assign F[4][4] = 9'b101001100;
assign F[4][5] = 9'b101001100;
assign F[4][6] = 9'b101001100;
assign F[4][7] = 9'b101001100;
assign F[4][8] = 9'b101001100;
assign F[4][9] = 9'b101001100;
assign F[4][10] = 9'b101001100;
assign F[4][11] = 9'b101001100;
assign F[4][12] = 9'b101001100;
assign F[4][13] = 9'b101001100;
assign F[4][14] = 9'b110010101;
assign F[4][15] = 9'b101110001;
assign F[4][16] = 9'b101001100;
assign F[4][17] = 9'b101001100;
assign F[4][18] = 9'b101001100;
assign F[4][19] = 9'b101001100;
assign F[4][20] = 9'b101001100;
assign F[4][21] = 9'b101001100;
assign F[4][22] = 9'b101001100;
assign F[4][23] = 9'b101001100;
assign F[4][24] = 9'b101001100;
assign F[4][25] = 9'b101001100;
assign F[4][26] = 9'b101101101;
assign F[4][27] = 9'b110010010;
assign F[5][2] = 9'b101001001;
assign F[5][3] = 9'b101001001;
assign F[5][4] = 9'b100100000;
assign F[5][5] = 9'b100100000;
assign F[5][6] = 9'b100100000;
assign F[5][14] = 9'b111111110;
assign F[5][15] = 9'b111111110;
assign F[5][23] = 9'b100100100;
assign F[5][24] = 9'b100100000;
assign F[5][25] = 9'b100100000;
assign F[5][26] = 9'b101001001;
assign F[5][27] = 9'b101001001;
assign F[6][1] = 9'b100100100;
assign F[6][2] = 9'b100100100;
assign F[6][3] = 9'b100100100;
assign F[6][4] = 9'b100100100;
assign F[6][5] = 9'b100100100;
assign F[6][6] = 9'b100100100;
assign F[6][7] = 9'b100100100;
assign F[6][13] = 9'b110011101;
assign F[6][14] = 9'b111111110;
assign F[6][15] = 9'b111111101;
assign F[6][16] = 9'b101110100;
assign F[6][22] = 9'b100100100;
assign F[6][23] = 9'b100100100;
assign F[6][24] = 9'b100100100;
assign F[6][25] = 9'b100100100;
assign F[6][26] = 9'b100100100;
assign F[6][27] = 9'b100100100;
assign F[6][28] = 9'b100100100;
assign F[7][1] = 9'b100100100;
assign F[7][2] = 9'b100100100;
assign F[7][3] = 9'b100100100;
assign F[7][4] = 9'b100100100;
assign F[7][5] = 9'b100100100;
assign F[7][6] = 9'b100100100;
assign F[7][7] = 9'b100100100;
assign F[7][13] = 9'b110010100;
assign F[7][14] = 9'b111111110;
assign F[7][15] = 9'b111111101;
assign F[7][16] = 9'b101110100;
assign F[7][21] = 9'b100100100;
assign F[7][22] = 9'b100100100;
assign F[7][23] = 9'b100100100;
assign F[7][24] = 9'b100100100;
assign F[7][25] = 9'b100100100;
assign F[7][26] = 9'b100100100;
assign F[7][27] = 9'b100100100;
assign F[7][28] = 9'b100100100;
assign F[8][0] = 9'b100100100;
assign F[8][1] = 9'b100100100;
assign F[8][2] = 9'b100100100;
assign F[8][3] = 9'b100100100;
assign F[8][4] = 9'b100100100;
assign F[8][5] = 9'b100100100;
assign F[8][6] = 9'b100100100;
assign F[8][7] = 9'b100100100;
assign F[8][13] = 9'b110011100;
assign F[8][14] = 9'b111111101;
assign F[8][15] = 9'b111111101;
assign F[8][16] = 9'b101110100;
assign F[8][21] = 9'b100100100;
assign F[8][22] = 9'b100100100;
assign F[8][23] = 9'b100100100;
assign F[8][24] = 9'b100100100;
assign F[8][25] = 9'b100100100;
assign F[8][26] = 9'b100100100;
assign F[8][27] = 9'b100100100;
assign F[8][28] = 9'b100100100;
assign F[9][0] = 9'b100100100;
assign F[9][1] = 9'b100100100;
assign F[9][2] = 9'b100100100;
assign F[9][3] = 9'b100100100;
assign F[9][4] = 9'b100100100;
assign F[9][5] = 9'b100100100;
assign F[9][6] = 9'b100100100;
assign F[9][7] = 9'b100100100;
assign F[9][8] = 9'b100100100;
assign F[9][12] = 9'b101001100;
assign F[9][13] = 9'b110011100;
assign F[9][14] = 9'b111111101;
assign F[9][15] = 9'b110111101;
assign F[9][16] = 9'b101110100;
assign F[9][17] = 9'b100101000;
assign F[9][21] = 9'b100100100;
assign F[9][22] = 9'b100100100;
assign F[9][23] = 9'b100100100;
assign F[9][24] = 9'b100100100;
assign F[9][25] = 9'b100100100;
assign F[9][26] = 9'b100100100;
assign F[9][27] = 9'b100100100;
assign F[9][28] = 9'b100100100;
assign F[10][0] = 9'b100100100;
assign F[10][1] = 9'b100100100;
assign F[10][2] = 9'b100100100;
assign F[10][3] = 9'b100100100;
assign F[10][4] = 9'b100100100;
assign F[10][5] = 9'b100100100;
assign F[10][6] = 9'b100100100;
assign F[10][7] = 9'b100100100;
assign F[10][8] = 9'b100100100;
assign F[10][9] = 9'b100100100;
assign F[10][10] = 9'b100100100;
assign F[10][11] = 9'b100100000;
assign F[10][12] = 9'b101001100;
assign F[10][13] = 9'b110011100;
assign F[10][14] = 9'b111111101;
assign F[10][15] = 9'b110111101;
assign F[10][16] = 9'b101110100;
assign F[10][17] = 9'b100101000;
assign F[10][18] = 9'b100100100;
assign F[10][19] = 9'b100100100;
assign F[10][20] = 9'b100100100;
assign F[10][21] = 9'b100100100;
assign F[10][22] = 9'b100100100;
assign F[10][23] = 9'b100100100;
assign F[10][24] = 9'b100100100;
assign F[10][25] = 9'b100100100;
assign F[10][26] = 9'b100100100;
assign F[10][27] = 9'b100100100;
assign F[10][28] = 9'b100100100;
assign F[10][29] = 9'b100100100;
assign F[11][0] = 9'b100100100;
assign F[11][1] = 9'b100100100;
assign F[11][2] = 9'b100100100;
assign F[11][3] = 9'b100100100;
assign F[11][4] = 9'b100100100;
assign F[11][5] = 9'b100100100;
assign F[11][6] = 9'b100100100;
assign F[11][7] = 9'b100100100;
assign F[11][8] = 9'b100100100;
assign F[11][12] = 9'b101110100;
assign F[11][13] = 9'b110011100;
assign F[11][14] = 9'b111111101;
assign F[11][15] = 9'b110111101;
assign F[11][16] = 9'b101110100;
assign F[11][21] = 9'b100100100;
assign F[11][22] = 9'b100100100;
assign F[11][23] = 9'b100100100;
assign F[11][24] = 9'b100100100;
assign F[11][25] = 9'b100100100;
assign F[11][26] = 9'b100100100;
assign F[11][27] = 9'b100100100;
assign F[11][28] = 9'b100100100;
assign F[11][29] = 9'b100100100;
assign F[12][0] = 9'b100100100;
assign F[12][1] = 9'b100100100;
assign F[12][2] = 9'b100100100;
assign F[12][3] = 9'b100100100;
assign F[12][4] = 9'b100100100;
assign F[12][5] = 9'b100100100;
assign F[12][6] = 9'b100100100;
assign F[12][7] = 9'b100100100;
assign F[12][8] = 9'b100100100;
assign F[12][10] = 9'b100100100;
assign F[12][11] = 9'b100000000;
assign F[12][12] = 9'b101001100;
assign F[12][13] = 9'b110011100;
assign F[12][14] = 9'b111111101;
assign F[12][15] = 9'b110111101;
assign F[12][16] = 9'b101110100;
assign F[12][17] = 9'b100101000;
assign F[12][18] = 9'b100100000;
assign F[12][19] = 9'b100100100;
assign F[12][21] = 9'b100100100;
assign F[12][22] = 9'b100100100;
assign F[12][23] = 9'b100100100;
assign F[12][24] = 9'b100100100;
assign F[12][25] = 9'b100100100;
assign F[12][26] = 9'b100100100;
assign F[12][27] = 9'b100100100;
assign F[12][28] = 9'b100100100;
assign F[12][29] = 9'b100100100;
assign F[13][0] = 9'b100100100;
assign F[13][1] = 9'b100100100;
assign F[13][2] = 9'b100100100;
assign F[13][3] = 9'b100100100;
assign F[13][4] = 9'b100100100;
assign F[13][5] = 9'b100100100;
assign F[13][6] = 9'b100100100;
assign F[13][7] = 9'b100100100;
assign F[13][8] = 9'b100100100;
assign F[13][9] = 9'b100100100;
assign F[13][10] = 9'b100100100;
assign F[13][12] = 9'b101110100;
assign F[13][13] = 9'b110011100;
assign F[13][14] = 9'b111111101;
assign F[13][15] = 9'b110111101;
assign F[13][16] = 9'b101110100;
assign F[13][19] = 9'b100100100;
assign F[13][20] = 9'b100100100;
assign F[13][21] = 9'b100100100;
assign F[13][22] = 9'b100100100;
assign F[13][23] = 9'b100100100;
assign F[13][24] = 9'b100100100;
assign F[13][25] = 9'b100100100;
assign F[13][26] = 9'b100100100;
assign F[13][27] = 9'b100100100;
assign F[13][28] = 9'b100100100;
assign F[14][0] = 9'b100100100;
assign F[14][1] = 9'b100100100;
assign F[14][2] = 9'b100100100;
assign F[14][3] = 9'b100100100;
assign F[14][4] = 9'b100100100;
assign F[14][5] = 9'b100100100;
assign F[14][6] = 9'b100100100;
assign F[14][7] = 9'b100100100;
assign F[14][12] = 9'b101110100;
assign F[14][13] = 9'b110011100;
assign F[14][14] = 9'b111111101;
assign F[14][15] = 9'b110111101;
assign F[14][16] = 9'b101110100;
assign F[14][21] = 9'b100100100;
assign F[14][22] = 9'b100100100;
assign F[14][23] = 9'b100100100;
assign F[14][24] = 9'b100100100;
assign F[14][25] = 9'b100100100;
assign F[14][26] = 9'b100100100;
assign F[14][27] = 9'b100100100;
assign F[14][28] = 9'b100100100;
assign F[15][1] = 9'b100100100;
assign F[15][2] = 9'b100100100;
assign F[15][3] = 9'b100100100;
assign F[15][4] = 9'b100100100;
assign F[15][5] = 9'b100100100;
assign F[15][6] = 9'b100100100;
assign F[15][7] = 9'b100100100;
assign F[15][12] = 9'b101110100;
assign F[15][13] = 9'b110011100;
assign F[15][14] = 9'b111111101;
assign F[15][15] = 9'b110111101;
assign F[15][16] = 9'b101110100;
assign F[15][17] = 9'b101110100;
assign F[15][21] = 9'b100100100;
assign F[15][22] = 9'b100100100;
assign F[15][23] = 9'b100100100;
assign F[15][24] = 9'b100100100;
assign F[15][25] = 9'b100100100;
assign F[15][26] = 9'b100100100;
assign F[15][27] = 9'b100100100;
assign F[15][28] = 9'b100100100;
assign F[16][1] = 9'b100100100;
assign F[16][2] = 9'b100100100;
assign F[16][3] = 9'b100100100;
assign F[16][4] = 9'b100100100;
assign F[16][5] = 9'b100100100;
assign F[16][6] = 9'b100100100;
assign F[16][7] = 9'b100100100;
assign F[16][12] = 9'b101110100;
assign F[16][13] = 9'b110011100;
assign F[16][14] = 9'b111111101;
assign F[16][15] = 9'b110111101;
assign F[16][16] = 9'b101111100;
assign F[16][17] = 9'b101110100;
assign F[16][22] = 9'b100100100;
assign F[16][23] = 9'b100100100;
assign F[16][24] = 9'b100100100;
assign F[16][25] = 9'b100100100;
assign F[16][26] = 9'b100100100;
assign F[16][27] = 9'b100100100;
assign F[16][28] = 9'b100100100;
assign F[17][2] = 9'b100100100;
assign F[17][3] = 9'b100100100;
assign F[17][4] = 9'b100100100;
assign F[17][5] = 9'b100100100;
assign F[17][6] = 9'b100100100;
assign F[17][12] = 9'b101110100;
assign F[17][13] = 9'b110011100;
assign F[17][14] = 9'b111111101;
assign F[17][15] = 9'b110111101;
assign F[17][16] = 9'b101111100;
assign F[17][17] = 9'b101110100;
assign F[17][22] = 9'b100100100;
assign F[17][23] = 9'b100100100;
assign F[17][24] = 9'b100100100;
assign F[17][25] = 9'b100100100;
assign F[17][26] = 9'b100100100;
assign F[17][27] = 9'b100100100;
assign F[18][12] = 9'b101110100;
assign F[18][13] = 9'b110011100;
assign F[18][14] = 9'b111111101;
assign F[18][15] = 9'b110111101;
assign F[18][16] = 9'b101111100;
assign F[18][17] = 9'b101110100;
assign F[19][12] = 9'b101110100;
assign F[19][13] = 9'b110011100;
assign F[19][14] = 9'b111111101;
assign F[19][15] = 9'b110111101;
assign F[19][16] = 9'b101111100;
assign F[19][17] = 9'b101110100;
assign F[20][12] = 9'b101110100;
assign F[20][13] = 9'b110011100;
assign F[20][14] = 9'b111111101;
assign F[20][15] = 9'b110111101;
assign F[20][16] = 9'b101111100;
assign F[20][17] = 9'b101110100;
assign F[21][12] = 9'b101110100;
assign F[21][13] = 9'b110011100;
assign F[21][14] = 9'b111111101;
assign F[21][15] = 9'b110111101;
assign F[21][16] = 9'b101111100;
assign F[21][17] = 9'b101110100;
assign F[22][12] = 9'b101110100;
assign F[22][13] = 9'b110011100;
assign F[22][14] = 9'b111111101;
assign F[22][15] = 9'b110111101;
assign F[22][16] = 9'b101110100;
assign F[22][17] = 9'b101110100;
assign F[23][12] = 9'b101110100;
assign F[23][13] = 9'b110010100;
assign F[23][14] = 9'b111111101;
assign F[23][15] = 9'b110111101;
assign F[23][16] = 9'b101110100;
assign F[23][17] = 9'b101110100;
assign F[24][9] = 9'b101010000;
assign F[24][10] = 9'b101010000;
assign F[24][11] = 9'b101110000;
assign F[24][12] = 9'b101110100;
assign F[24][13] = 9'b110010100;
assign F[24][14] = 9'b111111101;
assign F[24][15] = 9'b110111101;
assign F[24][16] = 9'b101110100;
assign F[24][17] = 9'b101110100;
assign F[24][18] = 9'b101010000;
assign F[24][19] = 9'b101010000;
assign F[24][20] = 9'b101010000;
assign F[25][7] = 9'b101111100;
assign F[25][8] = 9'b101010000;
assign F[25][9] = 9'b100101100;
assign F[25][10] = 9'b100101000;
assign F[25][11] = 9'b101010000;
assign F[25][12] = 9'b101110100;
assign F[25][13] = 9'b110010100;
assign F[25][14] = 9'b111111101;
assign F[25][15] = 9'b110111101;
assign F[25][16] = 9'b101110100;
assign F[25][17] = 9'b101110100;
assign F[25][18] = 9'b101001100;
assign F[25][19] = 9'b100101100;
assign F[25][20] = 9'b101001100;
assign F[25][21] = 9'b101110000;
assign F[26][7] = 9'b101110100;
assign F[26][8] = 9'b101110100;
assign F[26][9] = 9'b101001100;
assign F[26][10] = 9'b101001100;
assign F[26][11] = 9'b101010000;
assign F[26][12] = 9'b101110100;
assign F[26][13] = 9'b110010100;
assign F[26][14] = 9'b111111101;
assign F[26][15] = 9'b110111101;
assign F[26][16] = 9'b101110100;
assign F[26][17] = 9'b101110100;
assign F[26][18] = 9'b101001100;
assign F[26][19] = 9'b101001100;
assign F[26][20] = 9'b101001100;
assign F[26][21] = 9'b101111100;
assign F[26][22] = 9'b101110100;
assign F[27][7] = 9'b101110100;
assign F[27][8] = 9'b101110100;
assign F[27][9] = 9'b101110100;
assign F[27][10] = 9'b101110100;
assign F[27][11] = 9'b101110100;
assign F[27][12] = 9'b101110100;
assign F[27][13] = 9'b110010100;
assign F[27][14] = 9'b111111101;
assign F[27][15] = 9'b110111101;
assign F[27][16] = 9'b101110100;
assign F[27][17] = 9'b101110100;
assign F[27][18] = 9'b101110100;
assign F[27][19] = 9'b101110100;
assign F[27][20] = 9'b101110100;
assign F[27][21] = 9'b101110100;
assign F[27][22] = 9'b101110100;
assign F[28][7] = 9'b101110100;
assign F[28][8] = 9'b101110100;
assign F[28][9] = 9'b101001100;
assign F[28][10] = 9'b101110000;
assign F[28][11] = 9'b101110100;
assign F[28][12] = 9'b101110100;
assign F[28][13] = 9'b110010100;
assign F[28][14] = 9'b111111101;
assign F[28][15] = 9'b110111101;
assign F[28][16] = 9'b101110100;
assign F[28][17] = 9'b101110100;
assign F[28][18] = 9'b101110100;
assign F[28][19] = 9'b101001100;
assign F[28][20] = 9'b101010000;
assign F[28][21] = 9'b101111100;
assign F[28][22] = 9'b101110100;
assign F[29][7] = 9'b101110100;
assign F[29][8] = 9'b101110100;
assign F[29][9] = 9'b101001100;
assign F[29][10] = 9'b101001100;
assign F[29][11] = 9'b101110100;
assign F[29][12] = 9'b101110100;
assign F[29][13] = 9'b110010100;
assign F[29][14] = 9'b111111101;
assign F[29][15] = 9'b110111101;
assign F[29][16] = 9'b101110100;
assign F[29][17] = 9'b101110100;
assign F[29][18] = 9'b101110000;
assign F[29][19] = 9'b101001000;
assign F[29][20] = 9'b101010000;
assign F[29][21] = 9'b101111100;
assign F[29][22] = 9'b101110100;
assign F[30][7] = 9'b101110000;
assign F[30][8] = 9'b101110100;
assign F[30][9] = 9'b101001100;
assign F[30][10] = 9'b101001100;
assign F[30][11] = 9'b101110100;
assign F[30][12] = 9'b101110100;
assign F[30][13] = 9'b110011100;
assign F[30][14] = 9'b111111110;
assign F[30][15] = 9'b111111101;
assign F[30][16] = 9'b101110100;
assign F[30][17] = 9'b101110100;
assign F[30][18] = 9'b101110000;
assign F[30][19] = 9'b101001000;
assign F[30][20] = 9'b101010000;
assign F[30][21] = 9'b101111100;
assign F[30][22] = 9'b101110000;
assign F[31][7] = 9'b101110000;
assign F[31][8] = 9'b101110100;
assign F[31][9] = 9'b101001100;
assign F[31][10] = 9'b101001100;
assign F[31][11] = 9'b101110100;
assign F[31][12] = 9'b101110100;
assign F[31][13] = 9'b101110000;
assign F[31][14] = 9'b110010101;
assign F[31][15] = 9'b110010101;
assign F[31][16] = 9'b101110000;
assign F[31][17] = 9'b101110100;
assign F[31][18] = 9'b101110000;
assign F[31][19] = 9'b101001000;
assign F[31][20] = 9'b101010000;
assign F[31][21] = 9'b101111100;
assign F[31][22] = 9'b101001100;
assign F[32][7] = 9'b101001100;
assign F[32][8] = 9'b101111100;
assign F[32][9] = 9'b101001100;
assign F[32][10] = 9'b101001100;
assign F[32][11] = 9'b101110100;
assign F[32][12] = 9'b101010000;
assign F[32][13] = 9'b100101000;
assign F[32][14] = 9'b100101000;
assign F[32][15] = 9'b100101000;
assign F[32][16] = 9'b101001100;
assign F[32][17] = 9'b101110000;
assign F[32][18] = 9'b101110000;
assign F[32][19] = 9'b101001000;
assign F[32][20] = 9'b101110000;
assign F[32][21] = 9'b101111100;
assign F[32][22] = 9'b101001000;
assign F[33][7] = 9'b101001100;
assign F[33][8] = 9'b101110100;
assign F[33][9] = 9'b101110000;
assign F[33][10] = 9'b101010000;
assign F[33][11] = 9'b101110100;
assign F[33][12] = 9'b101010000;
assign F[33][13] = 9'b100101000;
assign F[33][14] = 9'b100101100;
assign F[33][15] = 9'b100101100;
assign F[33][16] = 9'b100101100;
assign F[33][17] = 9'b101110000;
assign F[33][18] = 9'b101110000;
assign F[33][19] = 9'b101010000;
assign F[33][20] = 9'b101110100;
assign F[33][21] = 9'b101110100;
assign F[33][22] = 9'b101001000;
assign F[34][7] = 9'b101001100;
assign F[34][8] = 9'b101110100;
assign F[34][9] = 9'b101110100;
assign F[34][10] = 9'b101110100;
assign F[34][11] = 9'b101110100;
assign F[34][12] = 9'b101010000;
assign F[34][13] = 9'b100101000;
assign F[34][14] = 9'b100101100;
assign F[34][15] = 9'b100101100;
assign F[34][16] = 9'b101001100;
assign F[34][17] = 9'b101110000;
assign F[34][18] = 9'b101110100;
assign F[34][19] = 9'b101110100;
assign F[34][20] = 9'b101110100;
assign F[34][21] = 9'b101110100;
assign F[34][22] = 9'b101001000;
assign F[35][7] = 9'b101001000;
assign F[35][8] = 9'b101110100;
assign F[35][9] = 9'b101110100;
assign F[35][10] = 9'b101110100;
assign F[35][11] = 9'b101110100;
assign F[35][12] = 9'b101010000;
assign F[35][13] = 9'b100101000;
assign F[35][14] = 9'b100101100;
assign F[35][15] = 9'b100101100;
assign F[35][16] = 9'b101001100;
assign F[35][17] = 9'b101110000;
assign F[35][18] = 9'b101110100;
assign F[35][19] = 9'b101110100;
assign F[35][20] = 9'b101110100;
assign F[35][21] = 9'b101110000;
assign F[35][22] = 9'b100100100;
assign F[36][7] = 9'b101001000;
assign F[36][8] = 9'b101110100;
assign F[36][9] = 9'b101110100;
assign F[36][10] = 9'b101110100;
assign F[36][11] = 9'b101110100;
assign F[36][12] = 9'b101010000;
assign F[36][13] = 9'b100101000;
assign F[36][14] = 9'b100101000;
assign F[36][15] = 9'b100101000;
assign F[36][16] = 9'b100101100;
assign F[36][17] = 9'b101110000;
assign F[36][18] = 9'b101110100;
assign F[36][19] = 9'b101110100;
assign F[36][20] = 9'b101110100;
assign F[36][21] = 9'b101110000;
assign F[36][22] = 9'b100100100;
assign F[37][7] = 9'b101001000;
assign F[37][8] = 9'b101110100;
assign F[37][9] = 9'b101110100;
assign F[37][10] = 9'b101110100;
assign F[37][11] = 9'b101110100;
assign F[37][12] = 9'b101010000;
assign F[37][13] = 9'b100101000;
assign F[37][14] = 9'b101001100;
assign F[37][15] = 9'b101001100;
assign F[37][16] = 9'b100101100;
assign F[37][17] = 9'b101110000;
assign F[37][18] = 9'b101110100;
assign F[37][19] = 9'b101110100;
assign F[37][20] = 9'b101110100;
assign F[37][21] = 9'b101110000;
assign F[37][22] = 9'b100100100;
assign F[38][7] = 9'b100100100;
assign F[38][8] = 9'b101110000;
assign F[38][9] = 9'b101110100;
assign F[38][10] = 9'b101110100;
assign F[38][11] = 9'b101110100;
assign F[38][12] = 9'b101110000;
assign F[38][13] = 9'b101110000;
assign F[38][14] = 9'b101110100;
assign F[38][15] = 9'b101110100;
assign F[38][16] = 9'b101110000;
assign F[38][17] = 9'b101110000;
assign F[38][18] = 9'b101110100;
assign F[38][19] = 9'b101110100;
assign F[38][20] = 9'b101110100;
assign F[38][21] = 9'b101001100;
assign F[38][22] = 9'b100100100;
assign F[39][7] = 9'b100100100;
assign F[39][8] = 9'b101110000;
assign F[39][9] = 9'b101110100;
assign F[39][10] = 9'b101110100;
assign F[39][11] = 9'b101110100;
assign F[39][12] = 9'b101110100;
assign F[39][13] = 9'b110010100;
assign F[39][14] = 9'b110010100;
assign F[39][15] = 9'b110010100;
assign F[39][16] = 9'b101110100;
assign F[39][17] = 9'b101110100;
assign F[39][18] = 9'b101110100;
assign F[39][19] = 9'b101110100;
assign F[39][20] = 9'b101110100;
assign F[39][21] = 9'b101001100;
assign F[39][22] = 9'b100100100;
assign F[40][7] = 9'b100100100;
assign F[40][8] = 9'b101110000;
assign F[40][9] = 9'b101110100;
assign F[40][10] = 9'b101110100;
assign F[40][11] = 9'b101110100;
assign F[40][12] = 9'b101110100;
assign F[40][13] = 9'b101110100;
assign F[40][14] = 9'b101110100;
assign F[40][15] = 9'b110010100;
assign F[40][16] = 9'b101110100;
assign F[40][17] = 9'b101110100;
assign F[40][18] = 9'b101110100;
assign F[40][19] = 9'b101110100;
assign F[40][20] = 9'b101110100;
assign F[40][21] = 9'b101001100;
assign F[40][22] = 9'b100100100;
assign F[41][7] = 9'b100100100;
assign F[41][8] = 9'b101001100;
assign F[41][9] = 9'b101110100;
assign F[41][10] = 9'b101110100;
assign F[41][11] = 9'b101110100;
assign F[41][12] = 9'b101110100;
assign F[41][13] = 9'b101110100;
assign F[41][14] = 9'b101110100;
assign F[41][15] = 9'b110010100;
assign F[41][16] = 9'b101110100;
assign F[41][17] = 9'b101110100;
assign F[41][18] = 9'b101110100;
assign F[41][19] = 9'b101110100;
assign F[41][20] = 9'b101110100;
assign F[41][21] = 9'b101001000;
assign F[41][22] = 9'b100100100;
assign F[42][7] = 9'b100100100;
assign F[42][8] = 9'b101001100;
assign F[42][9] = 9'b101110100;
assign F[42][10] = 9'b101110100;
assign F[42][11] = 9'b101110100;
assign F[42][12] = 9'b101110100;
assign F[42][13] = 9'b110010100;
assign F[42][14] = 9'b101110100;
assign F[42][15] = 9'b110010100;
assign F[42][16] = 9'b101110100;
assign F[42][17] = 9'b101110100;
assign F[42][18] = 9'b101110100;
assign F[42][19] = 9'b101110100;
assign F[42][20] = 9'b101110100;
assign F[42][21] = 9'b101001000;
assign F[42][22] = 9'b100100100;
assign F[43][7] = 9'b100100100;
assign F[43][8] = 9'b101001100;
assign F[43][9] = 9'b101110100;
assign F[43][10] = 9'b101110100;
assign F[43][11] = 9'b101110100;
assign F[43][12] = 9'b101110100;
assign F[43][13] = 9'b110010100;
assign F[43][14] = 9'b101110100;
assign F[43][15] = 9'b110010100;
assign F[43][16] = 9'b101110100;
assign F[43][17] = 9'b101110100;
assign F[43][18] = 9'b101110100;
assign F[43][19] = 9'b101110100;
assign F[43][20] = 9'b101110100;
assign F[43][21] = 9'b101001000;
assign F[43][22] = 9'b100100100;
assign F[44][7] = 9'b100100100;
assign F[44][8] = 9'b101001000;
assign F[44][9] = 9'b101110100;
assign F[44][10] = 9'b101110100;
assign F[44][11] = 9'b101110100;
assign F[44][12] = 9'b101110100;
assign F[44][13] = 9'b110010100;
assign F[44][14] = 9'b101110100;
assign F[44][15] = 9'b110010100;
assign F[44][16] = 9'b101110100;
assign F[44][17] = 9'b101110100;
assign F[44][18] = 9'b101110100;
assign F[44][19] = 9'b101110100;
assign F[44][20] = 9'b101110000;
assign F[44][21] = 9'b101001000;
assign F[44][22] = 9'b100100100;
assign F[45][7] = 9'b100100100;
assign F[45][8] = 9'b101001000;
assign F[45][9] = 9'b101110100;
assign F[45][10] = 9'b101110100;
assign F[45][11] = 9'b101110100;
assign F[45][12] = 9'b101110100;
assign F[45][13] = 9'b110010100;
assign F[45][14] = 9'b101110100;
assign F[45][15] = 9'b110010100;
assign F[45][16] = 9'b101110100;
assign F[45][17] = 9'b101110100;
assign F[45][18] = 9'b101110100;
assign F[45][19] = 9'b101110100;
assign F[45][20] = 9'b101110000;
assign F[45][21] = 9'b100100100;
assign F[45][22] = 9'b100100100;
assign F[46][7] = 9'b100100100;
assign F[46][8] = 9'b101001000;
assign F[46][9] = 9'b101110100;
assign F[46][10] = 9'b101110100;
assign F[46][11] = 9'b101110100;
assign F[46][12] = 9'b101110100;
assign F[46][13] = 9'b110010100;
assign F[46][14] = 9'b101110100;
assign F[46][15] = 9'b101110100;
assign F[46][16] = 9'b101110100;
assign F[46][17] = 9'b101110100;
assign F[46][18] = 9'b101110100;
assign F[46][19] = 9'b101110100;
assign F[46][20] = 9'b101110000;
assign F[46][21] = 9'b100100100;
assign F[46][22] = 9'b100100100;
assign F[47][7] = 9'b100100100;
assign F[47][8] = 9'b100101000;
assign F[47][9] = 9'b101110000;
assign F[47][10] = 9'b101110100;
assign F[47][11] = 9'b101110100;
assign F[47][12] = 9'b101110100;
assign F[47][13] = 9'b110010100;
assign F[47][14] = 9'b101110100;
assign F[47][15] = 9'b101110100;
assign F[47][16] = 9'b101110100;
assign F[47][17] = 9'b101110100;
assign F[47][18] = 9'b101110100;
assign F[47][19] = 9'b101110100;
assign F[47][20] = 9'b101001100;
assign F[47][21] = 9'b100100100;
assign F[47][22] = 9'b100100100;
assign F[48][7] = 9'b100100100;
assign F[48][8] = 9'b100100100;
assign F[48][9] = 9'b101110000;
assign F[48][10] = 9'b101110100;
assign F[48][11] = 9'b101110100;
assign F[48][12] = 9'b101110100;
assign F[48][13] = 9'b110010100;
assign F[48][14] = 9'b101110100;
assign F[48][15] = 9'b101110100;
assign F[48][16] = 9'b101110100;
assign F[48][17] = 9'b101110100;
assign F[48][18] = 9'b101110100;
assign F[48][19] = 9'b101110100;
assign F[48][20] = 9'b101001100;
assign F[48][21] = 9'b100100100;
assign F[48][22] = 9'b100100100;
assign F[49][7] = 9'b100100100;
assign F[49][8] = 9'b100100100;
assign F[49][9] = 9'b101110000;
assign F[49][10] = 9'b101110100;
assign F[49][11] = 9'b101110100;
assign F[49][12] = 9'b101110100;
assign F[49][13] = 9'b110010100;
assign F[49][14] = 9'b101110100;
assign F[49][15] = 9'b101110100;
assign F[49][16] = 9'b101110100;
assign F[49][17] = 9'b101110100;
assign F[49][18] = 9'b101110100;
assign F[49][19] = 9'b101110100;
assign F[49][20] = 9'b101001100;
assign F[49][21] = 9'b100100100;
assign F[49][22] = 9'b100100100;
assign F[50][7] = 9'b100100100;
assign F[50][8] = 9'b100100100;
assign F[50][9] = 9'b101001100;
assign F[50][10] = 9'b101110100;
assign F[50][11] = 9'b101110100;
assign F[50][12] = 9'b101110100;
assign F[50][13] = 9'b110010100;
assign F[50][14] = 9'b101110100;
assign F[50][15] = 9'b101110100;
assign F[50][16] = 9'b110010100;
assign F[50][17] = 9'b101110100;
assign F[50][18] = 9'b101110100;
assign F[50][19] = 9'b101110100;
assign F[50][20] = 9'b101001000;
assign F[50][21] = 9'b100100100;
assign F[50][22] = 9'b100100100;
assign F[51][7] = 9'b100100100;
assign F[51][8] = 9'b100100100;
assign F[51][9] = 9'b101001100;
assign F[51][10] = 9'b101110100;
assign F[51][11] = 9'b101110100;
assign F[51][12] = 9'b101110100;
assign F[51][13] = 9'b110010100;
assign F[51][14] = 9'b101110100;
assign F[51][15] = 9'b101110100;
assign F[51][16] = 9'b110010100;
assign F[51][17] = 9'b101110100;
assign F[51][18] = 9'b101110100;
assign F[51][19] = 9'b101110100;
assign F[51][20] = 9'b101001000;
assign F[51][21] = 9'b100100100;
assign F[51][22] = 9'b100100100;
assign F[52][7] = 9'b100100100;
assign F[52][8] = 9'b100100100;
assign F[52][9] = 9'b101001100;
assign F[52][10] = 9'b101110100;
assign F[52][11] = 9'b101110100;
assign F[52][12] = 9'b101110100;
assign F[52][13] = 9'b110010100;
assign F[52][14] = 9'b101110100;
assign F[52][15] = 9'b101110100;
assign F[52][16] = 9'b110010100;
assign F[52][17] = 9'b101110100;
assign F[52][18] = 9'b101110100;
assign F[52][19] = 9'b101110100;
assign F[52][20] = 9'b101001000;
assign F[52][21] = 9'b100100100;
assign F[52][22] = 9'b100100100;
assign F[53][7] = 9'b100100100;
assign F[53][8] = 9'b100100100;
assign F[53][9] = 9'b101001000;
assign F[53][10] = 9'b101110100;
assign F[53][11] = 9'b101110100;
assign F[53][12] = 9'b101110100;
assign F[53][13] = 9'b110010100;
assign F[53][14] = 9'b101110100;
assign F[53][15] = 9'b101110100;
assign F[53][16] = 9'b110010100;
assign F[53][17] = 9'b101110100;
assign F[53][18] = 9'b101110100;
assign F[53][19] = 9'b101110000;
assign F[53][20] = 9'b100101000;
assign F[53][21] = 9'b100100100;
assign F[53][22] = 9'b100100100;
assign F[54][7] = 9'b100100100;
assign F[54][8] = 9'b100100100;
assign F[54][9] = 9'b101001000;
assign F[54][10] = 9'b101110100;
assign F[54][11] = 9'b101110100;
assign F[54][12] = 9'b101110100;
assign F[54][13] = 9'b110010100;
assign F[54][14] = 9'b101110100;
assign F[54][15] = 9'b101110100;
assign F[54][16] = 9'b110010100;
assign F[54][17] = 9'b101110100;
assign F[54][18] = 9'b101110100;
assign F[54][19] = 9'b101110000;
assign F[54][20] = 9'b100100100;
assign F[54][21] = 9'b100100100;
assign F[54][22] = 9'b100100100;
assign F[55][7] = 9'b100100100;
assign F[55][8] = 9'b100100100;
assign F[55][9] = 9'b101001000;
assign F[55][10] = 9'b101110100;
assign F[55][11] = 9'b101110100;
assign F[55][12] = 9'b101110100;
assign F[55][13] = 9'b110010100;
assign F[55][14] = 9'b110010100;
assign F[55][15] = 9'b110010100;
assign F[55][16] = 9'b110010100;
assign F[55][17] = 9'b101110100;
assign F[55][18] = 9'b101110100;
assign F[55][19] = 9'b101110000;
assign F[55][20] = 9'b100100100;
assign F[55][21] = 9'b100100100;
assign F[55][22] = 9'b100100100;
assign F[55][24] = 9'b100100100;
assign F[56][1] = 9'b100100100;
assign F[56][2] = 9'b100100100;
assign F[56][3] = 9'b100100100;
assign F[56][4] = 9'b100100100;
assign F[56][5] = 9'b100100100;
assign F[56][6] = 9'b101001100;
assign F[56][7] = 9'b101001100;
assign F[56][8] = 9'b101001100;
assign F[56][9] = 9'b101001100;
assign F[56][10] = 9'b101001100;
assign F[56][11] = 9'b101010000;
assign F[56][12] = 9'b101010000;
assign F[56][13] = 9'b101010000;
assign F[56][14] = 9'b101010000;
assign F[56][15] = 9'b101010000;
assign F[56][16] = 9'b101010000;
assign F[56][17] = 9'b101001100;
assign F[56][18] = 9'b101010000;
assign F[56][19] = 9'b101001100;
assign F[56][20] = 9'b101001100;
assign F[56][21] = 9'b101001100;
assign F[56][22] = 9'b101001100;
assign F[56][23] = 9'b101001100;
assign F[56][24] = 9'b100100100;
assign F[56][25] = 9'b100100100;
assign F[56][26] = 9'b100100100;
assign F[56][27] = 9'b100100100;
assign F[56][28] = 9'b100100100;
assign F[57][0] = 9'b100100100;
assign F[57][1] = 9'b100100100;
assign F[57][2] = 9'b100100100;
assign F[57][3] = 9'b100100100;
assign F[57][4] = 9'b100100100;
assign F[57][5] = 9'b100101000;
assign F[57][6] = 9'b101010000;
assign F[57][7] = 9'b101001100;
assign F[57][8] = 9'b101001100;
assign F[57][9] = 9'b101001100;
assign F[57][10] = 9'b101001100;
assign F[57][11] = 9'b101001100;
assign F[57][12] = 9'b101001100;
assign F[57][13] = 9'b101001100;
assign F[57][14] = 9'b101001100;
assign F[57][15] = 9'b101001100;
assign F[57][16] = 9'b101001100;
assign F[57][17] = 9'b101001100;
assign F[57][18] = 9'b101001100;
assign F[57][19] = 9'b101001100;
assign F[57][20] = 9'b101001100;
assign F[57][21] = 9'b101001100;
assign F[57][22] = 9'b101010000;
assign F[57][23] = 9'b101001100;
assign F[57][24] = 9'b100100100;
assign F[57][25] = 9'b100100100;
assign F[57][26] = 9'b100100100;
assign F[57][27] = 9'b100100100;
assign F[57][28] = 9'b100100100;
assign F[57][29] = 9'b100100100;
assign F[58][0] = 9'b100100100;
assign F[58][1] = 9'b100100100;
assign F[58][2] = 9'b100100100;
assign F[58][3] = 9'b100100100;
assign F[58][4] = 9'b100100100;
assign F[58][5] = 9'b100100100;
assign F[58][6] = 9'b101001100;
assign F[58][7] = 9'b101001100;
assign F[58][8] = 9'b101001100;
assign F[58][9] = 9'b101001100;
assign F[58][10] = 9'b101001100;
assign F[58][11] = 9'b101001100;
assign F[58][12] = 9'b101001100;
assign F[58][13] = 9'b101001100;
assign F[58][14] = 9'b101001100;
assign F[58][15] = 9'b101001100;
assign F[58][16] = 9'b101001100;
assign F[58][17] = 9'b101001100;
assign F[58][18] = 9'b101001100;
assign F[58][19] = 9'b101001100;
assign F[58][20] = 9'b101001100;
assign F[58][21] = 9'b101001100;
assign F[58][22] = 9'b101001100;
assign F[58][23] = 9'b101001100;
assign F[58][24] = 9'b100100100;
assign F[58][25] = 9'b100100100;
assign F[58][26] = 9'b100100100;
assign F[58][27] = 9'b100100100;
assign F[58][28] = 9'b100100100;
assign F[58][29] = 9'b100100100;
assign F[59][0] = 9'b100100100;
assign F[59][1] = 9'b100100100;
assign F[59][2] = 9'b100100100;
assign F[59][3] = 9'b100100100;
assign F[59][4] = 9'b100100100;
assign F[59][5] = 9'b100100100;
assign F[59][6] = 9'b101001100;
assign F[59][7] = 9'b101001100;
assign F[59][8] = 9'b101001100;
assign F[59][9] = 9'b101001100;
assign F[59][10] = 9'b101001100;
assign F[59][11] = 9'b101001100;
assign F[59][12] = 9'b101001100;
assign F[59][13] = 9'b101001100;
assign F[59][14] = 9'b101001100;
assign F[59][15] = 9'b101001100;
assign F[59][16] = 9'b101001100;
assign F[59][17] = 9'b101001100;
assign F[59][18] = 9'b101001100;
assign F[59][19] = 9'b101001100;
assign F[59][20] = 9'b101001100;
assign F[59][21] = 9'b101001100;
assign F[59][22] = 9'b101001100;
assign F[59][23] = 9'b101001100;
assign F[59][24] = 9'b100100100;
assign F[59][25] = 9'b100100100;
assign F[59][26] = 9'b100100100;
assign F[59][27] = 9'b100100100;
assign F[59][28] = 9'b100100100;
assign F[59][29] = 9'b100100100;
assign F[60][0] = 9'b100100100;
assign F[60][1] = 9'b100100100;
assign F[60][2] = 9'b100100100;
assign F[60][3] = 9'b100100100;
assign F[60][4] = 9'b100100100;
assign F[60][5] = 9'b101001001;
assign F[60][6] = 9'b110111110;
assign F[60][7] = 9'b110111110;
assign F[60][8] = 9'b110111110;
assign F[60][9] = 9'b110111110;
assign F[60][10] = 9'b110111110;
assign F[60][11] = 9'b110111110;
assign F[60][12] = 9'b110111110;
assign F[60][13] = 9'b110111110;
assign F[60][14] = 9'b110111110;
assign F[60][15] = 9'b110111110;
assign F[60][16] = 9'b110111110;
assign F[60][17] = 9'b110111110;
assign F[60][18] = 9'b110111110;
assign F[60][19] = 9'b110111110;
assign F[60][20] = 9'b110111110;
assign F[60][21] = 9'b110111110;
assign F[60][22] = 9'b110111110;
assign F[60][23] = 9'b110111110;
assign F[60][24] = 9'b100100100;
assign F[60][25] = 9'b100100100;
assign F[60][26] = 9'b100100100;
assign F[60][27] = 9'b100100100;
assign F[60][28] = 9'b100100100;
assign F[60][29] = 9'b100100100;
assign F[61][0] = 9'b100100100;
assign F[61][1] = 9'b100100100;
assign F[61][2] = 9'b100100100;
assign F[61][3] = 9'b100100100;
assign F[61][4] = 9'b100100100;
assign F[61][5] = 9'b100100100;
assign F[61][6] = 9'b101001001;
assign F[61][7] = 9'b101001001;
assign F[61][8] = 9'b101101101;
assign F[61][9] = 9'b101101101;
assign F[61][10] = 9'b101101101;
assign F[61][11] = 9'b101101101;
assign F[61][12] = 9'b101101101;
assign F[61][13] = 9'b101101001;
assign F[61][14] = 9'b101101101;
assign F[61][15] = 9'b101101101;
assign F[61][16] = 9'b101101001;
assign F[61][17] = 9'b101101101;
assign F[61][18] = 9'b101101101;
assign F[61][19] = 9'b101101101;
assign F[61][20] = 9'b101101101;
assign F[61][21] = 9'b101101101;
assign F[61][22] = 9'b101001001;
assign F[61][23] = 9'b101001001;
assign F[61][24] = 9'b100100100;
assign F[61][25] = 9'b100100100;
assign F[61][26] = 9'b100100100;
assign F[61][27] = 9'b100100100;
assign F[61][28] = 9'b100100100;
assign F[61][29] = 9'b100100100;
assign F[62][0] = 9'b100100100;
assign F[62][1] = 9'b100100100;
assign F[62][2] = 9'b100100100;
assign F[62][3] = 9'b100100100;
assign F[62][4] = 9'b100100100;
assign F[62][5] = 9'b100100100;
assign F[62][6] = 9'b100000000;
assign F[62][7] = 9'b100000000;
assign F[62][8] = 9'b100100100;
assign F[62][9] = 9'b100100100;
assign F[62][10] = 9'b100100100;
assign F[62][11] = 9'b100100100;
assign F[62][12] = 9'b100100100;
assign F[62][13] = 9'b100000000;
assign F[62][14] = 9'b100100100;
assign F[62][15] = 9'b100100100;
assign F[62][16] = 9'b100000000;
assign F[62][17] = 9'b100100100;
assign F[62][18] = 9'b100100100;
assign F[62][19] = 9'b100100100;
assign F[62][20] = 9'b100100100;
assign F[62][21] = 9'b100100100;
assign F[62][22] = 9'b100000000;
assign F[62][23] = 9'b100000000;
assign F[62][24] = 9'b100100100;
assign F[62][25] = 9'b100100100;
assign F[62][26] = 9'b100100100;
assign F[62][27] = 9'b100100100;
assign F[62][28] = 9'b100100100;
assign F[62][29] = 9'b100100100;
assign F[63][0] = 9'b100100100;
assign F[63][1] = 9'b100100100;
assign F[63][2] = 9'b100100100;
assign F[63][3] = 9'b100100100;
assign F[63][4] = 9'b100100100;
assign F[63][5] = 9'b100100100;
assign F[63][6] = 9'b100100100;
assign F[63][7] = 9'b100100100;
assign F[63][8] = 9'b100100100;
assign F[63][9] = 9'b100100100;
assign F[63][10] = 9'b100100100;
assign F[63][11] = 9'b100100100;
assign F[63][12] = 9'b100100100;
assign F[63][13] = 9'b100100100;
assign F[63][14] = 9'b100100100;
assign F[63][15] = 9'b100100100;
assign F[63][16] = 9'b100100100;
assign F[63][17] = 9'b100100100;
assign F[63][18] = 9'b100100100;
assign F[63][19] = 9'b100100100;
assign F[63][20] = 9'b100100100;
assign F[63][21] = 9'b100100100;
assign F[63][22] = 9'b100100100;
assign F[63][23] = 9'b100100100;
assign F[63][24] = 9'b100100100;
assign F[63][25] = 9'b100100100;
assign F[63][26] = 9'b100100100;
assign F[63][27] = 9'b100100100;
assign F[63][28] = 9'b100100100;
assign F[63][29] = 9'b100100100;
assign F[64][0] = 9'b100100100;
assign F[64][1] = 9'b100100100;
assign F[64][2] = 9'b100100100;
assign F[64][3] = 9'b100100100;
assign F[64][4] = 9'b100100100;
assign F[64][5] = 9'b100100100;
assign F[64][6] = 9'b100100100;
assign F[64][7] = 9'b100100100;
assign F[64][8] = 9'b100100100;
assign F[64][9] = 9'b100100100;
assign F[64][10] = 9'b100100100;
assign F[64][11] = 9'b100100100;
assign F[64][12] = 9'b100100100;
assign F[64][13] = 9'b100100100;
assign F[64][14] = 9'b100100100;
assign F[64][15] = 9'b100100100;
assign F[64][16] = 9'b100100100;
assign F[64][17] = 9'b100100100;
assign F[64][18] = 9'b100100100;
assign F[64][19] = 9'b100100100;
assign F[64][20] = 9'b100100100;
assign F[64][21] = 9'b100100100;
assign F[64][22] = 9'b100100100;
assign F[64][23] = 9'b100100100;
assign F[64][24] = 9'b100100100;
assign F[64][25] = 9'b100100100;
assign F[64][26] = 9'b100100100;
assign F[64][27] = 9'b100100100;
assign F[64][28] = 9'b100100100;
assign F[64][29] = 9'b100100100;
assign F[65][0] = 9'b100100100;
assign F[65][1] = 9'b100100100;
assign F[65][2] = 9'b100100100;
assign F[65][3] = 9'b100100100;
assign F[65][4] = 9'b100100100;
assign F[65][5] = 9'b100100100;
assign F[65][6] = 9'b100100100;
assign F[65][7] = 9'b100100100;
assign F[65][8] = 9'b100100100;
assign F[65][9] = 9'b100100100;
assign F[65][10] = 9'b100100100;
assign F[65][11] = 9'b100100100;
assign F[65][12] = 9'b100100100;
assign F[65][13] = 9'b100100100;
assign F[65][14] = 9'b100100100;
assign F[65][15] = 9'b100100100;
assign F[65][16] = 9'b100100100;
assign F[65][17] = 9'b100100100;
assign F[65][18] = 9'b100100100;
assign F[65][19] = 9'b100100100;
assign F[65][20] = 9'b100100100;
assign F[65][21] = 9'b100100100;
assign F[65][22] = 9'b100100100;
assign F[65][23] = 9'b100100100;
assign F[65][24] = 9'b100100100;
assign F[65][25] = 9'b100100100;
assign F[65][26] = 9'b100100100;
assign F[65][27] = 9'b100100100;
assign F[65][28] = 9'b100100100;
assign F[65][29] = 9'b100100100;
assign F[66][0] = 9'b100100100;
assign F[66][1] = 9'b100100100;
assign F[66][2] = 9'b100100100;
assign F[66][3] = 9'b100100100;
assign F[66][4] = 9'b100100100;
assign F[66][5] = 9'b100100100;
assign F[66][6] = 9'b100100100;
assign F[66][7] = 9'b100100100;
assign F[66][22] = 9'b100100100;
assign F[66][23] = 9'b100100100;
assign F[66][24] = 9'b100100100;
assign F[66][25] = 9'b100100100;
assign F[66][26] = 9'b100100100;
assign F[66][27] = 9'b100100100;
assign F[66][28] = 9'b100100100;
assign F[66][29] = 9'b100100100;
assign F[67][1] = 9'b100100100;
assign F[67][2] = 9'b100100100;
assign F[67][3] = 9'b100100100;
assign F[67][4] = 9'b100100100;
assign F[67][5] = 9'b100100100;
assign F[67][6] = 9'b100100100;
assign F[67][23] = 9'b100100100;
assign F[67][24] = 9'b100100100;
assign F[67][25] = 9'b100100100;
assign F[67][26] = 9'b100100100;
assign F[67][27] = 9'b100100100;
assign F[67][28] = 9'b100100100;
//Total de Lineas = 1243
endmodule



