`timescale 1ns / 1ps
module prueba_3 (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (micromatri[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= micromatri[vcount- posy][hcount- posx][7:5];
				green <= micromatri[vcount- posy][hcount- posx][4:2];
            blue 	<= micromatri[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 100;
parameter RESOLUCION_Y = 50;
wire [8:0] micromatri[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign micromatri[0][0] = 9'b111111111;
assign micromatri[0][1] = 9'b111111111;
assign micromatri[0][2] = 9'b111111111;
assign micromatri[0][3] = 9'b111111111;
assign micromatri[0][4] = 9'b111111111;
assign micromatri[0][5] = 9'b111111111;
assign micromatri[0][6] = 9'b111111111;
assign micromatri[0][7] = 9'b111111111;
assign micromatri[0][8] = 9'b111111111;
assign micromatri[0][9] = 9'b111111111;
assign micromatri[0][10] = 9'b111111111;
assign micromatri[0][11] = 9'b111111111;
assign micromatri[0][12] = 9'b111111111;
assign micromatri[0][13] = 9'b111111111;
assign micromatri[0][14] = 9'b111111111;
assign micromatri[0][15] = 9'b111111111;
assign micromatri[0][16] = 9'b111111111;
assign micromatri[0][17] = 9'b111111111;
assign micromatri[0][18] = 9'b111111111;
assign micromatri[0][19] = 9'b111111111;
assign micromatri[0][20] = 9'b111111111;
assign micromatri[0][21] = 9'b111111111;
assign micromatri[0][22] = 9'b111111111;
assign micromatri[0][23] = 9'b111111111;
assign micromatri[0][24] = 9'b111111111;
assign micromatri[0][25] = 9'b111111111;
assign micromatri[0][26] = 9'b111111111;
assign micromatri[0][27] = 9'b111111111;
assign micromatri[0][28] = 9'b111111111;
assign micromatri[0][29] = 9'b111111111;
assign micromatri[0][30] = 9'b111111111;
assign micromatri[0][31] = 9'b111111111;
assign micromatri[0][32] = 9'b111111111;
assign micromatri[0][33] = 9'b111111111;
assign micromatri[0][34] = 9'b111111111;
assign micromatri[0][35] = 9'b111111111;
assign micromatri[0][36] = 9'b111111111;
assign micromatri[0][37] = 9'b111111111;
assign micromatri[0][38] = 9'b111111111;
assign micromatri[0][39] = 9'b111111111;
assign micromatri[0][40] = 9'b111111111;
assign micromatri[0][41] = 9'b111111111;
assign micromatri[0][42] = 9'b111111111;
assign micromatri[0][43] = 9'b111111111;
assign micromatri[0][44] = 9'b111111111;
assign micromatri[0][45] = 9'b111111111;
assign micromatri[0][46] = 9'b111111111;
assign micromatri[0][47] = 9'b111111111;
assign micromatri[0][48] = 9'b111111111;
assign micromatri[0][49] = 9'b111111111;
assign micromatri[0][50] = 9'b111111111;
assign micromatri[0][51] = 9'b111111111;
assign micromatri[0][52] = 9'b111111111;
assign micromatri[0][53] = 9'b111111111;
assign micromatri[0][54] = 9'b111111111;
assign micromatri[0][55] = 9'b111111111;
assign micromatri[0][56] = 9'b111111111;
assign micromatri[0][57] = 9'b111111111;
assign micromatri[0][58] = 9'b111111111;
assign micromatri[0][59] = 9'b111111111;
assign micromatri[0][60] = 9'b111111111;
assign micromatri[0][61] = 9'b111111111;
assign micromatri[0][62] = 9'b111111111;
assign micromatri[0][63] = 9'b111111111;
assign micromatri[0][64] = 9'b111111111;
assign micromatri[0][65] = 9'b111111111;
assign micromatri[0][66] = 9'b111111111;
assign micromatri[0][67] = 9'b111111111;
assign micromatri[0][68] = 9'b111111111;
assign micromatri[0][69] = 9'b111111111;
assign micromatri[0][70] = 9'b111111111;
assign micromatri[0][71] = 9'b111111111;
assign micromatri[0][72] = 9'b111111111;
assign micromatri[0][73] = 9'b111111111;
assign micromatri[0][74] = 9'b111111111;
assign micromatri[0][75] = 9'b111111111;
assign micromatri[0][76] = 9'b111111111;
assign micromatri[0][77] = 9'b111111111;
assign micromatri[0][78] = 9'b111111111;
assign micromatri[0][79] = 9'b111111111;
assign micromatri[0][80] = 9'b111111111;
assign micromatri[0][81] = 9'b111111111;
assign micromatri[0][82] = 9'b111111111;
assign micromatri[0][83] = 9'b111111111;
assign micromatri[0][84] = 9'b111111111;
assign micromatri[0][85] = 9'b111111111;
assign micromatri[0][86] = 9'b111111111;
assign micromatri[0][87] = 9'b111111111;
assign micromatri[0][88] = 9'b111111111;
assign micromatri[0][89] = 9'b111111111;
assign micromatri[0][90] = 9'b111111111;
assign micromatri[0][91] = 9'b111111111;
assign micromatri[0][92] = 9'b111111111;
assign micromatri[0][93] = 9'b111111111;
assign micromatri[0][94] = 9'b111111111;
assign micromatri[0][95] = 9'b111111111;
assign micromatri[0][96] = 9'b111111111;
assign micromatri[0][97] = 9'b111111111;
assign micromatri[0][98] = 9'b111111111;
assign micromatri[0][99] = 9'b111111111;
assign micromatri[1][0] = 9'b111111111;
assign micromatri[1][1] = 9'b111111111;
assign micromatri[1][2] = 9'b111111111;
assign micromatri[1][3] = 9'b111111111;
assign micromatri[1][4] = 9'b111111111;
assign micromatri[1][5] = 9'b111111111;
assign micromatri[1][6] = 9'b111111111;
assign micromatri[1][7] = 9'b111111111;
assign micromatri[1][8] = 9'b111111111;
assign micromatri[1][9] = 9'b111111111;
assign micromatri[1][10] = 9'b111111111;
assign micromatri[1][11] = 9'b111111111;
assign micromatri[1][12] = 9'b111111111;
assign micromatri[1][13] = 9'b111111111;
assign micromatri[1][14] = 9'b111111111;
assign micromatri[1][15] = 9'b111111111;
assign micromatri[1][16] = 9'b111111111;
assign micromatri[1][17] = 9'b111111111;
assign micromatri[1][18] = 9'b111111111;
assign micromatri[1][19] = 9'b111111111;
assign micromatri[1][20] = 9'b111111111;
assign micromatri[1][21] = 9'b111111111;
assign micromatri[1][22] = 9'b111111111;
assign micromatri[1][23] = 9'b111111111;
assign micromatri[1][24] = 9'b111111111;
assign micromatri[1][25] = 9'b111111111;
assign micromatri[1][26] = 9'b111111111;
assign micromatri[1][27] = 9'b111111111;
assign micromatri[1][28] = 9'b111111111;
assign micromatri[1][29] = 9'b111111111;
assign micromatri[1][30] = 9'b111111111;
assign micromatri[1][31] = 9'b111111111;
assign micromatri[1][32] = 9'b111111111;
assign micromatri[1][33] = 9'b111111111;
assign micromatri[1][34] = 9'b111111111;
assign micromatri[1][35] = 9'b111111111;
assign micromatri[1][36] = 9'b111111111;
assign micromatri[1][37] = 9'b111111111;
assign micromatri[1][38] = 9'b111111111;
assign micromatri[1][39] = 9'b111111111;
assign micromatri[1][40] = 9'b111111111;
assign micromatri[1][41] = 9'b111111111;
assign micromatri[1][42] = 9'b111111111;
assign micromatri[1][43] = 9'b111111111;
assign micromatri[1][44] = 9'b111111111;
assign micromatri[1][45] = 9'b111111111;
assign micromatri[1][46] = 9'b111111111;
assign micromatri[1][47] = 9'b111111111;
assign micromatri[1][48] = 9'b111111111;
assign micromatri[1][49] = 9'b111111111;
assign micromatri[1][50] = 9'b111111111;
assign micromatri[1][51] = 9'b111111111;
assign micromatri[1][52] = 9'b111111111;
assign micromatri[1][53] = 9'b111111111;
assign micromatri[1][54] = 9'b111111111;
assign micromatri[1][55] = 9'b111111111;
assign micromatri[1][56] = 9'b111111111;
assign micromatri[1][57] = 9'b111111111;
assign micromatri[1][58] = 9'b111111111;
assign micromatri[1][59] = 9'b111111111;
assign micromatri[1][60] = 9'b111111111;
assign micromatri[1][61] = 9'b111111111;
assign micromatri[1][62] = 9'b111111111;
assign micromatri[1][63] = 9'b111111111;
assign micromatri[1][64] = 9'b111111111;
assign micromatri[1][65] = 9'b111111111;
assign micromatri[1][66] = 9'b111111111;
assign micromatri[1][67] = 9'b111111111;
assign micromatri[1][68] = 9'b111111111;
assign micromatri[1][69] = 9'b111111111;
assign micromatri[1][70] = 9'b111111111;
assign micromatri[1][71] = 9'b111111111;
assign micromatri[1][72] = 9'b111111111;
assign micromatri[1][73] = 9'b111111111;
assign micromatri[1][74] = 9'b111111111;
assign micromatri[1][75] = 9'b111111111;
assign micromatri[1][76] = 9'b111111111;
assign micromatri[1][77] = 9'b111111111;
assign micromatri[1][78] = 9'b111111111;
assign micromatri[1][79] = 9'b111111111;
assign micromatri[1][80] = 9'b111111111;
assign micromatri[1][81] = 9'b111111111;
assign micromatri[1][82] = 9'b111111111;
assign micromatri[1][83] = 9'b111111111;
assign micromatri[1][84] = 9'b111111111;
assign micromatri[1][85] = 9'b111111111;
assign micromatri[1][86] = 9'b111111111;
assign micromatri[1][87] = 9'b111111111;
assign micromatri[1][88] = 9'b111111111;
assign micromatri[1][89] = 9'b111111111;
assign micromatri[1][90] = 9'b111111111;
assign micromatri[1][91] = 9'b111111111;
assign micromatri[1][92] = 9'b111111111;
assign micromatri[1][93] = 9'b111111111;
assign micromatri[1][94] = 9'b111111111;
assign micromatri[1][95] = 9'b111111111;
assign micromatri[1][96] = 9'b111111111;
assign micromatri[1][97] = 9'b111111111;
assign micromatri[1][98] = 9'b111111111;
assign micromatri[1][99] = 9'b111111111;
assign micromatri[2][0] = 9'b111111111;
assign micromatri[2][1] = 9'b111111111;
assign micromatri[2][2] = 9'b111111111;
assign micromatri[2][3] = 9'b111111111;
assign micromatri[2][4] = 9'b111111111;
assign micromatri[2][5] = 9'b111111111;
assign micromatri[2][6] = 9'b111111111;
assign micromatri[2][7] = 9'b111111111;
assign micromatri[2][8] = 9'b111111111;
assign micromatri[2][9] = 9'b111111111;
assign micromatri[2][10] = 9'b111111111;
assign micromatri[2][11] = 9'b111111111;
assign micromatri[2][12] = 9'b111111111;
assign micromatri[2][13] = 9'b111111111;
assign micromatri[2][14] = 9'b111111111;
assign micromatri[2][15] = 9'b111111111;
assign micromatri[2][16] = 9'b111111111;
assign micromatri[2][17] = 9'b111111111;
assign micromatri[2][18] = 9'b111111111;
assign micromatri[2][19] = 9'b111111111;
assign micromatri[2][20] = 9'b111111111;
assign micromatri[2][21] = 9'b111111111;
assign micromatri[2][22] = 9'b111111111;
assign micromatri[2][23] = 9'b111111111;
assign micromatri[2][24] = 9'b111111111;
assign micromatri[2][25] = 9'b111111111;
assign micromatri[2][26] = 9'b111111111;
assign micromatri[2][27] = 9'b111111111;
assign micromatri[2][28] = 9'b111111111;
assign micromatri[2][29] = 9'b111111111;
assign micromatri[2][30] = 9'b111111111;
assign micromatri[2][31] = 9'b111111111;
assign micromatri[2][32] = 9'b111111111;
assign micromatri[2][33] = 9'b111111111;
assign micromatri[2][34] = 9'b111111111;
assign micromatri[2][35] = 9'b111111111;
assign micromatri[2][36] = 9'b111111111;
assign micromatri[2][37] = 9'b111111111;
assign micromatri[2][38] = 9'b111111111;
assign micromatri[2][39] = 9'b111111111;
assign micromatri[2][40] = 9'b111111111;
assign micromatri[2][41] = 9'b111111111;
assign micromatri[2][42] = 9'b111111111;
assign micromatri[2][43] = 9'b111111111;
assign micromatri[2][44] = 9'b111111111;
assign micromatri[2][45] = 9'b111111111;
assign micromatri[2][46] = 9'b111111111;
assign micromatri[2][47] = 9'b111111111;
assign micromatri[2][48] = 9'b111111111;
assign micromatri[2][49] = 9'b111111111;
assign micromatri[2][50] = 9'b111111111;
assign micromatri[2][51] = 9'b111111111;
assign micromatri[2][52] = 9'b111111111;
assign micromatri[2][53] = 9'b111111111;
assign micromatri[2][54] = 9'b111111111;
assign micromatri[2][55] = 9'b111111111;
assign micromatri[2][56] = 9'b111111111;
assign micromatri[2][57] = 9'b111111111;
assign micromatri[2][58] = 9'b111111111;
assign micromatri[2][59] = 9'b111111111;
assign micromatri[2][60] = 9'b111111111;
assign micromatri[2][61] = 9'b111111111;
assign micromatri[2][62] = 9'b111111111;
assign micromatri[2][63] = 9'b111111111;
assign micromatri[2][64] = 9'b111111111;
assign micromatri[2][65] = 9'b111111111;
assign micromatri[2][66] = 9'b111111111;
assign micromatri[2][67] = 9'b111111111;
assign micromatri[2][68] = 9'b111111111;
assign micromatri[2][69] = 9'b111111111;
assign micromatri[2][70] = 9'b111111111;
assign micromatri[2][71] = 9'b111111111;
assign micromatri[2][72] = 9'b111111111;
assign micromatri[2][73] = 9'b111111111;
assign micromatri[2][74] = 9'b111111111;
assign micromatri[2][75] = 9'b111111111;
assign micromatri[2][76] = 9'b111111111;
assign micromatri[2][77] = 9'b111111111;
assign micromatri[2][78] = 9'b111111111;
assign micromatri[2][79] = 9'b111111111;
assign micromatri[2][80] = 9'b111111111;
assign micromatri[2][81] = 9'b111111111;
assign micromatri[2][82] = 9'b111111111;
assign micromatri[2][83] = 9'b111111111;
assign micromatri[2][84] = 9'b111111111;
assign micromatri[2][85] = 9'b111111111;
assign micromatri[2][86] = 9'b111111111;
assign micromatri[2][87] = 9'b111111111;
assign micromatri[2][88] = 9'b111111111;
assign micromatri[2][89] = 9'b111111111;
assign micromatri[2][90] = 9'b111111111;
assign micromatri[2][91] = 9'b111111111;
assign micromatri[2][92] = 9'b111111111;
assign micromatri[2][93] = 9'b111111111;
assign micromatri[2][94] = 9'b111111111;
assign micromatri[2][95] = 9'b111111111;
assign micromatri[2][96] = 9'b111111111;
assign micromatri[2][97] = 9'b111111111;
assign micromatri[2][98] = 9'b111111111;
assign micromatri[2][99] = 9'b111111111;
assign micromatri[3][0] = 9'b111111111;
assign micromatri[3][1] = 9'b111111111;
assign micromatri[3][2] = 9'b111111111;
assign micromatri[3][3] = 9'b111111111;
assign micromatri[3][4] = 9'b111111111;
assign micromatri[3][5] = 9'b111111111;
assign micromatri[3][6] = 9'b111111111;
assign micromatri[3][7] = 9'b111111111;
assign micromatri[3][8] = 9'b111111111;
assign micromatri[3][9] = 9'b111111111;
assign micromatri[3][10] = 9'b111111111;
assign micromatri[3][11] = 9'b111111111;
assign micromatri[3][12] = 9'b111111111;
assign micromatri[3][13] = 9'b111111111;
assign micromatri[3][14] = 9'b111111111;
assign micromatri[3][15] = 9'b111111111;
assign micromatri[3][16] = 9'b111111111;
assign micromatri[3][17] = 9'b111111111;
assign micromatri[3][18] = 9'b111111111;
assign micromatri[3][19] = 9'b111111111;
assign micromatri[3][20] = 9'b111111111;
assign micromatri[3][21] = 9'b111111111;
assign micromatri[3][22] = 9'b111111111;
assign micromatri[3][23] = 9'b111111111;
assign micromatri[3][24] = 9'b111111111;
assign micromatri[3][25] = 9'b111111111;
assign micromatri[3][26] = 9'b111111111;
assign micromatri[3][27] = 9'b111111111;
assign micromatri[3][28] = 9'b111111111;
assign micromatri[3][29] = 9'b111111111;
assign micromatri[3][30] = 9'b111111111;
assign micromatri[3][31] = 9'b111111111;
assign micromatri[3][32] = 9'b111111111;
assign micromatri[3][33] = 9'b111111111;
assign micromatri[3][34] = 9'b111111111;
assign micromatri[3][35] = 9'b111111111;
assign micromatri[3][36] = 9'b111111111;
assign micromatri[3][37] = 9'b111111111;
assign micromatri[3][38] = 9'b111111111;
assign micromatri[3][39] = 9'b111111111;
assign micromatri[3][40] = 9'b111111111;
assign micromatri[3][41] = 9'b111111111;
assign micromatri[3][42] = 9'b111111111;
assign micromatri[3][43] = 9'b111111111;
assign micromatri[3][44] = 9'b111111111;
assign micromatri[3][45] = 9'b111111111;
assign micromatri[3][46] = 9'b111111111;
assign micromatri[3][47] = 9'b111111111;
assign micromatri[3][48] = 9'b111111111;
assign micromatri[3][49] = 9'b111111111;
assign micromatri[3][50] = 9'b111111111;
assign micromatri[3][51] = 9'b111111111;
assign micromatri[3][52] = 9'b111111111;
assign micromatri[3][53] = 9'b111111111;
assign micromatri[3][54] = 9'b111111111;
assign micromatri[3][55] = 9'b111111111;
assign micromatri[3][56] = 9'b111111111;
assign micromatri[3][57] = 9'b111111111;
assign micromatri[3][58] = 9'b111111111;
assign micromatri[3][59] = 9'b111111111;
assign micromatri[3][60] = 9'b111111111;
assign micromatri[3][61] = 9'b111111111;
assign micromatri[3][62] = 9'b111111111;
assign micromatri[3][63] = 9'b111111111;
assign micromatri[3][64] = 9'b111111111;
assign micromatri[3][65] = 9'b111111111;
assign micromatri[3][66] = 9'b111111111;
assign micromatri[3][67] = 9'b111111111;
assign micromatri[3][68] = 9'b111111111;
assign micromatri[3][69] = 9'b111111111;
assign micromatri[3][70] = 9'b111111111;
assign micromatri[3][71] = 9'b111111111;
assign micromatri[3][72] = 9'b111111111;
assign micromatri[3][73] = 9'b111111111;
assign micromatri[3][74] = 9'b111111111;
assign micromatri[3][75] = 9'b111111111;
assign micromatri[3][76] = 9'b111111111;
assign micromatri[3][77] = 9'b111111111;
assign micromatri[3][78] = 9'b111111111;
assign micromatri[3][79] = 9'b111111111;
assign micromatri[3][80] = 9'b111111111;
assign micromatri[3][81] = 9'b111111111;
assign micromatri[3][82] = 9'b111111111;
assign micromatri[3][83] = 9'b111111111;
assign micromatri[3][84] = 9'b111111111;
assign micromatri[3][85] = 9'b111111111;
assign micromatri[3][86] = 9'b111111111;
assign micromatri[3][87] = 9'b111111111;
assign micromatri[3][88] = 9'b111111111;
assign micromatri[3][89] = 9'b111111111;
assign micromatri[3][90] = 9'b111111111;
assign micromatri[3][91] = 9'b111111111;
assign micromatri[3][92] = 9'b111111111;
assign micromatri[3][93] = 9'b111111111;
assign micromatri[3][94] = 9'b111111111;
assign micromatri[3][95] = 9'b111111111;
assign micromatri[3][96] = 9'b111111111;
assign micromatri[3][97] = 9'b111111111;
assign micromatri[3][98] = 9'b111111111;
assign micromatri[3][99] = 9'b111111111;
assign micromatri[4][0] = 9'b111111111;
assign micromatri[4][1] = 9'b111111111;
assign micromatri[4][2] = 9'b111111111;
assign micromatri[4][3] = 9'b111111111;
assign micromatri[4][4] = 9'b111111111;
assign micromatri[4][5] = 9'b111111111;
assign micromatri[4][6] = 9'b111111111;
assign micromatri[4][7] = 9'b111111111;
assign micromatri[4][8] = 9'b111111111;
assign micromatri[4][9] = 9'b111111111;
assign micromatri[4][10] = 9'b111111111;
assign micromatri[4][11] = 9'b111111111;
assign micromatri[4][12] = 9'b111111111;
assign micromatri[4][13] = 9'b111111111;
assign micromatri[4][14] = 9'b111111111;
assign micromatri[4][15] = 9'b111111111;
assign micromatri[4][16] = 9'b111111111;
assign micromatri[4][17] = 9'b111111111;
assign micromatri[4][18] = 9'b111111111;
assign micromatri[4][19] = 9'b111111111;
assign micromatri[4][20] = 9'b111111111;
assign micromatri[4][21] = 9'b111111111;
assign micromatri[4][22] = 9'b111111111;
assign micromatri[4][23] = 9'b111111111;
assign micromatri[4][24] = 9'b111111111;
assign micromatri[4][25] = 9'b111111111;
assign micromatri[4][26] = 9'b111111111;
assign micromatri[4][27] = 9'b111111111;
assign micromatri[4][28] = 9'b111111111;
assign micromatri[4][29] = 9'b111111111;
assign micromatri[4][30] = 9'b111111111;
assign micromatri[4][31] = 9'b111111111;
assign micromatri[4][32] = 9'b111111111;
assign micromatri[4][33] = 9'b111111111;
assign micromatri[4][34] = 9'b111111111;
assign micromatri[4][35] = 9'b111111111;
assign micromatri[4][36] = 9'b111111111;
assign micromatri[4][37] = 9'b111111111;
assign micromatri[4][38] = 9'b111111111;
assign micromatri[4][39] = 9'b111111111;
assign micromatri[4][40] = 9'b111111111;
assign micromatri[4][41] = 9'b111111111;
assign micromatri[4][42] = 9'b111111111;
assign micromatri[4][43] = 9'b111111111;
assign micromatri[4][44] = 9'b111111111;
assign micromatri[4][45] = 9'b111111111;
assign micromatri[4][46] = 9'b111111111;
assign micromatri[4][47] = 9'b111111111;
assign micromatri[4][48] = 9'b111111111;
assign micromatri[4][49] = 9'b111111111;
assign micromatri[4][50] = 9'b111111111;
assign micromatri[4][51] = 9'b111111111;
assign micromatri[4][52] = 9'b111111111;
assign micromatri[4][53] = 9'b111111111;
assign micromatri[4][54] = 9'b111111111;
assign micromatri[4][55] = 9'b111111111;
assign micromatri[4][56] = 9'b111111111;
assign micromatri[4][57] = 9'b111111111;
assign micromatri[4][58] = 9'b111111111;
assign micromatri[4][59] = 9'b111111111;
assign micromatri[4][60] = 9'b111111111;
assign micromatri[4][61] = 9'b111111111;
assign micromatri[4][62] = 9'b111111111;
assign micromatri[4][63] = 9'b111111111;
assign micromatri[4][64] = 9'b111111111;
assign micromatri[4][65] = 9'b111111111;
assign micromatri[4][66] = 9'b111111111;
assign micromatri[4][67] = 9'b111111111;
assign micromatri[4][68] = 9'b111111111;
assign micromatri[4][69] = 9'b111111111;
assign micromatri[4][70] = 9'b111111111;
assign micromatri[4][71] = 9'b111111111;
assign micromatri[4][72] = 9'b111111111;
assign micromatri[4][73] = 9'b111111111;
assign micromatri[4][74] = 9'b111111111;
assign micromatri[4][75] = 9'b111111111;
assign micromatri[4][76] = 9'b111111111;
assign micromatri[4][77] = 9'b111111111;
assign micromatri[4][78] = 9'b111111111;
assign micromatri[4][79] = 9'b111111111;
assign micromatri[4][80] = 9'b111111111;
assign micromatri[4][81] = 9'b111111111;
assign micromatri[4][82] = 9'b111111111;
assign micromatri[4][83] = 9'b111111111;
assign micromatri[4][84] = 9'b111111111;
assign micromatri[4][85] = 9'b111111111;
assign micromatri[4][86] = 9'b111111111;
assign micromatri[4][87] = 9'b111111111;
assign micromatri[4][88] = 9'b111111111;
assign micromatri[4][89] = 9'b111111111;
assign micromatri[4][90] = 9'b111111111;
assign micromatri[4][91] = 9'b111111111;
assign micromatri[4][92] = 9'b111111111;
assign micromatri[4][93] = 9'b111111111;
assign micromatri[4][94] = 9'b111111111;
assign micromatri[4][95] = 9'b111111111;
assign micromatri[4][96] = 9'b111111111;
assign micromatri[4][97] = 9'b111111111;
assign micromatri[4][98] = 9'b111111111;
assign micromatri[4][99] = 9'b111111111;
assign micromatri[5][0] = 9'b111111111;
assign micromatri[5][1] = 9'b111111111;
assign micromatri[5][2] = 9'b111111111;
assign micromatri[5][3] = 9'b111111111;
assign micromatri[5][4] = 9'b111111111;
assign micromatri[5][5] = 9'b111111111;
assign micromatri[5][6] = 9'b111111111;
assign micromatri[5][7] = 9'b111111111;
assign micromatri[5][8] = 9'b111111111;
assign micromatri[5][9] = 9'b111111111;
assign micromatri[5][10] = 9'b111111111;
assign micromatri[5][11] = 9'b111111111;
assign micromatri[5][12] = 9'b111111111;
assign micromatri[5][13] = 9'b111111111;
assign micromatri[5][14] = 9'b111111111;
assign micromatri[5][15] = 9'b111111111;
assign micromatri[5][16] = 9'b111111111;
assign micromatri[5][17] = 9'b111111111;
assign micromatri[5][18] = 9'b111111111;
assign micromatri[5][19] = 9'b111111111;
assign micromatri[5][20] = 9'b111111111;
assign micromatri[5][21] = 9'b111111111;
assign micromatri[5][22] = 9'b111111111;
assign micromatri[5][23] = 9'b111111111;
assign micromatri[5][24] = 9'b111111111;
assign micromatri[5][25] = 9'b111111111;
assign micromatri[5][26] = 9'b111111111;
assign micromatri[5][27] = 9'b111111111;
assign micromatri[5][28] = 9'b111111111;
assign micromatri[5][29] = 9'b111111111;
assign micromatri[5][30] = 9'b111111111;
assign micromatri[5][31] = 9'b111111111;
assign micromatri[5][32] = 9'b111111111;
assign micromatri[5][33] = 9'b111111111;
assign micromatri[5][34] = 9'b111111111;
assign micromatri[5][35] = 9'b111111111;
assign micromatri[5][36] = 9'b111111111;
assign micromatri[5][37] = 9'b111111111;
assign micromatri[5][38] = 9'b111111111;
assign micromatri[5][39] = 9'b111111111;
assign micromatri[5][40] = 9'b111111111;
assign micromatri[5][41] = 9'b111111111;
assign micromatri[5][42] = 9'b111111111;
assign micromatri[5][43] = 9'b111111111;
assign micromatri[5][44] = 9'b111111111;
assign micromatri[5][45] = 9'b111111111;
assign micromatri[5][46] = 9'b111111111;
assign micromatri[5][47] = 9'b111111111;
assign micromatri[5][48] = 9'b111111111;
assign micromatri[5][49] = 9'b111111111;
assign micromatri[5][50] = 9'b111111111;
assign micromatri[5][51] = 9'b111111111;
assign micromatri[5][52] = 9'b111111111;
assign micromatri[5][53] = 9'b111111111;
assign micromatri[5][54] = 9'b111111111;
assign micromatri[5][55] = 9'b111111111;
assign micromatri[5][56] = 9'b111111111;
assign micromatri[5][57] = 9'b111111111;
assign micromatri[5][58] = 9'b111111111;
assign micromatri[5][59] = 9'b111111111;
assign micromatri[5][60] = 9'b111111111;
assign micromatri[5][61] = 9'b111111111;
assign micromatri[5][62] = 9'b111111111;
assign micromatri[5][63] = 9'b111111111;
assign micromatri[5][64] = 9'b111111111;
assign micromatri[5][65] = 9'b111111111;
assign micromatri[5][66] = 9'b111111111;
assign micromatri[5][67] = 9'b111111111;
assign micromatri[5][68] = 9'b111111111;
assign micromatri[5][69] = 9'b111111111;
assign micromatri[5][70] = 9'b111111111;
assign micromatri[5][71] = 9'b111111111;
assign micromatri[5][72] = 9'b111111111;
assign micromatri[5][73] = 9'b111111111;
assign micromatri[5][74] = 9'b111111111;
assign micromatri[5][75] = 9'b111111111;
assign micromatri[5][76] = 9'b111111111;
assign micromatri[5][77] = 9'b111111111;
assign micromatri[5][78] = 9'b111111111;
assign micromatri[5][79] = 9'b111111111;
assign micromatri[5][80] = 9'b111111111;
assign micromatri[5][81] = 9'b111111111;
assign micromatri[5][82] = 9'b111111111;
assign micromatri[5][83] = 9'b111111111;
assign micromatri[5][84] = 9'b111111111;
assign micromatri[5][85] = 9'b111111111;
assign micromatri[5][86] = 9'b111111111;
assign micromatri[5][87] = 9'b111111111;
assign micromatri[5][88] = 9'b111111111;
assign micromatri[5][89] = 9'b111111111;
assign micromatri[5][90] = 9'b111111111;
assign micromatri[5][91] = 9'b111111111;
assign micromatri[5][92] = 9'b111111111;
assign micromatri[5][93] = 9'b111111111;
assign micromatri[5][94] = 9'b111111111;
assign micromatri[5][95] = 9'b111111111;
assign micromatri[5][96] = 9'b111111111;
assign micromatri[5][97] = 9'b111111111;
assign micromatri[5][98] = 9'b111111111;
assign micromatri[5][99] = 9'b111111111;
assign micromatri[6][0] = 9'b111111111;
assign micromatri[6][1] = 9'b111111111;
assign micromatri[6][2] = 9'b111111111;
assign micromatri[6][3] = 9'b111111111;
assign micromatri[6][4] = 9'b111111111;
assign micromatri[6][5] = 9'b111111111;
assign micromatri[6][6] = 9'b111111111;
assign micromatri[6][7] = 9'b111111111;
assign micromatri[6][8] = 9'b111111111;
assign micromatri[6][9] = 9'b111111111;
assign micromatri[6][10] = 9'b111111111;
assign micromatri[6][11] = 9'b111111111;
assign micromatri[6][12] = 9'b111111111;
assign micromatri[6][13] = 9'b111111111;
assign micromatri[6][14] = 9'b111111111;
assign micromatri[6][15] = 9'b111111111;
assign micromatri[6][16] = 9'b111111111;
assign micromatri[6][17] = 9'b111111111;
assign micromatri[6][18] = 9'b111111111;
assign micromatri[6][19] = 9'b111111111;
assign micromatri[6][20] = 9'b111111111;
assign micromatri[6][21] = 9'b111111111;
assign micromatri[6][22] = 9'b111111111;
assign micromatri[6][23] = 9'b111111111;
assign micromatri[6][24] = 9'b111111111;
assign micromatri[6][25] = 9'b111111111;
assign micromatri[6][26] = 9'b111111111;
assign micromatri[6][27] = 9'b111111111;
assign micromatri[6][28] = 9'b111111111;
assign micromatri[6][29] = 9'b111111111;
assign micromatri[6][30] = 9'b111111111;
assign micromatri[6][31] = 9'b111111111;
assign micromatri[6][32] = 9'b111111111;
assign micromatri[6][33] = 9'b111111111;
assign micromatri[6][34] = 9'b111111111;
assign micromatri[6][35] = 9'b111111111;
assign micromatri[6][36] = 9'b111111111;
assign micromatri[6][37] = 9'b111111111;
assign micromatri[6][38] = 9'b111111111;
assign micromatri[6][39] = 9'b111111111;
assign micromatri[6][40] = 9'b111111111;
assign micromatri[6][41] = 9'b111111111;
assign micromatri[6][42] = 9'b111111111;
assign micromatri[6][43] = 9'b111111111;
assign micromatri[6][44] = 9'b111111111;
assign micromatri[6][45] = 9'b111111111;
assign micromatri[6][46] = 9'b111111111;
assign micromatri[6][47] = 9'b111111111;
assign micromatri[6][48] = 9'b111111111;
assign micromatri[6][49] = 9'b111111111;
assign micromatri[6][50] = 9'b111111111;
assign micromatri[6][51] = 9'b111111111;
assign micromatri[6][52] = 9'b111111111;
assign micromatri[6][53] = 9'b111111111;
assign micromatri[6][54] = 9'b111111111;
assign micromatri[6][55] = 9'b111111111;
assign micromatri[6][56] = 9'b111111111;
assign micromatri[6][57] = 9'b111111111;
assign micromatri[6][58] = 9'b111111111;
assign micromatri[6][59] = 9'b111111111;
assign micromatri[6][60] = 9'b111111111;
assign micromatri[6][61] = 9'b111111111;
assign micromatri[6][62] = 9'b111111111;
assign micromatri[6][63] = 9'b111111111;
assign micromatri[6][64] = 9'b111111111;
assign micromatri[6][65] = 9'b111111111;
assign micromatri[6][66] = 9'b111111111;
assign micromatri[6][67] = 9'b111111111;
assign micromatri[6][68] = 9'b111111111;
assign micromatri[6][69] = 9'b111111111;
assign micromatri[6][70] = 9'b111111111;
assign micromatri[6][71] = 9'b111111111;
assign micromatri[6][72] = 9'b111111111;
assign micromatri[6][73] = 9'b111111111;
assign micromatri[6][74] = 9'b111111111;
assign micromatri[6][75] = 9'b111111111;
assign micromatri[6][76] = 9'b111111111;
assign micromatri[6][77] = 9'b111111111;
assign micromatri[6][78] = 9'b111111111;
assign micromatri[6][79] = 9'b111111111;
assign micromatri[6][80] = 9'b111111111;
assign micromatri[6][81] = 9'b111111111;
assign micromatri[6][82] = 9'b111111111;
assign micromatri[6][83] = 9'b111111111;
assign micromatri[6][84] = 9'b111111111;
assign micromatri[6][85] = 9'b111111111;
assign micromatri[6][86] = 9'b111111111;
assign micromatri[6][87] = 9'b111111111;
assign micromatri[6][88] = 9'b111111111;
assign micromatri[6][89] = 9'b111111111;
assign micromatri[6][90] = 9'b111111111;
assign micromatri[6][91] = 9'b111111111;
assign micromatri[6][92] = 9'b111111111;
assign micromatri[6][93] = 9'b111111111;
assign micromatri[6][94] = 9'b111111111;
assign micromatri[6][95] = 9'b111111111;
assign micromatri[6][96] = 9'b111111111;
assign micromatri[6][97] = 9'b111111111;
assign micromatri[6][98] = 9'b111111111;
assign micromatri[6][99] = 9'b111111111;
assign micromatri[7][0] = 9'b111111111;
assign micromatri[7][1] = 9'b111111111;
assign micromatri[7][2] = 9'b111111111;
assign micromatri[7][3] = 9'b111111111;
assign micromatri[7][4] = 9'b111111111;
assign micromatri[7][5] = 9'b111111111;
assign micromatri[7][6] = 9'b111111111;
assign micromatri[7][7] = 9'b111111111;
assign micromatri[7][8] = 9'b111111111;
assign micromatri[7][9] = 9'b111111111;
assign micromatri[7][10] = 9'b111111111;
assign micromatri[7][11] = 9'b111111111;
assign micromatri[7][12] = 9'b111111111;
assign micromatri[7][13] = 9'b111111111;
assign micromatri[7][14] = 9'b111111111;
assign micromatri[7][15] = 9'b111111111;
assign micromatri[7][16] = 9'b111111111;
assign micromatri[7][17] = 9'b111111111;
assign micromatri[7][18] = 9'b111111111;
assign micromatri[7][19] = 9'b111111111;
assign micromatri[7][20] = 9'b111111111;
assign micromatri[7][21] = 9'b111111111;
assign micromatri[7][22] = 9'b111111111;
assign micromatri[7][23] = 9'b111111111;
assign micromatri[7][24] = 9'b111111111;
assign micromatri[7][25] = 9'b111111111;
assign micromatri[7][26] = 9'b111111111;
assign micromatri[7][27] = 9'b111111111;
assign micromatri[7][28] = 9'b111111111;
assign micromatri[7][29] = 9'b111111111;
assign micromatri[7][30] = 9'b111111111;
assign micromatri[7][31] = 9'b111111111;
assign micromatri[7][32] = 9'b111111111;
assign micromatri[7][33] = 9'b111111111;
assign micromatri[7][34] = 9'b111111111;
assign micromatri[7][35] = 9'b111111111;
assign micromatri[7][36] = 9'b111111111;
assign micromatri[7][37] = 9'b111111111;
assign micromatri[7][38] = 9'b111111111;
assign micromatri[7][39] = 9'b111111111;
assign micromatri[7][40] = 9'b111111111;
assign micromatri[7][41] = 9'b111111111;
assign micromatri[7][42] = 9'b111111111;
assign micromatri[7][43] = 9'b111111111;
assign micromatri[7][44] = 9'b111111111;
assign micromatri[7][45] = 9'b111111111;
assign micromatri[7][46] = 9'b111111111;
assign micromatri[7][47] = 9'b111111111;
assign micromatri[7][48] = 9'b111111111;
assign micromatri[7][49] = 9'b111111111;
assign micromatri[7][50] = 9'b111111111;
assign micromatri[7][51] = 9'b111111111;
assign micromatri[7][52] = 9'b111111111;
assign micromatri[7][53] = 9'b111111111;
assign micromatri[7][54] = 9'b111111111;
assign micromatri[7][55] = 9'b111111111;
assign micromatri[7][56] = 9'b111111111;
assign micromatri[7][57] = 9'b111111111;
assign micromatri[7][58] = 9'b111111111;
assign micromatri[7][59] = 9'b111111111;
assign micromatri[7][60] = 9'b111111111;
assign micromatri[7][61] = 9'b111111111;
assign micromatri[7][62] = 9'b111111111;
assign micromatri[7][63] = 9'b111111111;
assign micromatri[7][64] = 9'b111111111;
assign micromatri[7][65] = 9'b111111111;
assign micromatri[7][66] = 9'b111111111;
assign micromatri[7][67] = 9'b111111111;
assign micromatri[7][68] = 9'b111111111;
assign micromatri[7][69] = 9'b111111111;
assign micromatri[7][70] = 9'b111111111;
assign micromatri[7][71] = 9'b111111111;
assign micromatri[7][72] = 9'b111111111;
assign micromatri[7][73] = 9'b111111111;
assign micromatri[7][74] = 9'b111111111;
assign micromatri[7][75] = 9'b111111111;
assign micromatri[7][76] = 9'b111111111;
assign micromatri[7][77] = 9'b111111111;
assign micromatri[7][78] = 9'b111111111;
assign micromatri[7][79] = 9'b111111111;
assign micromatri[7][80] = 9'b111111111;
assign micromatri[7][81] = 9'b111111111;
assign micromatri[7][82] = 9'b111111111;
assign micromatri[7][83] = 9'b111111111;
assign micromatri[7][84] = 9'b111111111;
assign micromatri[7][85] = 9'b111111111;
assign micromatri[7][86] = 9'b111111111;
assign micromatri[7][87] = 9'b111111111;
assign micromatri[7][88] = 9'b111111111;
assign micromatri[7][89] = 9'b111111111;
assign micromatri[7][90] = 9'b111111111;
assign micromatri[7][91] = 9'b111111111;
assign micromatri[7][92] = 9'b111111111;
assign micromatri[7][93] = 9'b111111111;
assign micromatri[7][94] = 9'b111111111;
assign micromatri[7][95] = 9'b111111111;
assign micromatri[7][96] = 9'b111111111;
assign micromatri[7][97] = 9'b111111111;
assign micromatri[7][98] = 9'b111111111;
assign micromatri[7][99] = 9'b111111111;
assign micromatri[8][0] = 9'b111111111;
assign micromatri[8][1] = 9'b111111111;
assign micromatri[8][2] = 9'b111111111;
assign micromatri[8][3] = 9'b111111111;
assign micromatri[8][4] = 9'b111111111;
assign micromatri[8][5] = 9'b111111111;
assign micromatri[8][6] = 9'b111111111;
assign micromatri[8][7] = 9'b111111111;
assign micromatri[8][8] = 9'b111111111;
assign micromatri[8][9] = 9'b111111111;
assign micromatri[8][10] = 9'b111111111;
assign micromatri[8][11] = 9'b111111111;
assign micromatri[8][12] = 9'b111111111;
assign micromatri[8][13] = 9'b111111111;
assign micromatri[8][14] = 9'b111111111;
assign micromatri[8][15] = 9'b111111111;
assign micromatri[8][16] = 9'b111111111;
assign micromatri[8][17] = 9'b111111111;
assign micromatri[8][18] = 9'b111111111;
assign micromatri[8][19] = 9'b111111111;
assign micromatri[8][20] = 9'b111111111;
assign micromatri[8][21] = 9'b111111111;
assign micromatri[8][22] = 9'b111111111;
assign micromatri[8][23] = 9'b111111111;
assign micromatri[8][24] = 9'b111111111;
assign micromatri[8][25] = 9'b111111111;
assign micromatri[8][26] = 9'b111111111;
assign micromatri[8][27] = 9'b111111111;
assign micromatri[8][28] = 9'b111111111;
assign micromatri[8][29] = 9'b111111111;
assign micromatri[8][30] = 9'b111111111;
assign micromatri[8][31] = 9'b111111111;
assign micromatri[8][32] = 9'b111111111;
assign micromatri[8][33] = 9'b111111111;
assign micromatri[8][34] = 9'b111111111;
assign micromatri[8][35] = 9'b111111111;
assign micromatri[8][36] = 9'b111111111;
assign micromatri[8][37] = 9'b111111111;
assign micromatri[8][38] = 9'b111111111;
assign micromatri[8][39] = 9'b111111111;
assign micromatri[8][40] = 9'b111111111;
assign micromatri[8][41] = 9'b111111111;
assign micromatri[8][42] = 9'b111111111;
assign micromatri[8][43] = 9'b111111111;
assign micromatri[8][44] = 9'b111111111;
assign micromatri[8][45] = 9'b111111111;
assign micromatri[8][46] = 9'b111111111;
assign micromatri[8][47] = 9'b111111111;
assign micromatri[8][48] = 9'b111111111;
assign micromatri[8][49] = 9'b111111111;
assign micromatri[8][50] = 9'b111111111;
assign micromatri[8][51] = 9'b111111111;
assign micromatri[8][52] = 9'b111111111;
assign micromatri[8][53] = 9'b111111111;
assign micromatri[8][54] = 9'b111111111;
assign micromatri[8][55] = 9'b111111111;
assign micromatri[8][56] = 9'b111111111;
assign micromatri[8][57] = 9'b111111111;
assign micromatri[8][58] = 9'b111111111;
assign micromatri[8][59] = 9'b111111111;
assign micromatri[8][60] = 9'b111111111;
assign micromatri[8][61] = 9'b111111111;
assign micromatri[8][62] = 9'b111111111;
assign micromatri[8][63] = 9'b111111111;
assign micromatri[8][64] = 9'b111111111;
assign micromatri[8][65] = 9'b111111111;
assign micromatri[8][66] = 9'b111111111;
assign micromatri[8][67] = 9'b111111111;
assign micromatri[8][68] = 9'b111111111;
assign micromatri[8][69] = 9'b111111111;
assign micromatri[8][70] = 9'b111111111;
assign micromatri[8][71] = 9'b111111111;
assign micromatri[8][72] = 9'b111111111;
assign micromatri[8][73] = 9'b111111111;
assign micromatri[8][74] = 9'b111111111;
assign micromatri[8][75] = 9'b111111111;
assign micromatri[8][76] = 9'b111111111;
assign micromatri[8][77] = 9'b111111111;
assign micromatri[8][78] = 9'b111111111;
assign micromatri[8][79] = 9'b111111111;
assign micromatri[8][80] = 9'b111111111;
assign micromatri[8][81] = 9'b111111111;
assign micromatri[8][82] = 9'b111111111;
assign micromatri[8][83] = 9'b111111111;
assign micromatri[8][84] = 9'b111111111;
assign micromatri[8][85] = 9'b111111111;
assign micromatri[8][86] = 9'b111111111;
assign micromatri[8][87] = 9'b111111111;
assign micromatri[8][88] = 9'b111111111;
assign micromatri[8][89] = 9'b111111111;
assign micromatri[8][90] = 9'b111111111;
assign micromatri[8][91] = 9'b111111111;
assign micromatri[8][92] = 9'b111111111;
assign micromatri[8][93] = 9'b111111111;
assign micromatri[8][94] = 9'b111111111;
assign micromatri[8][95] = 9'b111111111;
assign micromatri[8][96] = 9'b111111111;
assign micromatri[8][97] = 9'b111111111;
assign micromatri[8][98] = 9'b111111111;
assign micromatri[8][99] = 9'b111111111;
assign micromatri[9][0] = 9'b111111111;
assign micromatri[9][1] = 9'b111111111;
assign micromatri[9][2] = 9'b111111111;
assign micromatri[9][3] = 9'b111111111;
assign micromatri[9][4] = 9'b111111111;
assign micromatri[9][5] = 9'b111111111;
assign micromatri[9][6] = 9'b111111111;
assign micromatri[9][7] = 9'b111111111;
assign micromatri[9][8] = 9'b111111111;
assign micromatri[9][9] = 9'b111111111;
assign micromatri[9][10] = 9'b111111111;
assign micromatri[9][11] = 9'b111111111;
assign micromatri[9][12] = 9'b111111111;
assign micromatri[9][13] = 9'b111111111;
assign micromatri[9][14] = 9'b111111111;
assign micromatri[9][15] = 9'b111111111;
assign micromatri[9][16] = 9'b111111111;
assign micromatri[9][17] = 9'b111111111;
assign micromatri[9][18] = 9'b111111111;
assign micromatri[9][19] = 9'b111111111;
assign micromatri[9][20] = 9'b111111111;
assign micromatri[9][21] = 9'b111111111;
assign micromatri[9][22] = 9'b111111111;
assign micromatri[9][23] = 9'b111111111;
assign micromatri[9][24] = 9'b111111111;
assign micromatri[9][25] = 9'b111111111;
assign micromatri[9][26] = 9'b111111111;
assign micromatri[9][27] = 9'b111111111;
assign micromatri[9][28] = 9'b111111111;
assign micromatri[9][29] = 9'b111111111;
assign micromatri[9][30] = 9'b111111111;
assign micromatri[9][31] = 9'b111111111;
assign micromatri[9][32] = 9'b111111111;
assign micromatri[9][33] = 9'b111111111;
assign micromatri[9][34] = 9'b111111111;
assign micromatri[9][35] = 9'b111111111;
assign micromatri[9][36] = 9'b111111111;
assign micromatri[9][37] = 9'b111111111;
assign micromatri[9][38] = 9'b111111111;
assign micromatri[9][39] = 9'b111111111;
assign micromatri[9][40] = 9'b111111111;
assign micromatri[9][41] = 9'b111111111;
assign micromatri[9][42] = 9'b111111111;
assign micromatri[9][43] = 9'b111111111;
assign micromatri[9][44] = 9'b111111111;
assign micromatri[9][45] = 9'b111111111;
assign micromatri[9][46] = 9'b111111111;
assign micromatri[9][47] = 9'b111111111;
assign micromatri[9][48] = 9'b111111111;
assign micromatri[9][49] = 9'b111111111;
assign micromatri[9][50] = 9'b111111111;
assign micromatri[9][51] = 9'b111111111;
assign micromatri[9][52] = 9'b111111111;
assign micromatri[9][53] = 9'b111111111;
assign micromatri[9][54] = 9'b111111111;
assign micromatri[9][55] = 9'b111111111;
assign micromatri[9][56] = 9'b111111111;
assign micromatri[9][57] = 9'b111111111;
assign micromatri[9][58] = 9'b111111111;
assign micromatri[9][59] = 9'b111111111;
assign micromatri[9][60] = 9'b111111111;
assign micromatri[9][61] = 9'b111111111;
assign micromatri[9][62] = 9'b111111111;
assign micromatri[9][63] = 9'b111111111;
assign micromatri[9][64] = 9'b111111111;
assign micromatri[9][65] = 9'b111111111;
assign micromatri[9][66] = 9'b111111111;
assign micromatri[9][67] = 9'b111111111;
assign micromatri[9][68] = 9'b111111111;
assign micromatri[9][69] = 9'b111111111;
assign micromatri[9][70] = 9'b111111111;
assign micromatri[9][71] = 9'b111111111;
assign micromatri[9][72] = 9'b111111111;
assign micromatri[9][73] = 9'b111111111;
assign micromatri[9][74] = 9'b111111111;
assign micromatri[9][75] = 9'b111111111;
assign micromatri[9][76] = 9'b111111111;
assign micromatri[9][77] = 9'b111111111;
assign micromatri[9][78] = 9'b111111111;
assign micromatri[9][79] = 9'b111111111;
assign micromatri[9][80] = 9'b111111111;
assign micromatri[9][81] = 9'b111111111;
assign micromatri[9][82] = 9'b111111111;
assign micromatri[9][83] = 9'b111111111;
assign micromatri[9][84] = 9'b111111111;
assign micromatri[9][85] = 9'b111111111;
assign micromatri[9][86] = 9'b111111111;
assign micromatri[9][87] = 9'b111111111;
assign micromatri[9][88] = 9'b111111111;
assign micromatri[9][89] = 9'b111111111;
assign micromatri[9][90] = 9'b111111111;
assign micromatri[9][91] = 9'b111111111;
assign micromatri[9][92] = 9'b111111111;
assign micromatri[9][93] = 9'b111111111;
assign micromatri[9][94] = 9'b111111111;
assign micromatri[9][95] = 9'b111111111;
assign micromatri[9][96] = 9'b111111111;
assign micromatri[9][97] = 9'b111111111;
assign micromatri[9][98] = 9'b111111111;
assign micromatri[9][99] = 9'b111111111;
assign micromatri[10][0] = 9'b111111111;
assign micromatri[10][1] = 9'b111111111;
assign micromatri[10][2] = 9'b111111111;
assign micromatri[10][3] = 9'b111111111;
assign micromatri[10][4] = 9'b111111111;
assign micromatri[10][5] = 9'b111111111;
assign micromatri[10][6] = 9'b111111111;
assign micromatri[10][7] = 9'b111111111;
assign micromatri[10][8] = 9'b111111111;
assign micromatri[10][9] = 9'b111111111;
assign micromatri[10][10] = 9'b111111111;
assign micromatri[10][11] = 9'b111111111;
assign micromatri[10][12] = 9'b111111111;
assign micromatri[10][13] = 9'b111111111;
assign micromatri[10][14] = 9'b111111111;
assign micromatri[10][15] = 9'b111111111;
assign micromatri[10][16] = 9'b111111111;
assign micromatri[10][17] = 9'b111111111;
assign micromatri[10][18] = 9'b111111111;
assign micromatri[10][19] = 9'b111111111;
assign micromatri[10][20] = 9'b111111111;
assign micromatri[10][21] = 9'b111111111;
assign micromatri[10][22] = 9'b111111111;
assign micromatri[10][23] = 9'b111111111;
assign micromatri[10][24] = 9'b111111111;
assign micromatri[10][25] = 9'b111111111;
assign micromatri[10][26] = 9'b111111111;
assign micromatri[10][27] = 9'b111111111;
assign micromatri[10][28] = 9'b111111111;
assign micromatri[10][29] = 9'b111111111;
assign micromatri[10][30] = 9'b111111111;
assign micromatri[10][31] = 9'b111111111;
assign micromatri[10][32] = 9'b111111111;
assign micromatri[10][33] = 9'b111111111;
assign micromatri[10][34] = 9'b111111111;
assign micromatri[10][35] = 9'b111111111;
assign micromatri[10][36] = 9'b111111111;
assign micromatri[10][37] = 9'b111111111;
assign micromatri[10][38] = 9'b111111111;
assign micromatri[10][39] = 9'b111111111;
assign micromatri[10][40] = 9'b111111111;
assign micromatri[10][41] = 9'b111111111;
assign micromatri[10][42] = 9'b111111111;
assign micromatri[10][43] = 9'b111111111;
assign micromatri[10][44] = 9'b111111111;
assign micromatri[10][45] = 9'b111111111;
assign micromatri[10][46] = 9'b111111111;
assign micromatri[10][47] = 9'b111111111;
assign micromatri[10][48] = 9'b111111111;
assign micromatri[10][49] = 9'b111111111;
assign micromatri[10][50] = 9'b111111111;
assign micromatri[10][51] = 9'b111111111;
assign micromatri[10][52] = 9'b111111111;
assign micromatri[10][53] = 9'b111111111;
assign micromatri[10][54] = 9'b111111111;
assign micromatri[10][55] = 9'b111111111;
assign micromatri[10][56] = 9'b111111111;
assign micromatri[10][57] = 9'b111111111;
assign micromatri[10][58] = 9'b111111111;
assign micromatri[10][59] = 9'b111111111;
assign micromatri[10][60] = 9'b111111111;
assign micromatri[10][61] = 9'b111111111;
assign micromatri[10][62] = 9'b111111111;
assign micromatri[10][63] = 9'b111111111;
assign micromatri[10][64] = 9'b111111111;
assign micromatri[10][65] = 9'b111111111;
assign micromatri[10][66] = 9'b111111111;
assign micromatri[10][67] = 9'b111111111;
assign micromatri[10][68] = 9'b111111111;
assign micromatri[10][69] = 9'b111111111;
assign micromatri[10][70] = 9'b111111111;
assign micromatri[10][71] = 9'b111111111;
assign micromatri[10][72] = 9'b111111111;
assign micromatri[10][73] = 9'b111111111;
assign micromatri[10][74] = 9'b111111111;
assign micromatri[10][75] = 9'b111111111;
assign micromatri[10][76] = 9'b111111111;
assign micromatri[10][77] = 9'b111111111;
assign micromatri[10][78] = 9'b111111111;
assign micromatri[10][79] = 9'b111111111;
assign micromatri[10][80] = 9'b111111111;
assign micromatri[10][81] = 9'b111111111;
assign micromatri[10][82] = 9'b111111111;
assign micromatri[10][83] = 9'b111111111;
assign micromatri[10][84] = 9'b111111111;
assign micromatri[10][85] = 9'b111111111;
assign micromatri[10][86] = 9'b111111111;
assign micromatri[10][87] = 9'b111111111;
assign micromatri[10][88] = 9'b111111111;
assign micromatri[10][89] = 9'b111111111;
assign micromatri[10][90] = 9'b111111111;
assign micromatri[10][91] = 9'b111111111;
assign micromatri[10][92] = 9'b111111111;
assign micromatri[10][93] = 9'b111111111;
assign micromatri[10][94] = 9'b111111111;
assign micromatri[10][95] = 9'b111111111;
assign micromatri[10][96] = 9'b111111111;
assign micromatri[10][97] = 9'b111111111;
assign micromatri[10][98] = 9'b111111111;
assign micromatri[10][99] = 9'b111111111;
assign micromatri[11][0] = 9'b111111111;
assign micromatri[11][1] = 9'b111111111;
assign micromatri[11][2] = 9'b111111111;
assign micromatri[11][3] = 9'b111111111;
assign micromatri[11][4] = 9'b111111111;
assign micromatri[11][5] = 9'b111111111;
assign micromatri[11][6] = 9'b111111111;
assign micromatri[11][7] = 9'b111111111;
assign micromatri[11][8] = 9'b111111111;
assign micromatri[11][9] = 9'b111111111;
assign micromatri[11][10] = 9'b111111111;
assign micromatri[11][11] = 9'b111111111;
assign micromatri[11][12] = 9'b111111111;
assign micromatri[11][13] = 9'b111111111;
assign micromatri[11][14] = 9'b111111111;
assign micromatri[11][15] = 9'b111111111;
assign micromatri[11][16] = 9'b111111111;
assign micromatri[11][17] = 9'b111111111;
assign micromatri[11][18] = 9'b111111111;
assign micromatri[11][19] = 9'b111111111;
assign micromatri[11][20] = 9'b111111111;
assign micromatri[11][21] = 9'b111111111;
assign micromatri[11][22] = 9'b111111111;
assign micromatri[11][23] = 9'b111111111;
assign micromatri[11][24] = 9'b111111111;
assign micromatri[11][25] = 9'b111111111;
assign micromatri[11][26] = 9'b111111111;
assign micromatri[11][27] = 9'b111111111;
assign micromatri[11][28] = 9'b111111111;
assign micromatri[11][29] = 9'b111111111;
assign micromatri[11][30] = 9'b111111111;
assign micromatri[11][31] = 9'b111111111;
assign micromatri[11][32] = 9'b111111111;
assign micromatri[11][33] = 9'b111111111;
assign micromatri[11][34] = 9'b111111111;
assign micromatri[11][35] = 9'b111111111;
assign micromatri[11][36] = 9'b111111111;
assign micromatri[11][37] = 9'b111111111;
assign micromatri[11][38] = 9'b111111111;
assign micromatri[11][39] = 9'b111111111;
assign micromatri[11][40] = 9'b111111111;
assign micromatri[11][41] = 9'b111111111;
assign micromatri[11][42] = 9'b111111111;
assign micromatri[11][43] = 9'b111111111;
assign micromatri[11][44] = 9'b111111111;
assign micromatri[11][45] = 9'b111111111;
assign micromatri[11][46] = 9'b111111111;
assign micromatri[11][47] = 9'b111111111;
assign micromatri[11][48] = 9'b111111111;
assign micromatri[11][49] = 9'b111111111;
assign micromatri[11][50] = 9'b111111111;
assign micromatri[11][51] = 9'b111111111;
assign micromatri[11][52] = 9'b111111111;
assign micromatri[11][53] = 9'b111111111;
assign micromatri[11][54] = 9'b111111111;
assign micromatri[11][55] = 9'b111111111;
assign micromatri[11][56] = 9'b111111111;
assign micromatri[11][57] = 9'b111111111;
assign micromatri[11][58] = 9'b111111111;
assign micromatri[11][59] = 9'b111111111;
assign micromatri[11][60] = 9'b111111111;
assign micromatri[11][61] = 9'b111111111;
assign micromatri[11][62] = 9'b111111111;
assign micromatri[11][63] = 9'b111111111;
assign micromatri[11][64] = 9'b111111111;
assign micromatri[11][65] = 9'b111111111;
assign micromatri[11][66] = 9'b111111111;
assign micromatri[11][67] = 9'b111111111;
assign micromatri[11][68] = 9'b111111111;
assign micromatri[11][69] = 9'b111111111;
assign micromatri[11][70] = 9'b111111111;
assign micromatri[11][71] = 9'b111111111;
assign micromatri[11][72] = 9'b111111111;
assign micromatri[11][73] = 9'b111111111;
assign micromatri[11][74] = 9'b111111111;
assign micromatri[11][75] = 9'b111111111;
assign micromatri[11][76] = 9'b111111111;
assign micromatri[11][77] = 9'b111111111;
assign micromatri[11][78] = 9'b111111111;
assign micromatri[11][79] = 9'b111111111;
assign micromatri[11][80] = 9'b111111111;
assign micromatri[11][81] = 9'b111111111;
assign micromatri[11][82] = 9'b111111111;
assign micromatri[11][83] = 9'b111111111;
assign micromatri[11][84] = 9'b111111111;
assign micromatri[11][85] = 9'b111111111;
assign micromatri[11][86] = 9'b111111111;
assign micromatri[11][87] = 9'b111111111;
assign micromatri[11][88] = 9'b111111111;
assign micromatri[11][89] = 9'b111111111;
assign micromatri[11][90] = 9'b111111111;
assign micromatri[11][91] = 9'b111111111;
assign micromatri[11][92] = 9'b111111111;
assign micromatri[11][93] = 9'b111111111;
assign micromatri[11][94] = 9'b111111111;
assign micromatri[11][95] = 9'b111111111;
assign micromatri[11][96] = 9'b111111111;
assign micromatri[11][97] = 9'b111111111;
assign micromatri[11][98] = 9'b111111111;
assign micromatri[11][99] = 9'b111111111;
assign micromatri[12][0] = 9'b111111111;
assign micromatri[12][1] = 9'b111111111;
assign micromatri[12][2] = 9'b111111111;
assign micromatri[12][3] = 9'b111111111;
assign micromatri[12][4] = 9'b111111111;
assign micromatri[12][5] = 9'b111111111;
assign micromatri[12][6] = 9'b111111111;
assign micromatri[12][7] = 9'b111111111;
assign micromatri[12][8] = 9'b111111111;
assign micromatri[12][9] = 9'b111111111;
assign micromatri[12][10] = 9'b111111111;
assign micromatri[12][11] = 9'b111111111;
assign micromatri[12][12] = 9'b111111111;
assign micromatri[12][13] = 9'b111111111;
assign micromatri[12][14] = 9'b111111111;
assign micromatri[12][15] = 9'b111111111;
assign micromatri[12][16] = 9'b111111111;
assign micromatri[12][17] = 9'b111111111;
assign micromatri[12][18] = 9'b111111111;
assign micromatri[12][19] = 9'b111111111;
assign micromatri[12][20] = 9'b111111111;
assign micromatri[12][21] = 9'b111111111;
assign micromatri[12][22] = 9'b111111111;
assign micromatri[12][23] = 9'b111111111;
assign micromatri[12][24] = 9'b111111111;
assign micromatri[12][25] = 9'b111111111;
assign micromatri[12][26] = 9'b111111111;
assign micromatri[12][27] = 9'b111111111;
assign micromatri[12][28] = 9'b111111111;
assign micromatri[12][29] = 9'b111111111;
assign micromatri[12][30] = 9'b111111111;
assign micromatri[12][31] = 9'b111111111;
assign micromatri[12][32] = 9'b111111111;
assign micromatri[12][33] = 9'b111111111;
assign micromatri[12][34] = 9'b111111111;
assign micromatri[12][35] = 9'b111111111;
assign micromatri[12][36] = 9'b111111111;
assign micromatri[12][37] = 9'b111111111;
assign micromatri[12][38] = 9'b111111111;
assign micromatri[12][39] = 9'b111111111;
assign micromatri[12][40] = 9'b111111111;
assign micromatri[12][41] = 9'b111111111;
assign micromatri[12][42] = 9'b111111111;
assign micromatri[12][43] = 9'b111111111;
assign micromatri[12][44] = 9'b111111111;
assign micromatri[12][45] = 9'b111111111;
assign micromatri[12][46] = 9'b111111111;
assign micromatri[12][47] = 9'b111111111;
assign micromatri[12][48] = 9'b111111111;
assign micromatri[12][49] = 9'b111111111;
assign micromatri[12][50] = 9'b111111111;
assign micromatri[12][51] = 9'b111111111;
assign micromatri[12][52] = 9'b111111111;
assign micromatri[12][53] = 9'b111111111;
assign micromatri[12][54] = 9'b111111111;
assign micromatri[12][55] = 9'b111111111;
assign micromatri[12][56] = 9'b111111111;
assign micromatri[12][57] = 9'b111111111;
assign micromatri[12][58] = 9'b111111111;
assign micromatri[12][59] = 9'b111111111;
assign micromatri[12][60] = 9'b111111111;
assign micromatri[12][61] = 9'b111111111;
assign micromatri[12][62] = 9'b111111111;
assign micromatri[12][63] = 9'b111111111;
assign micromatri[12][64] = 9'b111111111;
assign micromatri[12][65] = 9'b111111111;
assign micromatri[12][66] = 9'b111111111;
assign micromatri[12][67] = 9'b111111111;
assign micromatri[12][68] = 9'b111111111;
assign micromatri[12][69] = 9'b111111111;
assign micromatri[12][70] = 9'b111111111;
assign micromatri[12][71] = 9'b111111111;
assign micromatri[12][72] = 9'b111111111;
assign micromatri[12][73] = 9'b111111111;
assign micromatri[12][74] = 9'b111111111;
assign micromatri[12][75] = 9'b111111111;
assign micromatri[12][76] = 9'b111111111;
assign micromatri[12][77] = 9'b111111111;
assign micromatri[12][78] = 9'b111111111;
assign micromatri[12][79] = 9'b111111111;
assign micromatri[12][80] = 9'b111111111;
assign micromatri[12][81] = 9'b111111111;
assign micromatri[12][82] = 9'b111111111;
assign micromatri[12][83] = 9'b111111111;
assign micromatri[12][84] = 9'b111111111;
assign micromatri[12][85] = 9'b111111111;
assign micromatri[12][86] = 9'b111111111;
assign micromatri[12][87] = 9'b111111111;
assign micromatri[12][88] = 9'b111111111;
assign micromatri[12][89] = 9'b111111111;
assign micromatri[12][90] = 9'b111111111;
assign micromatri[12][91] = 9'b111111111;
assign micromatri[12][92] = 9'b111111111;
assign micromatri[12][93] = 9'b111111111;
assign micromatri[12][94] = 9'b111111111;
assign micromatri[12][95] = 9'b111111111;
assign micromatri[12][96] = 9'b111111111;
assign micromatri[12][97] = 9'b111111111;
assign micromatri[12][98] = 9'b111111111;
assign micromatri[12][99] = 9'b111111111;
assign micromatri[13][0] = 9'b111111111;
assign micromatri[13][1] = 9'b111111111;
assign micromatri[13][2] = 9'b111111111;
assign micromatri[13][3] = 9'b111111111;
assign micromatri[13][4] = 9'b111111111;
assign micromatri[13][5] = 9'b111111111;
assign micromatri[13][6] = 9'b111111111;
assign micromatri[13][7] = 9'b111111111;
assign micromatri[13][8] = 9'b111111111;
assign micromatri[13][9] = 9'b111111111;
assign micromatri[13][10] = 9'b111111111;
assign micromatri[13][11] = 9'b111111111;
assign micromatri[13][12] = 9'b111111111;
assign micromatri[13][13] = 9'b111111111;
assign micromatri[13][14] = 9'b111111111;
assign micromatri[13][15] = 9'b111111111;
assign micromatri[13][16] = 9'b111111111;
assign micromatri[13][17] = 9'b111111111;
assign micromatri[13][18] = 9'b111111111;
assign micromatri[13][19] = 9'b111111111;
assign micromatri[13][20] = 9'b111111111;
assign micromatri[13][21] = 9'b111111111;
assign micromatri[13][22] = 9'b111111111;
assign micromatri[13][23] = 9'b111111111;
assign micromatri[13][24] = 9'b111111111;
assign micromatri[13][25] = 9'b111111111;
assign micromatri[13][26] = 9'b111111111;
assign micromatri[13][27] = 9'b111111111;
assign micromatri[13][28] = 9'b111111111;
assign micromatri[13][29] = 9'b111111111;
assign micromatri[13][30] = 9'b111111111;
assign micromatri[13][31] = 9'b111111111;
assign micromatri[13][32] = 9'b111111111;
assign micromatri[13][33] = 9'b111111111;
assign micromatri[13][34] = 9'b111111111;
assign micromatri[13][35] = 9'b111111111;
assign micromatri[13][36] = 9'b111111111;
assign micromatri[13][37] = 9'b111111111;
assign micromatri[13][38] = 9'b111111111;
assign micromatri[13][39] = 9'b111111111;
assign micromatri[13][40] = 9'b111111111;
assign micromatri[13][41] = 9'b111111111;
assign micromatri[13][42] = 9'b111111111;
assign micromatri[13][43] = 9'b111111111;
assign micromatri[13][44] = 9'b111111111;
assign micromatri[13][45] = 9'b111111111;
assign micromatri[13][46] = 9'b111111111;
assign micromatri[13][47] = 9'b111111111;
assign micromatri[13][48] = 9'b111111111;
assign micromatri[13][49] = 9'b111111111;
assign micromatri[13][50] = 9'b111111111;
assign micromatri[13][51] = 9'b111111111;
assign micromatri[13][52] = 9'b111111111;
assign micromatri[13][53] = 9'b111111111;
assign micromatri[13][54] = 9'b111111111;
assign micromatri[13][55] = 9'b111111111;
assign micromatri[13][56] = 9'b111111111;
assign micromatri[13][57] = 9'b111111111;
assign micromatri[13][58] = 9'b111111111;
assign micromatri[13][59] = 9'b111111111;
assign micromatri[13][60] = 9'b111111111;
assign micromatri[13][61] = 9'b111111111;
assign micromatri[13][62] = 9'b111111111;
assign micromatri[13][63] = 9'b111111111;
assign micromatri[13][64] = 9'b111111111;
assign micromatri[13][65] = 9'b111111111;
assign micromatri[13][66] = 9'b111111111;
assign micromatri[13][67] = 9'b111111111;
assign micromatri[13][68] = 9'b111111111;
assign micromatri[13][69] = 9'b111111111;
assign micromatri[13][70] = 9'b111111111;
assign micromatri[13][71] = 9'b111111111;
assign micromatri[13][72] = 9'b111111111;
assign micromatri[13][73] = 9'b111111111;
assign micromatri[13][74] = 9'b111111111;
assign micromatri[13][75] = 9'b111111111;
assign micromatri[13][76] = 9'b111111111;
assign micromatri[13][77] = 9'b111111111;
assign micromatri[13][78] = 9'b111111111;
assign micromatri[13][79] = 9'b111111111;
assign micromatri[13][80] = 9'b111111111;
assign micromatri[13][81] = 9'b111111111;
assign micromatri[13][82] = 9'b111111111;
assign micromatri[13][83] = 9'b111111111;
assign micromatri[13][84] = 9'b111111111;
assign micromatri[13][85] = 9'b111111111;
assign micromatri[13][86] = 9'b111111111;
assign micromatri[13][87] = 9'b111111111;
assign micromatri[13][88] = 9'b111111111;
assign micromatri[13][89] = 9'b111111111;
assign micromatri[13][90] = 9'b111111111;
assign micromatri[13][91] = 9'b111111111;
assign micromatri[13][92] = 9'b111111111;
assign micromatri[13][93] = 9'b111111111;
assign micromatri[13][94] = 9'b111111111;
assign micromatri[13][95] = 9'b111111111;
assign micromatri[13][96] = 9'b111111111;
assign micromatri[13][97] = 9'b111111111;
assign micromatri[13][98] = 9'b111111111;
assign micromatri[13][99] = 9'b111111111;
assign micromatri[14][0] = 9'b111111111;
assign micromatri[14][1] = 9'b111111111;
assign micromatri[14][2] = 9'b111111111;
assign micromatri[14][3] = 9'b111111111;
assign micromatri[14][4] = 9'b111111111;
assign micromatri[14][5] = 9'b111111111;
assign micromatri[14][6] = 9'b111111111;
assign micromatri[14][7] = 9'b111111111;
assign micromatri[14][8] = 9'b111111111;
assign micromatri[14][9] = 9'b111111111;
assign micromatri[14][10] = 9'b111111111;
assign micromatri[14][11] = 9'b111111111;
assign micromatri[14][12] = 9'b111111111;
assign micromatri[14][13] = 9'b111111111;
assign micromatri[14][14] = 9'b111111111;
assign micromatri[14][15] = 9'b111111111;
assign micromatri[14][16] = 9'b111111111;
assign micromatri[14][17] = 9'b111111111;
assign micromatri[14][18] = 9'b111111111;
assign micromatri[14][19] = 9'b111111111;
assign micromatri[14][20] = 9'b111111111;
assign micromatri[14][21] = 9'b111111111;
assign micromatri[14][22] = 9'b111111111;
assign micromatri[14][23] = 9'b111111111;
assign micromatri[14][24] = 9'b111111111;
assign micromatri[14][25] = 9'b111111111;
assign micromatri[14][26] = 9'b111111111;
assign micromatri[14][27] = 9'b111111111;
assign micromatri[14][28] = 9'b111111111;
assign micromatri[14][29] = 9'b111111111;
assign micromatri[14][30] = 9'b111111111;
assign micromatri[14][31] = 9'b111111111;
assign micromatri[14][32] = 9'b111111111;
assign micromatri[14][33] = 9'b111111111;
assign micromatri[14][34] = 9'b111111111;
assign micromatri[14][35] = 9'b111111111;
assign micromatri[14][36] = 9'b111111111;
assign micromatri[14][37] = 9'b111111111;
assign micromatri[14][38] = 9'b111111111;
assign micromatri[14][39] = 9'b111111111;
assign micromatri[14][40] = 9'b111111111;
assign micromatri[14][41] = 9'b111111111;
assign micromatri[14][42] = 9'b111111111;
assign micromatri[14][43] = 9'b111111111;
assign micromatri[14][44] = 9'b111111111;
assign micromatri[14][45] = 9'b111111111;
assign micromatri[14][46] = 9'b111111111;
assign micromatri[14][47] = 9'b111111111;
assign micromatri[14][48] = 9'b111111111;
assign micromatri[14][49] = 9'b111111111;
assign micromatri[14][50] = 9'b111111111;
assign micromatri[14][51] = 9'b111111111;
assign micromatri[14][52] = 9'b111111111;
assign micromatri[14][53] = 9'b111111111;
assign micromatri[14][54] = 9'b111111111;
assign micromatri[14][55] = 9'b111111111;
assign micromatri[14][56] = 9'b111111111;
assign micromatri[14][57] = 9'b111111111;
assign micromatri[14][58] = 9'b111111111;
assign micromatri[14][59] = 9'b111111111;
assign micromatri[14][60] = 9'b111111111;
assign micromatri[14][61] = 9'b111111111;
assign micromatri[14][62] = 9'b111111111;
assign micromatri[14][63] = 9'b111111111;
assign micromatri[14][64] = 9'b111111111;
assign micromatri[14][65] = 9'b111111111;
assign micromatri[14][66] = 9'b111111111;
assign micromatri[14][67] = 9'b111111111;
assign micromatri[14][68] = 9'b111111111;
assign micromatri[14][69] = 9'b111111111;
assign micromatri[14][70] = 9'b111111111;
assign micromatri[14][71] = 9'b111111111;
assign micromatri[14][72] = 9'b111111111;
assign micromatri[14][73] = 9'b111111111;
assign micromatri[14][74] = 9'b111111111;
assign micromatri[14][75] = 9'b111111111;
assign micromatri[14][76] = 9'b111111111;
assign micromatri[14][77] = 9'b111111111;
assign micromatri[14][78] = 9'b111111111;
assign micromatri[14][79] = 9'b111111111;
assign micromatri[14][80] = 9'b111111111;
assign micromatri[14][81] = 9'b111111111;
assign micromatri[14][82] = 9'b111111111;
assign micromatri[14][83] = 9'b111111111;
assign micromatri[14][84] = 9'b111111111;
assign micromatri[14][85] = 9'b111111111;
assign micromatri[14][86] = 9'b111111111;
assign micromatri[14][87] = 9'b111111111;
assign micromatri[14][88] = 9'b111111111;
assign micromatri[14][89] = 9'b111111111;
assign micromatri[14][90] = 9'b111111111;
assign micromatri[14][91] = 9'b111111111;
assign micromatri[14][92] = 9'b111111111;
assign micromatri[14][93] = 9'b111111111;
assign micromatri[14][94] = 9'b111111111;
assign micromatri[14][95] = 9'b111111111;
assign micromatri[14][96] = 9'b111111111;
assign micromatri[14][97] = 9'b111111111;
assign micromatri[14][98] = 9'b111111111;
assign micromatri[14][99] = 9'b111111111;
assign micromatri[15][0] = 9'b111111111;
assign micromatri[15][1] = 9'b111111111;
assign micromatri[15][2] = 9'b111111111;
assign micromatri[15][3] = 9'b111111111;
assign micromatri[15][4] = 9'b111111111;
assign micromatri[15][5] = 9'b111111111;
assign micromatri[15][6] = 9'b111111111;
assign micromatri[15][7] = 9'b111111111;
assign micromatri[15][8] = 9'b111111111;
assign micromatri[15][9] = 9'b111111111;
assign micromatri[15][10] = 9'b111111111;
assign micromatri[15][11] = 9'b111111111;
assign micromatri[15][12] = 9'b111111111;
assign micromatri[15][13] = 9'b111111111;
assign micromatri[15][14] = 9'b111111111;
assign micromatri[15][15] = 9'b111111111;
assign micromatri[15][16] = 9'b111111111;
assign micromatri[15][17] = 9'b111111111;
assign micromatri[15][18] = 9'b111111111;
assign micromatri[15][19] = 9'b111111111;
assign micromatri[15][20] = 9'b111111111;
assign micromatri[15][21] = 9'b111111111;
assign micromatri[15][22] = 9'b111111111;
assign micromatri[15][23] = 9'b111111111;
assign micromatri[15][24] = 9'b111111111;
assign micromatri[15][25] = 9'b111111111;
assign micromatri[15][26] = 9'b111111111;
assign micromatri[15][27] = 9'b111111111;
assign micromatri[15][28] = 9'b111111111;
assign micromatri[15][29] = 9'b111111111;
assign micromatri[15][30] = 9'b111111111;
assign micromatri[15][31] = 9'b111111111;
assign micromatri[15][32] = 9'b111111111;
assign micromatri[15][33] = 9'b111111111;
assign micromatri[15][34] = 9'b111111111;
assign micromatri[15][35] = 9'b111111111;
assign micromatri[15][36] = 9'b111111111;
assign micromatri[15][37] = 9'b111111111;
assign micromatri[15][38] = 9'b111111111;
assign micromatri[15][39] = 9'b111111111;
assign micromatri[15][40] = 9'b111111111;
assign micromatri[15][41] = 9'b111111111;
assign micromatri[15][42] = 9'b111111111;
assign micromatri[15][43] = 9'b111111111;
assign micromatri[15][44] = 9'b111111111;
assign micromatri[15][45] = 9'b111111111;
assign micromatri[15][46] = 9'b111111111;
assign micromatri[15][47] = 9'b111111111;
assign micromatri[15][48] = 9'b111111111;
assign micromatri[15][49] = 9'b111111111;
assign micromatri[15][50] = 9'b111111111;
assign micromatri[15][51] = 9'b111111111;
assign micromatri[15][52] = 9'b111111111;
assign micromatri[15][53] = 9'b111111111;
assign micromatri[15][54] = 9'b111111111;
assign micromatri[15][55] = 9'b111111111;
assign micromatri[15][56] = 9'b111111111;
assign micromatri[15][57] = 9'b111111111;
assign micromatri[15][58] = 9'b111111111;
assign micromatri[15][59] = 9'b111111111;
assign micromatri[15][60] = 9'b111111111;
assign micromatri[15][61] = 9'b110010001;
assign micromatri[15][62] = 9'b110010010;
assign micromatri[15][63] = 9'b110010001;
assign micromatri[15][64] = 9'b111111111;
assign micromatri[15][65] = 9'b111111111;
assign micromatri[15][66] = 9'b111111111;
assign micromatri[15][67] = 9'b111111111;
assign micromatri[15][68] = 9'b111111111;
assign micromatri[15][69] = 9'b111111111;
assign micromatri[15][70] = 9'b111111111;
assign micromatri[15][71] = 9'b111111111;
assign micromatri[15][72] = 9'b111111111;
assign micromatri[15][73] = 9'b111111111;
assign micromatri[15][74] = 9'b111111111;
assign micromatri[15][75] = 9'b111111111;
assign micromatri[15][76] = 9'b111111111;
assign micromatri[15][77] = 9'b111111111;
assign micromatri[15][78] = 9'b111111111;
assign micromatri[15][79] = 9'b111111111;
assign micromatri[15][80] = 9'b111111111;
assign micromatri[15][81] = 9'b111111111;
assign micromatri[15][82] = 9'b111111111;
assign micromatri[15][83] = 9'b111111111;
assign micromatri[15][84] = 9'b111111111;
assign micromatri[15][85] = 9'b111111111;
assign micromatri[15][86] = 9'b111111111;
assign micromatri[15][87] = 9'b111111111;
assign micromatri[15][88] = 9'b111111111;
assign micromatri[15][89] = 9'b111111111;
assign micromatri[15][90] = 9'b111111111;
assign micromatri[15][91] = 9'b111111111;
assign micromatri[15][92] = 9'b111111111;
assign micromatri[15][93] = 9'b111111111;
assign micromatri[15][94] = 9'b111111111;
assign micromatri[15][95] = 9'b111111111;
assign micromatri[15][96] = 9'b111111111;
assign micromatri[15][97] = 9'b111111111;
assign micromatri[15][98] = 9'b111111111;
assign micromatri[15][99] = 9'b111111111;
assign micromatri[16][0] = 9'b111111111;
assign micromatri[16][1] = 9'b111111111;
assign micromatri[16][2] = 9'b111111111;
assign micromatri[16][3] = 9'b111111111;
assign micromatri[16][4] = 9'b111111111;
assign micromatri[16][5] = 9'b111111111;
assign micromatri[16][6] = 9'b111111111;
assign micromatri[16][7] = 9'b111111111;
assign micromatri[16][8] = 9'b111111111;
assign micromatri[16][9] = 9'b111111111;
assign micromatri[16][10] = 9'b111111111;
assign micromatri[16][11] = 9'b111111111;
assign micromatri[16][12] = 9'b111111111;
assign micromatri[16][13] = 9'b111111111;
assign micromatri[16][14] = 9'b111111111;
assign micromatri[16][15] = 9'b111111111;
assign micromatri[16][16] = 9'b111111111;
assign micromatri[16][17] = 9'b111111111;
assign micromatri[16][18] = 9'b111111111;
assign micromatri[16][19] = 9'b111111111;
assign micromatri[16][20] = 9'b111111111;
assign micromatri[16][21] = 9'b111111111;
assign micromatri[16][22] = 9'b111111111;
assign micromatri[16][23] = 9'b111111111;
assign micromatri[16][24] = 9'b111111111;
assign micromatri[16][25] = 9'b110110110;
assign micromatri[16][26] = 9'b110010001;
assign micromatri[16][27] = 9'b110010001;
assign micromatri[16][28] = 9'b110001101;
assign micromatri[16][29] = 9'b111111111;
assign micromatri[16][30] = 9'b111111111;
assign micromatri[16][31] = 9'b111111111;
assign micromatri[16][32] = 9'b101101101;
assign micromatri[16][33] = 9'b110010010;
assign micromatri[16][34] = 9'b110010010;
assign micromatri[16][35] = 9'b111111111;
assign micromatri[16][36] = 9'b111111111;
assign micromatri[16][37] = 9'b111111111;
assign micromatri[16][38] = 9'b111111111;
assign micromatri[16][39] = 9'b111111111;
assign micromatri[16][40] = 9'b111111111;
assign micromatri[16][41] = 9'b111111111;
assign micromatri[16][42] = 9'b111111111;
assign micromatri[16][43] = 9'b111111111;
assign micromatri[16][44] = 9'b111111111;
assign micromatri[16][45] = 9'b111111111;
assign micromatri[16][46] = 9'b111111111;
assign micromatri[16][47] = 9'b110010010;
assign micromatri[16][48] = 9'b110010110;
assign micromatri[16][49] = 9'b110010110;
assign micromatri[16][50] = 9'b110010110;
assign micromatri[16][51] = 9'b110010010;
assign micromatri[16][52] = 9'b110010010;
assign micromatri[16][53] = 9'b111111111;
assign micromatri[16][54] = 9'b111111111;
assign micromatri[16][55] = 9'b111111111;
assign micromatri[16][56] = 9'b111111111;
assign micromatri[16][57] = 9'b111111111;
assign micromatri[16][58] = 9'b111111111;
assign micromatri[16][59] = 9'b111111111;
assign micromatri[16][60] = 9'b110001101;
assign micromatri[16][61] = 9'b111110111;
assign micromatri[16][62] = 9'b111110111;
assign micromatri[16][63] = 9'b111110111;
assign micromatri[16][64] = 9'b110001101;
assign micromatri[16][65] = 9'b111111111;
assign micromatri[16][66] = 9'b111111111;
assign micromatri[16][67] = 9'b111111111;
assign micromatri[16][68] = 9'b111111111;
assign micromatri[16][69] = 9'b111111111;
assign micromatri[16][70] = 9'b111111111;
assign micromatri[16][71] = 9'b110010001;
assign micromatri[16][72] = 9'b110001110;
assign micromatri[16][73] = 9'b110010010;
assign micromatri[16][74] = 9'b110110010;
assign micromatri[16][75] = 9'b110110010;
assign micromatri[16][76] = 9'b110010010;
assign micromatri[16][77] = 9'b110001101;
assign micromatri[16][78] = 9'b110010010;
assign micromatri[16][79] = 9'b111111111;
assign micromatri[16][80] = 9'b111111111;
assign micromatri[16][81] = 9'b111111111;
assign micromatri[16][82] = 9'b111111111;
assign micromatri[16][83] = 9'b111111111;
assign micromatri[16][84] = 9'b111111111;
assign micromatri[16][85] = 9'b111111111;
assign micromatri[16][86] = 9'b111111111;
assign micromatri[16][87] = 9'b111111111;
assign micromatri[16][88] = 9'b111111111;
assign micromatri[16][89] = 9'b111111111;
assign micromatri[16][90] = 9'b111111111;
assign micromatri[16][91] = 9'b111111111;
assign micromatri[16][92] = 9'b111111111;
assign micromatri[16][93] = 9'b111111111;
assign micromatri[16][94] = 9'b111111111;
assign micromatri[16][95] = 9'b111111111;
assign micromatri[16][96] = 9'b111111111;
assign micromatri[16][97] = 9'b111111111;
assign micromatri[16][98] = 9'b111111111;
assign micromatri[16][99] = 9'b111111111;
assign micromatri[17][0] = 9'b111111111;
assign micromatri[17][1] = 9'b111111111;
assign micromatri[17][2] = 9'b111111111;
assign micromatri[17][3] = 9'b111111111;
assign micromatri[17][4] = 9'b111111111;
assign micromatri[17][5] = 9'b111111111;
assign micromatri[17][6] = 9'b111111111;
assign micromatri[17][7] = 9'b111111111;
assign micromatri[17][8] = 9'b111111111;
assign micromatri[17][9] = 9'b111111111;
assign micromatri[17][10] = 9'b111111111;
assign micromatri[17][11] = 9'b111111111;
assign micromatri[17][12] = 9'b111111111;
assign micromatri[17][13] = 9'b111111111;
assign micromatri[17][14] = 9'b111111111;
assign micromatri[17][15] = 9'b111111111;
assign micromatri[17][16] = 9'b111111111;
assign micromatri[17][17] = 9'b111111111;
assign micromatri[17][18] = 9'b111111111;
assign micromatri[17][19] = 9'b111111111;
assign micromatri[17][20] = 9'b111111111;
assign micromatri[17][21] = 9'b111111111;
assign micromatri[17][22] = 9'b110010010;
assign micromatri[17][23] = 9'b110010001;
assign micromatri[17][24] = 9'b110110010;
assign micromatri[17][25] = 9'b111110010;
assign micromatri[17][26] = 9'b111110011;
assign micromatri[17][27] = 9'b111110111;
assign micromatri[17][28] = 9'b111110111;
assign micromatri[17][29] = 9'b110001101;
assign micromatri[17][30] = 9'b111111111;
assign micromatri[17][31] = 9'b110110110;
assign micromatri[17][32] = 9'b110110011;
assign micromatri[17][33] = 9'b111110111;
assign micromatri[17][34] = 9'b110110011;
assign micromatri[17][35] = 9'b110010010;
assign micromatri[17][36] = 9'b110001101;
assign micromatri[17][37] = 9'b110010010;
assign micromatri[17][38] = 9'b111111111;
assign micromatri[17][39] = 9'b111111111;
assign micromatri[17][40] = 9'b111111111;
assign micromatri[17][41] = 9'b110001101;
assign micromatri[17][42] = 9'b110110011;
assign micromatri[17][43] = 9'b110010010;
assign micromatri[17][44] = 9'b110010010;
assign micromatri[17][45] = 9'b110010001;
assign micromatri[17][46] = 9'b111111111;
assign micromatri[17][47] = 9'b110010010;
assign micromatri[17][48] = 9'b111111111;
assign micromatri[17][49] = 9'b111111111;
assign micromatri[17][50] = 9'b111111111;
assign micromatri[17][51] = 9'b111111111;
assign micromatri[17][52] = 9'b110010010;
assign micromatri[17][53] = 9'b111111111;
assign micromatri[17][54] = 9'b111111111;
assign micromatri[17][55] = 9'b111111111;
assign micromatri[17][56] = 9'b111111111;
assign micromatri[17][57] = 9'b111111111;
assign micromatri[17][58] = 9'b111111111;
assign micromatri[17][59] = 9'b110010001;
assign micromatri[17][60] = 9'b111110111;
assign micromatri[17][61] = 9'b111110111;
assign micromatri[17][62] = 9'b111110111;
assign micromatri[17][63] = 9'b111111111;
assign micromatri[17][64] = 9'b111110011;
assign micromatri[17][65] = 9'b101101101;
assign micromatri[17][66] = 9'b111111111;
assign micromatri[17][67] = 9'b111111111;
assign micromatri[17][68] = 9'b111111111;
assign micromatri[17][69] = 9'b110010001;
assign micromatri[17][70] = 9'b110001110;
assign micromatri[17][71] = 9'b111110011;
assign micromatri[17][72] = 9'b111110111;
assign micromatri[17][73] = 9'b111110111;
assign micromatri[17][74] = 9'b111110111;
assign micromatri[17][75] = 9'b111110111;
assign micromatri[17][76] = 9'b111110111;
assign micromatri[17][77] = 9'b111110111;
assign micromatri[17][78] = 9'b110110010;
assign micromatri[17][79] = 9'b110001101;
assign micromatri[17][80] = 9'b111111111;
assign micromatri[17][81] = 9'b111111111;
assign micromatri[17][82] = 9'b111111111;
assign micromatri[17][83] = 9'b111111111;
assign micromatri[17][84] = 9'b111111111;
assign micromatri[17][85] = 9'b111111111;
assign micromatri[17][86] = 9'b111111111;
assign micromatri[17][87] = 9'b111111111;
assign micromatri[17][88] = 9'b111111111;
assign micromatri[17][89] = 9'b111111111;
assign micromatri[17][90] = 9'b111111111;
assign micromatri[17][91] = 9'b111111111;
assign micromatri[17][92] = 9'b111111111;
assign micromatri[17][93] = 9'b111111111;
assign micromatri[17][94] = 9'b111111111;
assign micromatri[17][95] = 9'b111111111;
assign micromatri[17][96] = 9'b111111111;
assign micromatri[17][97] = 9'b111111111;
assign micromatri[17][98] = 9'b111111111;
assign micromatri[17][99] = 9'b111111111;
assign micromatri[18][0] = 9'b111111111;
assign micromatri[18][1] = 9'b111111111;
assign micromatri[18][2] = 9'b111111111;
assign micromatri[18][3] = 9'b111111111;
assign micromatri[18][4] = 9'b111111111;
assign micromatri[18][5] = 9'b111111111;
assign micromatri[18][6] = 9'b111111111;
assign micromatri[18][7] = 9'b111111111;
assign micromatri[18][8] = 9'b111111111;
assign micromatri[18][9] = 9'b111111111;
assign micromatri[18][10] = 9'b111111111;
assign micromatri[18][11] = 9'b111111111;
assign micromatri[18][12] = 9'b111111111;
assign micromatri[18][13] = 9'b111111111;
assign micromatri[18][14] = 9'b111111111;
assign micromatri[18][15] = 9'b111111111;
assign micromatri[18][16] = 9'b111111111;
assign micromatri[18][17] = 9'b111111111;
assign micromatri[18][18] = 9'b111111111;
assign micromatri[18][19] = 9'b111111111;
assign micromatri[18][20] = 9'b111111111;
assign micromatri[18][21] = 9'b111111111;
assign micromatri[18][22] = 9'b110001101;
assign micromatri[18][23] = 9'b111110111;
assign micromatri[18][24] = 9'b111111111;
assign micromatri[18][25] = 9'b111111111;
assign micromatri[18][26] = 9'b111110111;
assign micromatri[18][27] = 9'b111110111;
assign micromatri[18][28] = 9'b111111111;
assign micromatri[18][29] = 9'b110001101;
assign micromatri[18][30] = 9'b110110010;
assign micromatri[18][31] = 9'b110010010;
assign micromatri[18][32] = 9'b111110011;
assign micromatri[18][33] = 9'b111110111;
assign micromatri[18][34] = 9'b111110111;
assign micromatri[18][35] = 9'b111110111;
assign micromatri[18][36] = 9'b111110111;
assign micromatri[18][37] = 9'b111110011;
assign micromatri[18][38] = 9'b110001101;
assign micromatri[18][39] = 9'b111111111;
assign micromatri[18][40] = 9'b111111111;
assign micromatri[18][41] = 9'b110010010;
assign micromatri[18][42] = 9'b111110111;
assign micromatri[18][43] = 9'b111110111;
assign micromatri[18][44] = 9'b111110111;
assign micromatri[18][45] = 9'b110010010;
assign micromatri[18][46] = 9'b110010010;
assign micromatri[18][47] = 9'b110010010;
assign micromatri[18][48] = 9'b111111111;
assign micromatri[18][49] = 9'b111111111;
assign micromatri[18][50] = 9'b111111111;
assign micromatri[18][51] = 9'b111111111;
assign micromatri[18][52] = 9'b110010010;
assign micromatri[18][53] = 9'b110111111;
assign micromatri[18][54] = 9'b111111111;
assign micromatri[18][55] = 9'b111111111;
assign micromatri[18][56] = 9'b111111111;
assign micromatri[18][57] = 9'b111111111;
assign micromatri[18][58] = 9'b111111111;
assign micromatri[18][59] = 9'b110010010;
assign micromatri[18][60] = 9'b111110111;
assign micromatri[18][61] = 9'b111110111;
assign micromatri[18][62] = 9'b111110111;
assign micromatri[18][63] = 9'b111110111;
assign micromatri[18][64] = 9'b111110111;
assign micromatri[18][65] = 9'b110010001;
assign micromatri[18][66] = 9'b111111111;
assign micromatri[18][67] = 9'b111111111;
assign micromatri[18][68] = 9'b110010001;
assign micromatri[18][69] = 9'b110110011;
assign micromatri[18][70] = 9'b111110111;
assign micromatri[18][71] = 9'b111110111;
assign micromatri[18][72] = 9'b111110111;
assign micromatri[18][73] = 9'b111110111;
assign micromatri[18][74] = 9'b111110111;
assign micromatri[18][75] = 9'b111110111;
assign micromatri[18][76] = 9'b111110111;
assign micromatri[18][77] = 9'b111110111;
assign micromatri[18][78] = 9'b111110111;
assign micromatri[18][79] = 9'b111110011;
assign micromatri[18][80] = 9'b110001101;
assign micromatri[18][81] = 9'b111111111;
assign micromatri[18][82] = 9'b111111111;
assign micromatri[18][83] = 9'b111111111;
assign micromatri[18][84] = 9'b111111111;
assign micromatri[18][85] = 9'b111111111;
assign micromatri[18][86] = 9'b111111111;
assign micromatri[18][87] = 9'b111111111;
assign micromatri[18][88] = 9'b111111111;
assign micromatri[18][89] = 9'b111111111;
assign micromatri[18][90] = 9'b111111111;
assign micromatri[18][91] = 9'b111111111;
assign micromatri[18][92] = 9'b111111111;
assign micromatri[18][93] = 9'b111111111;
assign micromatri[18][94] = 9'b111111111;
assign micromatri[18][95] = 9'b111111111;
assign micromatri[18][96] = 9'b111111111;
assign micromatri[18][97] = 9'b111111111;
assign micromatri[18][98] = 9'b111111111;
assign micromatri[18][99] = 9'b111111111;
assign micromatri[19][0] = 9'b111111111;
assign micromatri[19][1] = 9'b111111111;
assign micromatri[19][2] = 9'b111111111;
assign micromatri[19][3] = 9'b111111111;
assign micromatri[19][4] = 9'b111111111;
assign micromatri[19][5] = 9'b111111111;
assign micromatri[19][6] = 9'b111111111;
assign micromatri[19][7] = 9'b111111111;
assign micromatri[19][8] = 9'b111111111;
assign micromatri[19][9] = 9'b111111111;
assign micromatri[19][10] = 9'b111111111;
assign micromatri[19][11] = 9'b111111111;
assign micromatri[19][12] = 9'b111111111;
assign micromatri[19][13] = 9'b111111111;
assign micromatri[19][14] = 9'b111111111;
assign micromatri[19][15] = 9'b111111111;
assign micromatri[19][16] = 9'b111111111;
assign micromatri[19][17] = 9'b111111111;
assign micromatri[19][18] = 9'b111111111;
assign micromatri[19][19] = 9'b111111111;
assign micromatri[19][20] = 9'b111111111;
assign micromatri[19][21] = 9'b111111111;
assign micromatri[19][22] = 9'b110110110;
assign micromatri[19][23] = 9'b111110010;
assign micromatri[19][24] = 9'b111111111;
assign micromatri[19][25] = 9'b111110111;
assign micromatri[19][26] = 9'b111110111;
assign micromatri[19][27] = 9'b111110111;
assign micromatri[19][28] = 9'b111111111;
assign micromatri[19][29] = 9'b111110010;
assign micromatri[19][30] = 9'b110010010;
assign micromatri[19][31] = 9'b110001101;
assign micromatri[19][32] = 9'b111110011;
assign micromatri[19][33] = 9'b111110111;
assign micromatri[19][34] = 9'b111110111;
assign micromatri[19][35] = 9'b111110111;
assign micromatri[19][36] = 9'b111110111;
assign micromatri[19][37] = 9'b111110111;
assign micromatri[19][38] = 9'b110001110;
assign micromatri[19][39] = 9'b110110110;
assign micromatri[19][40] = 9'b111111111;
assign micromatri[19][41] = 9'b110010010;
assign micromatri[19][42] = 9'b111110011;
assign micromatri[19][43] = 9'b111110111;
assign micromatri[19][44] = 9'b111110111;
assign micromatri[19][45] = 9'b110010010;
assign micromatri[19][46] = 9'b110110010;
assign micromatri[19][47] = 9'b110010010;
assign micromatri[19][48] = 9'b111111111;
assign micromatri[19][49] = 9'b111111111;
assign micromatri[19][50] = 9'b111111111;
assign micromatri[19][51] = 9'b111111111;
assign micromatri[19][52] = 9'b110010110;
assign micromatri[19][53] = 9'b111111111;
assign micromatri[19][54] = 9'b111111111;
assign micromatri[19][55] = 9'b111111111;
assign micromatri[19][56] = 9'b111111111;
assign micromatri[19][57] = 9'b111111111;
assign micromatri[19][58] = 9'b111111111;
assign micromatri[19][59] = 9'b110010001;
assign micromatri[19][60] = 9'b111110010;
assign micromatri[19][61] = 9'b111111111;
assign micromatri[19][62] = 9'b111110111;
assign micromatri[19][63] = 9'b111111111;
assign micromatri[19][64] = 9'b111110010;
assign micromatri[19][65] = 9'b110110010;
assign micromatri[19][66] = 9'b111111111;
assign micromatri[19][67] = 9'b110010001;
assign micromatri[19][68] = 9'b110110011;
assign micromatri[19][69] = 9'b111110111;
assign micromatri[19][70] = 9'b111110111;
assign micromatri[19][71] = 9'b111110111;
assign micromatri[19][72] = 9'b111110111;
assign micromatri[19][73] = 9'b111110111;
assign micromatri[19][74] = 9'b111110111;
assign micromatri[19][75] = 9'b111110111;
assign micromatri[19][76] = 9'b111110111;
assign micromatri[19][77] = 9'b111110111;
assign micromatri[19][78] = 9'b111110111;
assign micromatri[19][79] = 9'b111110111;
assign micromatri[19][80] = 9'b110110011;
assign micromatri[19][81] = 9'b101101101;
assign micromatri[19][82] = 9'b111111111;
assign micromatri[19][83] = 9'b111111111;
assign micromatri[19][84] = 9'b111111111;
assign micromatri[19][85] = 9'b111111111;
assign micromatri[19][86] = 9'b111111111;
assign micromatri[19][87] = 9'b111111111;
assign micromatri[19][88] = 9'b111111111;
assign micromatri[19][89] = 9'b111111111;
assign micromatri[19][90] = 9'b111111111;
assign micromatri[19][91] = 9'b111111111;
assign micromatri[19][92] = 9'b111111111;
assign micromatri[19][93] = 9'b111111111;
assign micromatri[19][94] = 9'b111111111;
assign micromatri[19][95] = 9'b111111111;
assign micromatri[19][96] = 9'b111111111;
assign micromatri[19][97] = 9'b111111111;
assign micromatri[19][98] = 9'b111111111;
assign micromatri[19][99] = 9'b111111111;
assign micromatri[20][0] = 9'b111111111;
assign micromatri[20][1] = 9'b111111111;
assign micromatri[20][2] = 9'b111111111;
assign micromatri[20][3] = 9'b111111111;
assign micromatri[20][4] = 9'b111111111;
assign micromatri[20][5] = 9'b111111111;
assign micromatri[20][6] = 9'b111111111;
assign micromatri[20][7] = 9'b111111111;
assign micromatri[20][8] = 9'b111111111;
assign micromatri[20][9] = 9'b111111111;
assign micromatri[20][10] = 9'b111111111;
assign micromatri[20][11] = 9'b111111111;
assign micromatri[20][12] = 9'b111111111;
assign micromatri[20][13] = 9'b111111111;
assign micromatri[20][14] = 9'b111111111;
assign micromatri[20][15] = 9'b111111111;
assign micromatri[20][16] = 9'b111111111;
assign micromatri[20][17] = 9'b111111111;
assign micromatri[20][18] = 9'b111111111;
assign micromatri[20][19] = 9'b111111111;
assign micromatri[20][20] = 9'b111111111;
assign micromatri[20][21] = 9'b111111111;
assign micromatri[20][22] = 9'b111111111;
assign micromatri[20][23] = 9'b110001101;
assign micromatri[20][24] = 9'b111111111;
assign micromatri[20][25] = 9'b111110111;
assign micromatri[20][26] = 9'b111110111;
assign micromatri[20][27] = 9'b111110111;
assign micromatri[20][28] = 9'b111110111;
assign micromatri[20][29] = 9'b111110011;
assign micromatri[20][30] = 9'b110110010;
assign micromatri[20][31] = 9'b110010001;
assign micromatri[20][32] = 9'b111110011;
assign micromatri[20][33] = 9'b111110111;
assign micromatri[20][34] = 9'b111110111;
assign micromatri[20][35] = 9'b111110111;
assign micromatri[20][36] = 9'b111110111;
assign micromatri[20][37] = 9'b111110111;
assign micromatri[20][38] = 9'b110010010;
assign micromatri[20][39] = 9'b111111111;
assign micromatri[20][40] = 9'b111111111;
assign micromatri[20][41] = 9'b110010010;
assign micromatri[20][42] = 9'b111110011;
assign micromatri[20][43] = 9'b111110111;
assign micromatri[20][44] = 9'b111110111;
assign micromatri[20][45] = 9'b110010010;
assign micromatri[20][46] = 9'b111110111;
assign micromatri[20][47] = 9'b110010010;
assign micromatri[20][48] = 9'b111111111;
assign micromatri[20][49] = 9'b111111111;
assign micromatri[20][50] = 9'b111111111;
assign micromatri[20][51] = 9'b111111111;
assign micromatri[20][52] = 9'b110010110;
assign micromatri[20][53] = 9'b111111111;
assign micromatri[20][54] = 9'b111111111;
assign micromatri[20][55] = 9'b111111111;
assign micromatri[20][56] = 9'b111111111;
assign micromatri[20][57] = 9'b111111111;
assign micromatri[20][58] = 9'b111111111;
assign micromatri[20][59] = 9'b111111111;
assign micromatri[20][60] = 9'b110010001;
assign micromatri[20][61] = 9'b110110010;
assign micromatri[20][62] = 9'b111110011;
assign micromatri[20][63] = 9'b110110001;
assign micromatri[20][64] = 9'b110001101;
assign micromatri[20][65] = 9'b111111111;
assign micromatri[20][66] = 9'b110110110;
assign micromatri[20][67] = 9'b101101101;
assign micromatri[20][68] = 9'b111110111;
assign micromatri[20][69] = 9'b111110111;
assign micromatri[20][70] = 9'b111110111;
assign micromatri[20][71] = 9'b111110111;
assign micromatri[20][72] = 9'b111110111;
assign micromatri[20][73] = 9'b111110111;
assign micromatri[20][74] = 9'b111110111;
assign micromatri[20][75] = 9'b111110111;
assign micromatri[20][76] = 9'b111110111;
assign micromatri[20][77] = 9'b111110111;
assign micromatri[20][78] = 9'b111110111;
assign micromatri[20][79] = 9'b111110111;
assign micromatri[20][80] = 9'b111111111;
assign micromatri[20][81] = 9'b110001101;
assign micromatri[20][82] = 9'b110010010;
assign micromatri[20][83] = 9'b111111111;
assign micromatri[20][84] = 9'b111111111;
assign micromatri[20][85] = 9'b111111111;
assign micromatri[20][86] = 9'b111111111;
assign micromatri[20][87] = 9'b111111111;
assign micromatri[20][88] = 9'b111111111;
assign micromatri[20][89] = 9'b111111111;
assign micromatri[20][90] = 9'b111111111;
assign micromatri[20][91] = 9'b111111111;
assign micromatri[20][92] = 9'b111111111;
assign micromatri[20][93] = 9'b111111111;
assign micromatri[20][94] = 9'b111111111;
assign micromatri[20][95] = 9'b111111111;
assign micromatri[20][96] = 9'b111111111;
assign micromatri[20][97] = 9'b111111111;
assign micromatri[20][98] = 9'b111111111;
assign micromatri[20][99] = 9'b111111111;
assign micromatri[21][0] = 9'b111111111;
assign micromatri[21][1] = 9'b111111111;
assign micromatri[21][2] = 9'b111111111;
assign micromatri[21][3] = 9'b111111111;
assign micromatri[21][4] = 9'b111111111;
assign micromatri[21][5] = 9'b111111111;
assign micromatri[21][6] = 9'b111111111;
assign micromatri[21][7] = 9'b111111111;
assign micromatri[21][8] = 9'b111111111;
assign micromatri[21][9] = 9'b111111111;
assign micromatri[21][10] = 9'b111111111;
assign micromatri[21][11] = 9'b111111111;
assign micromatri[21][12] = 9'b111111111;
assign micromatri[21][13] = 9'b111111111;
assign micromatri[21][14] = 9'b111111111;
assign micromatri[21][15] = 9'b111111111;
assign micromatri[21][16] = 9'b111111111;
assign micromatri[21][17] = 9'b111111111;
assign micromatri[21][18] = 9'b111111111;
assign micromatri[21][19] = 9'b111111111;
assign micromatri[21][20] = 9'b111111111;
assign micromatri[21][21] = 9'b111111111;
assign micromatri[21][22] = 9'b111111111;
assign micromatri[21][23] = 9'b110010001;
assign micromatri[21][24] = 9'b111110111;
assign micromatri[21][25] = 9'b111110111;
assign micromatri[21][26] = 9'b111110111;
assign micromatri[21][27] = 9'b111110111;
assign micromatri[21][28] = 9'b111110111;
assign micromatri[21][29] = 9'b111110111;
assign micromatri[21][30] = 9'b110110010;
assign micromatri[21][31] = 9'b110010010;
assign micromatri[21][32] = 9'b111110011;
assign micromatri[21][33] = 9'b111110111;
assign micromatri[21][34] = 9'b111110111;
assign micromatri[21][35] = 9'b111110111;
assign micromatri[21][36] = 9'b111110111;
assign micromatri[21][37] = 9'b111110111;
assign micromatri[21][38] = 9'b110010010;
assign micromatri[21][39] = 9'b111111111;
assign micromatri[21][40] = 9'b111111111;
assign micromatri[21][41] = 9'b110110010;
assign micromatri[21][42] = 9'b111110011;
assign micromatri[21][43] = 9'b111110111;
assign micromatri[21][44] = 9'b111110111;
assign micromatri[21][45] = 9'b110001110;
assign micromatri[21][46] = 9'b111110111;
assign micromatri[21][47] = 9'b110010010;
assign micromatri[21][48] = 9'b111111111;
assign micromatri[21][49] = 9'b111111111;
assign micromatri[21][50] = 9'b111111111;
assign micromatri[21][51] = 9'b111111111;
assign micromatri[21][52] = 9'b110010110;
assign micromatri[21][53] = 9'b111111111;
assign micromatri[21][54] = 9'b111111111;
assign micromatri[21][55] = 9'b111111111;
assign micromatri[21][56] = 9'b111111111;
assign micromatri[21][57] = 9'b111111111;
assign micromatri[21][58] = 9'b111111111;
assign micromatri[21][59] = 9'b110110110;
assign micromatri[21][60] = 9'b110010001;
assign micromatri[21][61] = 9'b101101001;
assign micromatri[21][62] = 9'b101101001;
assign micromatri[21][63] = 9'b101101101;
assign micromatri[21][64] = 9'b110001101;
assign micromatri[21][65] = 9'b110110010;
assign micromatri[21][66] = 9'b110001101;
assign micromatri[21][67] = 9'b110110011;
assign micromatri[21][68] = 9'b111110111;
assign micromatri[21][69] = 9'b111110111;
assign micromatri[21][70] = 9'b111110111;
assign micromatri[21][71] = 9'b111110111;
assign micromatri[21][72] = 9'b111110111;
assign micromatri[21][73] = 9'b111110111;
assign micromatri[21][74] = 9'b111110111;
assign micromatri[21][75] = 9'b111110111;
assign micromatri[21][76] = 9'b111110111;
assign micromatri[21][77] = 9'b111110111;
assign micromatri[21][78] = 9'b111110111;
assign micromatri[21][79] = 9'b111110111;
assign micromatri[21][80] = 9'b111110111;
assign micromatri[21][81] = 9'b111110011;
assign micromatri[21][82] = 9'b110001101;
assign micromatri[21][83] = 9'b111111111;
assign micromatri[21][84] = 9'b111111111;
assign micromatri[21][85] = 9'b111111111;
assign micromatri[21][86] = 9'b111111111;
assign micromatri[21][87] = 9'b111111111;
assign micromatri[21][88] = 9'b111111111;
assign micromatri[21][89] = 9'b111111111;
assign micromatri[21][90] = 9'b111111111;
assign micromatri[21][91] = 9'b111111111;
assign micromatri[21][92] = 9'b111111111;
assign micromatri[21][93] = 9'b111111111;
assign micromatri[21][94] = 9'b111111111;
assign micromatri[21][95] = 9'b111111111;
assign micromatri[21][96] = 9'b111111111;
assign micromatri[21][97] = 9'b111111111;
assign micromatri[21][98] = 9'b111111111;
assign micromatri[21][99] = 9'b111111111;
assign micromatri[22][0] = 9'b111111111;
assign micromatri[22][1] = 9'b111111111;
assign micromatri[22][2] = 9'b111111111;
assign micromatri[22][3] = 9'b111111111;
assign micromatri[22][4] = 9'b111111111;
assign micromatri[22][5] = 9'b111111111;
assign micromatri[22][6] = 9'b111111111;
assign micromatri[22][7] = 9'b111111111;
assign micromatri[22][8] = 9'b111111111;
assign micromatri[22][9] = 9'b111111111;
assign micromatri[22][10] = 9'b111111111;
assign micromatri[22][11] = 9'b111111111;
assign micromatri[22][12] = 9'b111111111;
assign micromatri[22][13] = 9'b111111111;
assign micromatri[22][14] = 9'b111111111;
assign micromatri[22][15] = 9'b111111111;
assign micromatri[22][16] = 9'b111111111;
assign micromatri[22][17] = 9'b111111111;
assign micromatri[22][18] = 9'b111111111;
assign micromatri[22][19] = 9'b111111111;
assign micromatri[22][20] = 9'b111111111;
assign micromatri[22][21] = 9'b111111111;
assign micromatri[22][22] = 9'b111111111;
assign micromatri[22][23] = 9'b110110110;
assign micromatri[22][24] = 9'b111110010;
assign micromatri[22][25] = 9'b111110111;
assign micromatri[22][26] = 9'b111110111;
assign micromatri[22][27] = 9'b111110111;
assign micromatri[22][28] = 9'b111110111;
assign micromatri[22][29] = 9'b111110111;
assign micromatri[22][30] = 9'b110110010;
assign micromatri[22][31] = 9'b110010010;
assign micromatri[22][32] = 9'b111110011;
assign micromatri[22][33] = 9'b111110111;
assign micromatri[22][34] = 9'b111110111;
assign micromatri[22][35] = 9'b111110111;
assign micromatri[22][36] = 9'b111110111;
assign micromatri[22][37] = 9'b111110111;
assign micromatri[22][38] = 9'b110010010;
assign micromatri[22][39] = 9'b111111111;
assign micromatri[22][40] = 9'b111111111;
assign micromatri[22][41] = 9'b110010010;
assign micromatri[22][42] = 9'b111110011;
assign micromatri[22][43] = 9'b111110111;
assign micromatri[22][44] = 9'b111110111;
assign micromatri[22][45] = 9'b110001110;
assign micromatri[22][46] = 9'b111111111;
assign micromatri[22][47] = 9'b110010001;
assign micromatri[22][48] = 9'b111111111;
assign micromatri[22][49] = 9'b111111111;
assign micromatri[22][50] = 9'b111111111;
assign micromatri[22][51] = 9'b111111111;
assign micromatri[22][52] = 9'b110010110;
assign micromatri[22][53] = 9'b111111111;
assign micromatri[22][54] = 9'b111111111;
assign micromatri[22][55] = 9'b111111111;
assign micromatri[22][56] = 9'b111111111;
assign micromatri[22][57] = 9'b111111111;
assign micromatri[22][58] = 9'b111111111;
assign micromatri[22][59] = 9'b110010001;
assign micromatri[22][60] = 9'b111110111;
assign micromatri[22][61] = 9'b111111111;
assign micromatri[22][62] = 9'b111111111;
assign micromatri[22][63] = 9'b111111111;
assign micromatri[22][64] = 9'b111110111;
assign micromatri[22][65] = 9'b110001101;
assign micromatri[22][66] = 9'b110001101;
assign micromatri[22][67] = 9'b111110111;
assign micromatri[22][68] = 9'b111110111;
assign micromatri[22][69] = 9'b111110111;
assign micromatri[22][70] = 9'b111110111;
assign micromatri[22][71] = 9'b111110111;
assign micromatri[22][72] = 9'b111110111;
assign micromatri[22][73] = 9'b110001110;
assign micromatri[22][74] = 9'b110001101;
assign micromatri[22][75] = 9'b110001110;
assign micromatri[22][76] = 9'b111110111;
assign micromatri[22][77] = 9'b111110111;
assign micromatri[22][78] = 9'b111110111;
assign micromatri[22][79] = 9'b111110111;
assign micromatri[22][80] = 9'b111110111;
assign micromatri[22][81] = 9'b111110111;
assign micromatri[22][82] = 9'b110001110;
assign micromatri[22][83] = 9'b111111111;
assign micromatri[22][84] = 9'b111111111;
assign micromatri[22][85] = 9'b111111111;
assign micromatri[22][86] = 9'b111111111;
assign micromatri[22][87] = 9'b111111111;
assign micromatri[22][88] = 9'b111111111;
assign micromatri[22][89] = 9'b111111111;
assign micromatri[22][90] = 9'b111111111;
assign micromatri[22][91] = 9'b111111111;
assign micromatri[22][92] = 9'b111111111;
assign micromatri[22][93] = 9'b111111111;
assign micromatri[22][94] = 9'b111111111;
assign micromatri[22][95] = 9'b111111111;
assign micromatri[22][96] = 9'b111111111;
assign micromatri[22][97] = 9'b111111111;
assign micromatri[22][98] = 9'b111111111;
assign micromatri[22][99] = 9'b111111111;
assign micromatri[23][0] = 9'b111111111;
assign micromatri[23][1] = 9'b111111111;
assign micromatri[23][2] = 9'b111111111;
assign micromatri[23][3] = 9'b111111111;
assign micromatri[23][4] = 9'b111111111;
assign micromatri[23][5] = 9'b111111111;
assign micromatri[23][6] = 9'b111111111;
assign micromatri[23][7] = 9'b111111111;
assign micromatri[23][8] = 9'b111111111;
assign micromatri[23][9] = 9'b111111111;
assign micromatri[23][10] = 9'b111111111;
assign micromatri[23][11] = 9'b111111111;
assign micromatri[23][12] = 9'b111111111;
assign micromatri[23][13] = 9'b111111111;
assign micromatri[23][14] = 9'b111111111;
assign micromatri[23][15] = 9'b111111111;
assign micromatri[23][16] = 9'b111111111;
assign micromatri[23][17] = 9'b111111111;
assign micromatri[23][18] = 9'b111111111;
assign micromatri[23][19] = 9'b111111111;
assign micromatri[23][20] = 9'b111111111;
assign micromatri[23][21] = 9'b111111111;
assign micromatri[23][22] = 9'b111111111;
assign micromatri[23][23] = 9'b111111111;
assign micromatri[23][24] = 9'b111110010;
assign micromatri[23][25] = 9'b111111111;
assign micromatri[23][26] = 9'b111110111;
assign micromatri[23][27] = 9'b111110111;
assign micromatri[23][28] = 9'b111110111;
assign micromatri[23][29] = 9'b111110111;
assign micromatri[23][30] = 9'b110110010;
assign micromatri[23][31] = 9'b110110010;
assign micromatri[23][32] = 9'b111110011;
assign micromatri[23][33] = 9'b111110111;
assign micromatri[23][34] = 9'b111110111;
assign micromatri[23][35] = 9'b111110111;
assign micromatri[23][36] = 9'b111110111;
assign micromatri[23][37] = 9'b111110111;
assign micromatri[23][38] = 9'b110001110;
assign micromatri[23][39] = 9'b111110111;
assign micromatri[23][40] = 9'b111111111;
assign micromatri[23][41] = 9'b110010010;
assign micromatri[23][42] = 9'b111110111;
assign micromatri[23][43] = 9'b111110111;
assign micromatri[23][44] = 9'b111110111;
assign micromatri[23][45] = 9'b110001110;
assign micromatri[23][46] = 9'b111111111;
assign micromatri[23][47] = 9'b101110001;
assign micromatri[23][48] = 9'b111111111;
assign micromatri[23][49] = 9'b111111111;
assign micromatri[23][50] = 9'b111111111;
assign micromatri[23][51] = 9'b111111111;
assign micromatri[23][52] = 9'b110010110;
assign micromatri[23][53] = 9'b111111111;
assign micromatri[23][54] = 9'b111111111;
assign micromatri[23][55] = 9'b111111111;
assign micromatri[23][56] = 9'b111111111;
assign micromatri[23][57] = 9'b111111111;
assign micromatri[23][58] = 9'b111111111;
assign micromatri[23][59] = 9'b110010010;
assign micromatri[23][60] = 9'b111110111;
assign micromatri[23][61] = 9'b111110111;
assign micromatri[23][62] = 9'b111110111;
assign micromatri[23][63] = 9'b111110111;
assign micromatri[23][64] = 9'b111110111;
assign micromatri[23][65] = 9'b110010001;
assign micromatri[23][66] = 9'b110010010;
assign micromatri[23][67] = 9'b111110111;
assign micromatri[23][68] = 9'b111110111;
assign micromatri[23][69] = 9'b111110111;
assign micromatri[23][70] = 9'b111110111;
assign micromatri[23][71] = 9'b111110111;
assign micromatri[23][72] = 9'b110001110;
assign micromatri[23][73] = 9'b110110010;
assign micromatri[23][74] = 9'b111111111;
assign micromatri[23][75] = 9'b110010010;
assign micromatri[23][76] = 9'b110001101;
assign micromatri[23][77] = 9'b111110111;
assign micromatri[23][78] = 9'b111110111;
assign micromatri[23][79] = 9'b111110111;
assign micromatri[23][80] = 9'b111110111;
assign micromatri[23][81] = 9'b111110111;
assign micromatri[23][82] = 9'b110010010;
assign micromatri[23][83] = 9'b111110111;
assign micromatri[23][84] = 9'b111111111;
assign micromatri[23][85] = 9'b111111111;
assign micromatri[23][86] = 9'b111111111;
assign micromatri[23][87] = 9'b111111111;
assign micromatri[23][88] = 9'b111111111;
assign micromatri[23][89] = 9'b111111111;
assign micromatri[23][90] = 9'b111111111;
assign micromatri[23][91] = 9'b111111111;
assign micromatri[23][92] = 9'b111111111;
assign micromatri[23][93] = 9'b111111111;
assign micromatri[23][94] = 9'b111111111;
assign micromatri[23][95] = 9'b111111111;
assign micromatri[23][96] = 9'b111111111;
assign micromatri[23][97] = 9'b111111111;
assign micromatri[23][98] = 9'b111111111;
assign micromatri[23][99] = 9'b111111111;
assign micromatri[24][0] = 9'b111111111;
assign micromatri[24][1] = 9'b111111111;
assign micromatri[24][2] = 9'b111111111;
assign micromatri[24][3] = 9'b111111111;
assign micromatri[24][4] = 9'b111111111;
assign micromatri[24][5] = 9'b111111111;
assign micromatri[24][6] = 9'b111111111;
assign micromatri[24][7] = 9'b111111111;
assign micromatri[24][8] = 9'b111111111;
assign micromatri[24][9] = 9'b111111111;
assign micromatri[24][10] = 9'b111111111;
assign micromatri[24][11] = 9'b111111111;
assign micromatri[24][12] = 9'b111111111;
assign micromatri[24][13] = 9'b111111111;
assign micromatri[24][14] = 9'b111111111;
assign micromatri[24][15] = 9'b110110110;
assign micromatri[24][16] = 9'b110001101;
assign micromatri[24][17] = 9'b110110010;
assign micromatri[24][18] = 9'b110110010;
assign micromatri[24][19] = 9'b110110010;
assign micromatri[24][20] = 9'b110001101;
assign micromatri[24][21] = 9'b111111111;
assign micromatri[24][22] = 9'b111111111;
assign micromatri[24][23] = 9'b111111111;
assign micromatri[24][24] = 9'b111110010;
assign micromatri[24][25] = 9'b111111111;
assign micromatri[24][26] = 9'b111110111;
assign micromatri[24][27] = 9'b111110111;
assign micromatri[24][28] = 9'b111110111;
assign micromatri[24][29] = 9'b111110111;
assign micromatri[24][30] = 9'b110110010;
assign micromatri[24][31] = 9'b110110010;
assign micromatri[24][32] = 9'b110110011;
assign micromatri[24][33] = 9'b111110111;
assign micromatri[24][34] = 9'b111110111;
assign micromatri[24][35] = 9'b111110111;
assign micromatri[24][36] = 9'b111110111;
assign micromatri[24][37] = 9'b111110111;
assign micromatri[24][38] = 9'b110001110;
assign micromatri[24][39] = 9'b111110111;
assign micromatri[24][40] = 9'b111111111;
assign micromatri[24][41] = 9'b110010010;
assign micromatri[24][42] = 9'b111110111;
assign micromatri[24][43] = 9'b111110111;
assign micromatri[24][44] = 9'b111110111;
assign micromatri[24][45] = 9'b110010010;
assign micromatri[24][46] = 9'b111111111;
assign micromatri[24][47] = 9'b101110001;
assign micromatri[24][48] = 9'b111111111;
assign micromatri[24][49] = 9'b111111111;
assign micromatri[24][50] = 9'b111111111;
assign micromatri[24][51] = 9'b111111111;
assign micromatri[24][52] = 9'b110010110;
assign micromatri[24][53] = 9'b111111111;
assign micromatri[24][54] = 9'b111111111;
assign micromatri[24][55] = 9'b111111111;
assign micromatri[24][56] = 9'b111111111;
assign micromatri[24][57] = 9'b111111111;
assign micromatri[24][58] = 9'b111111111;
assign micromatri[24][59] = 9'b110010010;
assign micromatri[24][60] = 9'b111110111;
assign micromatri[24][61] = 9'b111110111;
assign micromatri[24][62] = 9'b111110111;
assign micromatri[24][63] = 9'b111110111;
assign micromatri[24][64] = 9'b111110111;
assign micromatri[24][65] = 9'b110010001;
assign micromatri[24][66] = 9'b110010010;
assign micromatri[24][67] = 9'b111110111;
assign micromatri[24][68] = 9'b111110111;
assign micromatri[24][69] = 9'b111110111;
assign micromatri[24][70] = 9'b111110111;
assign micromatri[24][71] = 9'b111110011;
assign micromatri[24][72] = 9'b110010010;
assign micromatri[24][73] = 9'b111111111;
assign micromatri[24][74] = 9'b111110111;
assign micromatri[24][75] = 9'b111111111;
assign micromatri[24][76] = 9'b110010001;
assign micromatri[24][77] = 9'b111110011;
assign micromatri[24][78] = 9'b111110111;
assign micromatri[24][79] = 9'b111110111;
assign micromatri[24][80] = 9'b111110111;
assign micromatri[24][81] = 9'b111110111;
assign micromatri[24][82] = 9'b110010010;
assign micromatri[24][83] = 9'b111111111;
assign micromatri[24][84] = 9'b111111111;
assign micromatri[24][85] = 9'b111111111;
assign micromatri[24][86] = 9'b111111111;
assign micromatri[24][87] = 9'b111111111;
assign micromatri[24][88] = 9'b111111111;
assign micromatri[24][89] = 9'b111111111;
assign micromatri[24][90] = 9'b111111111;
assign micromatri[24][91] = 9'b111111111;
assign micromatri[24][92] = 9'b111111111;
assign micromatri[24][93] = 9'b111111111;
assign micromatri[24][94] = 9'b111111111;
assign micromatri[24][95] = 9'b111111111;
assign micromatri[24][96] = 9'b111111111;
assign micromatri[24][97] = 9'b111111111;
assign micromatri[24][98] = 9'b111111111;
assign micromatri[24][99] = 9'b111111111;
assign micromatri[25][0] = 9'b111111111;
assign micromatri[25][1] = 9'b111111111;
assign micromatri[25][2] = 9'b111111111;
assign micromatri[25][3] = 9'b111111111;
assign micromatri[25][4] = 9'b111111111;
assign micromatri[25][5] = 9'b111111111;
assign micromatri[25][6] = 9'b111111111;
assign micromatri[25][7] = 9'b111111111;
assign micromatri[25][8] = 9'b111111111;
assign micromatri[25][9] = 9'b111111111;
assign micromatri[25][10] = 9'b111111111;
assign micromatri[25][11] = 9'b111111111;
assign micromatri[25][12] = 9'b111111111;
assign micromatri[25][13] = 9'b111111111;
assign micromatri[25][14] = 9'b111111111;
assign micromatri[25][15] = 9'b110110110;
assign micromatri[25][16] = 9'b111110011;
assign micromatri[25][17] = 9'b111111111;
assign micromatri[25][18] = 9'b111111111;
assign micromatri[25][19] = 9'b111111111;
assign micromatri[25][20] = 9'b110110010;
assign micromatri[25][21] = 9'b110010001;
assign micromatri[25][22] = 9'b111111111;
assign micromatri[25][23] = 9'b110010010;
assign micromatri[25][24] = 9'b111110011;
assign micromatri[25][25] = 9'b111110111;
assign micromatri[25][26] = 9'b111110111;
assign micromatri[25][27] = 9'b111110111;
assign micromatri[25][28] = 9'b111110111;
assign micromatri[25][29] = 9'b111110011;
assign micromatri[25][30] = 9'b110110010;
assign micromatri[25][31] = 9'b111110111;
assign micromatri[25][32] = 9'b110001110;
assign micromatri[25][33] = 9'b111110111;
assign micromatri[25][34] = 9'b111110111;
assign micromatri[25][35] = 9'b111110111;
assign micromatri[25][36] = 9'b111110111;
assign micromatri[25][37] = 9'b111110111;
assign micromatri[25][38] = 9'b110110011;
assign micromatri[25][39] = 9'b110010001;
assign micromatri[25][40] = 9'b101101101;
assign micromatri[25][41] = 9'b110110011;
assign micromatri[25][42] = 9'b111110111;
assign micromatri[25][43] = 9'b111110111;
assign micromatri[25][44] = 9'b111110011;
assign micromatri[25][45] = 9'b110010010;
assign micromatri[25][46] = 9'b111111111;
assign micromatri[25][47] = 9'b101110001;
assign micromatri[25][48] = 9'b111111111;
assign micromatri[25][49] = 9'b111111111;
assign micromatri[25][50] = 9'b111111111;
assign micromatri[25][51] = 9'b111111111;
assign micromatri[25][52] = 9'b110010010;
assign micromatri[25][53] = 9'b110010010;
assign micromatri[25][54] = 9'b110010010;
assign micromatri[25][55] = 9'b110010010;
assign micromatri[25][56] = 9'b110010110;
assign micromatri[25][57] = 9'b110010001;
assign micromatri[25][58] = 9'b111111111;
assign micromatri[25][59] = 9'b110110010;
assign micromatri[25][60] = 9'b111110111;
assign micromatri[25][61] = 9'b111110111;
assign micromatri[25][62] = 9'b111110111;
assign micromatri[25][63] = 9'b111110111;
assign micromatri[25][64] = 9'b111110111;
assign micromatri[25][65] = 9'b110010001;
assign micromatri[25][66] = 9'b110010010;
assign micromatri[25][67] = 9'b111110111;
assign micromatri[25][68] = 9'b111110111;
assign micromatri[25][69] = 9'b111110111;
assign micromatri[25][70] = 9'b111110111;
assign micromatri[25][71] = 9'b111110011;
assign micromatri[25][72] = 9'b110010010;
assign micromatri[25][73] = 9'b111111111;
assign micromatri[25][74] = 9'b111111111;
assign micromatri[25][75] = 9'b111111111;
assign micromatri[25][76] = 9'b110110010;
assign micromatri[25][77] = 9'b111110011;
assign micromatri[25][78] = 9'b111110111;
assign micromatri[25][79] = 9'b111110111;
assign micromatri[25][80] = 9'b111110111;
assign micromatri[25][81] = 9'b111110111;
assign micromatri[25][82] = 9'b110001110;
assign micromatri[25][83] = 9'b111111111;
assign micromatri[25][84] = 9'b111111111;
assign micromatri[25][85] = 9'b111111111;
assign micromatri[25][86] = 9'b111111111;
assign micromatri[25][87] = 9'b111111111;
assign micromatri[25][88] = 9'b111111111;
assign micromatri[25][89] = 9'b111111111;
assign micromatri[25][90] = 9'b111111111;
assign micromatri[25][91] = 9'b111111111;
assign micromatri[25][92] = 9'b111111111;
assign micromatri[25][93] = 9'b111111111;
assign micromatri[25][94] = 9'b111111111;
assign micromatri[25][95] = 9'b111111111;
assign micromatri[25][96] = 9'b111111111;
assign micromatri[25][97] = 9'b111111111;
assign micromatri[25][98] = 9'b111111111;
assign micromatri[25][99] = 9'b111111111;
assign micromatri[26][0] = 9'b111111111;
assign micromatri[26][1] = 9'b111111111;
assign micromatri[26][2] = 9'b111111111;
assign micromatri[26][3] = 9'b111111111;
assign micromatri[26][4] = 9'b111111111;
assign micromatri[26][5] = 9'b111111111;
assign micromatri[26][6] = 9'b111111111;
assign micromatri[26][7] = 9'b111111111;
assign micromatri[26][8] = 9'b111111111;
assign micromatri[26][9] = 9'b111111111;
assign micromatri[26][10] = 9'b111111111;
assign micromatri[26][11] = 9'b111111111;
assign micromatri[26][12] = 9'b111111111;
assign micromatri[26][13] = 9'b111111111;
assign micromatri[26][14] = 9'b111111111;
assign micromatri[26][15] = 9'b110110110;
assign micromatri[26][16] = 9'b111110010;
assign micromatri[26][17] = 9'b111111111;
assign micromatri[26][18] = 9'b111110111;
assign micromatri[26][19] = 9'b111110111;
assign micromatri[26][20] = 9'b111110111;
assign micromatri[26][21] = 9'b110001101;
assign micromatri[26][22] = 9'b110001101;
assign micromatri[26][23] = 9'b110110010;
assign micromatri[26][24] = 9'b111111111;
assign micromatri[26][25] = 9'b111110111;
assign micromatri[26][26] = 9'b111110111;
assign micromatri[26][27] = 9'b111110111;
assign micromatri[26][28] = 9'b111111111;
assign micromatri[26][29] = 9'b111110010;
assign micromatri[26][30] = 9'b111110010;
assign micromatri[26][31] = 9'b111111111;
assign micromatri[26][32] = 9'b101101101;
assign micromatri[26][33] = 9'b111110111;
assign micromatri[26][34] = 9'b111110111;
assign micromatri[26][35] = 9'b111110111;
assign micromatri[26][36] = 9'b111110111;
assign micromatri[26][37] = 9'b111110111;
assign micromatri[26][38] = 9'b111110111;
assign micromatri[26][39] = 9'b110010010;
assign micromatri[26][40] = 9'b110110011;
assign micromatri[26][41] = 9'b111110111;
assign micromatri[26][42] = 9'b111110111;
assign micromatri[26][43] = 9'b111110111;
assign micromatri[26][44] = 9'b110110011;
assign micromatri[26][45] = 9'b110110010;
assign micromatri[26][46] = 9'b111111111;
assign micromatri[26][47] = 9'b110010001;
assign micromatri[26][48] = 9'b111111111;
assign micromatri[26][49] = 9'b111111111;
assign micromatri[26][50] = 9'b111111111;
assign micromatri[26][51] = 9'b111111111;
assign micromatri[26][52] = 9'b111111111;
assign micromatri[26][53] = 9'b111111111;
assign micromatri[26][54] = 9'b111111111;
assign micromatri[26][55] = 9'b111111111;
assign micromatri[26][56] = 9'b111111111;
assign micromatri[26][57] = 9'b110011111;
assign micromatri[26][58] = 9'b110010010;
assign micromatri[26][59] = 9'b110110010;
assign micromatri[26][60] = 9'b111110111;
assign micromatri[26][61] = 9'b111110111;
assign micromatri[26][62] = 9'b111110111;
assign micromatri[26][63] = 9'b111110111;
assign micromatri[26][64] = 9'b111110111;
assign micromatri[26][65] = 9'b110110010;
assign micromatri[26][66] = 9'b110010010;
assign micromatri[26][67] = 9'b111110011;
assign micromatri[26][68] = 9'b111110111;
assign micromatri[26][69] = 9'b111110111;
assign micromatri[26][70] = 9'b111110111;
assign micromatri[26][71] = 9'b111110111;
assign micromatri[26][72] = 9'b110001101;
assign micromatri[26][73] = 9'b110110110;
assign micromatri[26][74] = 9'b111111111;
assign micromatri[26][75] = 9'b111111111;
assign micromatri[26][76] = 9'b110001101;
assign micromatri[26][77] = 9'b111110111;
assign micromatri[26][78] = 9'b111110111;
assign micromatri[26][79] = 9'b111110111;
assign micromatri[26][80] = 9'b111110111;
assign micromatri[26][81] = 9'b111110011;
assign micromatri[26][82] = 9'b110010010;
assign micromatri[26][83] = 9'b111111111;
assign micromatri[26][84] = 9'b111111111;
assign micromatri[26][85] = 9'b111111111;
assign micromatri[26][86] = 9'b111111111;
assign micromatri[26][87] = 9'b111111111;
assign micromatri[26][88] = 9'b111111111;
assign micromatri[26][89] = 9'b111111111;
assign micromatri[26][90] = 9'b111111111;
assign micromatri[26][91] = 9'b111111111;
assign micromatri[26][92] = 9'b111111111;
assign micromatri[26][93] = 9'b111111111;
assign micromatri[26][94] = 9'b111111111;
assign micromatri[26][95] = 9'b111111111;
assign micromatri[26][96] = 9'b111111111;
assign micromatri[26][97] = 9'b111111111;
assign micromatri[26][98] = 9'b111111111;
assign micromatri[26][99] = 9'b111111111;
assign micromatri[27][0] = 9'b111111111;
assign micromatri[27][1] = 9'b111111111;
assign micromatri[27][2] = 9'b111111111;
assign micromatri[27][3] = 9'b111111111;
assign micromatri[27][4] = 9'b111111111;
assign micromatri[27][5] = 9'b111111111;
assign micromatri[27][6] = 9'b111111111;
assign micromatri[27][7] = 9'b111111111;
assign micromatri[27][8] = 9'b111111111;
assign micromatri[27][9] = 9'b111111111;
assign micromatri[27][10] = 9'b111111111;
assign micromatri[27][11] = 9'b111111111;
assign micromatri[27][12] = 9'b111111111;
assign micromatri[27][13] = 9'b111111111;
assign micromatri[27][14] = 9'b111111111;
assign micromatri[27][15] = 9'b111111111;
assign micromatri[27][16] = 9'b110110010;
assign micromatri[27][17] = 9'b111111111;
assign micromatri[27][18] = 9'b111110111;
assign micromatri[27][19] = 9'b111110111;
assign micromatri[27][20] = 9'b111110111;
assign micromatri[27][21] = 9'b111110111;
assign micromatri[27][22] = 9'b111110111;
assign micromatri[27][23] = 9'b111110111;
assign micromatri[27][24] = 9'b111110111;
assign micromatri[27][25] = 9'b111110111;
assign micromatri[27][26] = 9'b111110111;
assign micromatri[27][27] = 9'b111110111;
assign micromatri[27][28] = 9'b111111111;
assign micromatri[27][29] = 9'b110001101;
assign micromatri[27][30] = 9'b111111111;
assign micromatri[27][31] = 9'b111111111;
assign micromatri[27][32] = 9'b110010001;
assign micromatri[27][33] = 9'b111110011;
assign micromatri[27][34] = 9'b111110111;
assign micromatri[27][35] = 9'b111110111;
assign micromatri[27][36] = 9'b111110111;
assign micromatri[27][37] = 9'b111110111;
assign micromatri[27][38] = 9'b111110111;
assign micromatri[27][39] = 9'b111110111;
assign micromatri[27][40] = 9'b111110111;
assign micromatri[27][41] = 9'b111110111;
assign micromatri[27][42] = 9'b111110111;
assign micromatri[27][43] = 9'b111110111;
assign micromatri[27][44] = 9'b110001110;
assign micromatri[27][45] = 9'b111110111;
assign micromatri[27][46] = 9'b111111111;
assign micromatri[27][47] = 9'b110010001;
assign micromatri[27][48] = 9'b111111111;
assign micromatri[27][49] = 9'b111111111;
assign micromatri[27][50] = 9'b111111111;
assign micromatri[27][51] = 9'b111111111;
assign micromatri[27][52] = 9'b111111111;
assign micromatri[27][53] = 9'b111111111;
assign micromatri[27][54] = 9'b111111111;
assign micromatri[27][55] = 9'b111111111;
assign micromatri[27][56] = 9'b111111111;
assign micromatri[27][57] = 9'b110111111;
assign micromatri[27][58] = 9'b110010010;
assign micromatri[27][59] = 9'b110010010;
assign micromatri[27][60] = 9'b111110111;
assign micromatri[27][61] = 9'b111110111;
assign micromatri[27][62] = 9'b111110111;
assign micromatri[27][63] = 9'b111110111;
assign micromatri[27][64] = 9'b111110111;
assign micromatri[27][65] = 9'b110110010;
assign micromatri[27][66] = 9'b110110010;
assign micromatri[27][67] = 9'b110001110;
assign micromatri[27][68] = 9'b111110111;
assign micromatri[27][69] = 9'b111110111;
assign micromatri[27][70] = 9'b111110111;
assign micromatri[27][71] = 9'b111110111;
assign micromatri[27][72] = 9'b111110011;
assign micromatri[27][73] = 9'b101101101;
assign micromatri[27][74] = 9'b110010010;
assign micromatri[27][75] = 9'b110001101;
assign micromatri[27][76] = 9'b111110011;
assign micromatri[27][77] = 9'b111110111;
assign micromatri[27][78] = 9'b111110111;
assign micromatri[27][79] = 9'b111110111;
assign micromatri[27][80] = 9'b111110111;
assign micromatri[27][81] = 9'b110001110;
assign micromatri[27][82] = 9'b110110011;
assign micromatri[27][83] = 9'b111111111;
assign micromatri[27][84] = 9'b111111111;
assign micromatri[27][85] = 9'b111111111;
assign micromatri[27][86] = 9'b111111111;
assign micromatri[27][87] = 9'b111111111;
assign micromatri[27][88] = 9'b111111111;
assign micromatri[27][89] = 9'b111111111;
assign micromatri[27][90] = 9'b111111111;
assign micromatri[27][91] = 9'b111111111;
assign micromatri[27][92] = 9'b111111111;
assign micromatri[27][93] = 9'b111111111;
assign micromatri[27][94] = 9'b111111111;
assign micromatri[27][95] = 9'b111111111;
assign micromatri[27][96] = 9'b111111111;
assign micromatri[27][97] = 9'b111111111;
assign micromatri[27][98] = 9'b111111111;
assign micromatri[27][99] = 9'b111111111;
assign micromatri[28][0] = 9'b111111111;
assign micromatri[28][1] = 9'b111111111;
assign micromatri[28][2] = 9'b111111111;
assign micromatri[28][3] = 9'b111111111;
assign micromatri[28][4] = 9'b111111111;
assign micromatri[28][5] = 9'b111111111;
assign micromatri[28][6] = 9'b111111111;
assign micromatri[28][7] = 9'b111111111;
assign micromatri[28][8] = 9'b111111111;
assign micromatri[28][9] = 9'b111111111;
assign micromatri[28][10] = 9'b111111111;
assign micromatri[28][11] = 9'b111111111;
assign micromatri[28][12] = 9'b111111111;
assign micromatri[28][13] = 9'b111111111;
assign micromatri[28][14] = 9'b111111111;
assign micromatri[28][15] = 9'b111111111;
assign micromatri[28][16] = 9'b110001101;
assign micromatri[28][17] = 9'b111110111;
assign micromatri[28][18] = 9'b111110111;
assign micromatri[28][19] = 9'b111110111;
assign micromatri[28][20] = 9'b111110111;
assign micromatri[28][21] = 9'b111110111;
assign micromatri[28][22] = 9'b111110111;
assign micromatri[28][23] = 9'b111110111;
assign micromatri[28][24] = 9'b111110111;
assign micromatri[28][25] = 9'b111110111;
assign micromatri[28][26] = 9'b111110111;
assign micromatri[28][27] = 9'b111111111;
assign micromatri[28][28] = 9'b111110011;
assign micromatri[28][29] = 9'b110010001;
assign micromatri[28][30] = 9'b111111111;
assign micromatri[28][31] = 9'b111111111;
assign micromatri[28][32] = 9'b111111111;
assign micromatri[28][33] = 9'b110001110;
assign micromatri[28][34] = 9'b111110111;
assign micromatri[28][35] = 9'b111110111;
assign micromatri[28][36] = 9'b111110111;
assign micromatri[28][37] = 9'b111110111;
assign micromatri[28][38] = 9'b111110111;
assign micromatri[28][39] = 9'b111110111;
assign micromatri[28][40] = 9'b111110111;
assign micromatri[28][41] = 9'b111110111;
assign micromatri[28][42] = 9'b111110111;
assign micromatri[28][43] = 9'b111110111;
assign micromatri[28][44] = 9'b110001101;
assign micromatri[28][45] = 9'b111111111;
assign micromatri[28][46] = 9'b111111111;
assign micromatri[28][47] = 9'b110010110;
assign micromatri[28][48] = 9'b111111111;
assign micromatri[28][49] = 9'b111111111;
assign micromatri[28][50] = 9'b111111111;
assign micromatri[28][51] = 9'b111111111;
assign micromatri[28][52] = 9'b111111111;
assign micromatri[28][53] = 9'b111111111;
assign micromatri[28][54] = 9'b111111111;
assign micromatri[28][55] = 9'b111111111;
assign micromatri[28][56] = 9'b111111111;
assign micromatri[28][57] = 9'b110111111;
assign micromatri[28][58] = 9'b110111111;
assign micromatri[28][59] = 9'b110110010;
assign micromatri[28][60] = 9'b111110111;
assign micromatri[28][61] = 9'b111110111;
assign micromatri[28][62] = 9'b111110111;
assign micromatri[28][63] = 9'b111110111;
assign micromatri[28][64] = 9'b111110111;
assign micromatri[28][65] = 9'b110110010;
assign micromatri[28][66] = 9'b111111111;
assign micromatri[28][67] = 9'b101101101;
assign micromatri[28][68] = 9'b111110111;
assign micromatri[28][69] = 9'b111110111;
assign micromatri[28][70] = 9'b111110111;
assign micromatri[28][71] = 9'b111110111;
assign micromatri[28][72] = 9'b111110111;
assign micromatri[28][73] = 9'b111110111;
assign micromatri[28][74] = 9'b111110011;
assign micromatri[28][75] = 9'b111110111;
assign micromatri[28][76] = 9'b111110111;
assign micromatri[28][77] = 9'b111110111;
assign micromatri[28][78] = 9'b111110111;
assign micromatri[28][79] = 9'b111110111;
assign micromatri[28][80] = 9'b111110011;
assign micromatri[28][81] = 9'b110001101;
assign micromatri[28][82] = 9'b111111111;
assign micromatri[28][83] = 9'b111110111;
assign micromatri[28][84] = 9'b111111111;
assign micromatri[28][85] = 9'b111111111;
assign micromatri[28][86] = 9'b111111111;
assign micromatri[28][87] = 9'b111111111;
assign micromatri[28][88] = 9'b111111111;
assign micromatri[28][89] = 9'b111111111;
assign micromatri[28][90] = 9'b111111111;
assign micromatri[28][91] = 9'b111111111;
assign micromatri[28][92] = 9'b111111111;
assign micromatri[28][93] = 9'b111111111;
assign micromatri[28][94] = 9'b111111111;
assign micromatri[28][95] = 9'b111111111;
assign micromatri[28][96] = 9'b111111111;
assign micromatri[28][97] = 9'b111111111;
assign micromatri[28][98] = 9'b111111111;
assign micromatri[28][99] = 9'b111111111;
assign micromatri[29][0] = 9'b111111111;
assign micromatri[29][1] = 9'b111111111;
assign micromatri[29][2] = 9'b111111111;
assign micromatri[29][3] = 9'b111111111;
assign micromatri[29][4] = 9'b111111111;
assign micromatri[29][5] = 9'b111111111;
assign micromatri[29][6] = 9'b111111111;
assign micromatri[29][7] = 9'b111111111;
assign micromatri[29][8] = 9'b111111111;
assign micromatri[29][9] = 9'b111111111;
assign micromatri[29][10] = 9'b111111111;
assign micromatri[29][11] = 9'b111111111;
assign micromatri[29][12] = 9'b111111111;
assign micromatri[29][13] = 9'b111111111;
assign micromatri[29][14] = 9'b111111111;
assign micromatri[29][15] = 9'b111111111;
assign micromatri[29][16] = 9'b110110110;
assign micromatri[29][17] = 9'b110110010;
assign micromatri[29][18] = 9'b111111111;
assign micromatri[29][19] = 9'b111110111;
assign micromatri[29][20] = 9'b111110111;
assign micromatri[29][21] = 9'b111110111;
assign micromatri[29][22] = 9'b111110111;
assign micromatri[29][23] = 9'b111110111;
assign micromatri[29][24] = 9'b111110111;
assign micromatri[29][25] = 9'b111110111;
assign micromatri[29][26] = 9'b111110111;
assign micromatri[29][27] = 9'b111111111;
assign micromatri[29][28] = 9'b110001101;
assign micromatri[29][29] = 9'b111111111;
assign micromatri[29][30] = 9'b111111111;
assign micromatri[29][31] = 9'b111111111;
assign micromatri[29][32] = 9'b111111111;
assign micromatri[29][33] = 9'b110001101;
assign micromatri[29][34] = 9'b111110011;
assign micromatri[29][35] = 9'b111110111;
assign micromatri[29][36] = 9'b111110111;
assign micromatri[29][37] = 9'b111110111;
assign micromatri[29][38] = 9'b111110111;
assign micromatri[29][39] = 9'b111110111;
assign micromatri[29][40] = 9'b111110111;
assign micromatri[29][41] = 9'b111110111;
assign micromatri[29][42] = 9'b111110111;
assign micromatri[29][43] = 9'b110001110;
assign micromatri[29][44] = 9'b110110010;
assign micromatri[29][45] = 9'b111111111;
assign micromatri[29][46] = 9'b111111111;
assign micromatri[29][47] = 9'b110110110;
assign micromatri[29][48] = 9'b111111111;
assign micromatri[29][49] = 9'b111111111;
assign micromatri[29][50] = 9'b111111111;
assign micromatri[29][51] = 9'b111111111;
assign micromatri[29][52] = 9'b111111111;
assign micromatri[29][53] = 9'b111111111;
assign micromatri[29][54] = 9'b111111111;
assign micromatri[29][55] = 9'b111111111;
assign micromatri[29][56] = 9'b111111111;
assign micromatri[29][57] = 9'b110111111;
assign micromatri[29][58] = 9'b110111111;
assign micromatri[29][59] = 9'b110110010;
assign micromatri[29][60] = 9'b111110111;
assign micromatri[29][61] = 9'b111110111;
assign micromatri[29][62] = 9'b111110111;
assign micromatri[29][63] = 9'b111110111;
assign micromatri[29][64] = 9'b111110111;
assign micromatri[29][65] = 9'b110110010;
assign micromatri[29][66] = 9'b111111111;
assign micromatri[29][67] = 9'b110110110;
assign micromatri[29][68] = 9'b110001110;
assign micromatri[29][69] = 9'b111110111;
assign micromatri[29][70] = 9'b111110111;
assign micromatri[29][71] = 9'b111110111;
assign micromatri[29][72] = 9'b111110111;
assign micromatri[29][73] = 9'b111110111;
assign micromatri[29][74] = 9'b111110111;
assign micromatri[29][75] = 9'b111110111;
assign micromatri[29][76] = 9'b111110111;
assign micromatri[29][77] = 9'b111110111;
assign micromatri[29][78] = 9'b111110111;
assign micromatri[29][79] = 9'b111110111;
assign micromatri[29][80] = 9'b110001101;
assign micromatri[29][81] = 9'b111110111;
assign micromatri[29][82] = 9'b111111111;
assign micromatri[29][83] = 9'b111111111;
assign micromatri[29][84] = 9'b111111111;
assign micromatri[29][85] = 9'b111111111;
assign micromatri[29][86] = 9'b111111111;
assign micromatri[29][87] = 9'b111111111;
assign micromatri[29][88] = 9'b111111111;
assign micromatri[29][89] = 9'b111111111;
assign micromatri[29][90] = 9'b111111111;
assign micromatri[29][91] = 9'b111111111;
assign micromatri[29][92] = 9'b111111111;
assign micromatri[29][93] = 9'b111111111;
assign micromatri[29][94] = 9'b111111111;
assign micromatri[29][95] = 9'b111111111;
assign micromatri[29][96] = 9'b111111111;
assign micromatri[29][97] = 9'b111111111;
assign micromatri[29][98] = 9'b111111111;
assign micromatri[29][99] = 9'b111111111;
assign micromatri[30][0] = 9'b111111111;
assign micromatri[30][1] = 9'b111111111;
assign micromatri[30][2] = 9'b111111111;
assign micromatri[30][3] = 9'b111111111;
assign micromatri[30][4] = 9'b111111111;
assign micromatri[30][5] = 9'b111111111;
assign micromatri[30][6] = 9'b111111111;
assign micromatri[30][7] = 9'b111111111;
assign micromatri[30][8] = 9'b111111111;
assign micromatri[30][9] = 9'b111111111;
assign micromatri[30][10] = 9'b111111111;
assign micromatri[30][11] = 9'b111111111;
assign micromatri[30][12] = 9'b111111111;
assign micromatri[30][13] = 9'b111111111;
assign micromatri[30][14] = 9'b111111111;
assign micromatri[30][15] = 9'b111111111;
assign micromatri[30][16] = 9'b111111111;
assign micromatri[30][17] = 9'b110010001;
assign micromatri[30][18] = 9'b111110010;
assign micromatri[30][19] = 9'b111111111;
assign micromatri[30][20] = 9'b111110111;
assign micromatri[30][21] = 9'b111110111;
assign micromatri[30][22] = 9'b111110111;
assign micromatri[30][23] = 9'b111110111;
assign micromatri[30][24] = 9'b111110111;
assign micromatri[30][25] = 9'b111111111;
assign micromatri[30][26] = 9'b111111111;
assign micromatri[30][27] = 9'b110001101;
assign micromatri[30][28] = 9'b110110010;
assign micromatri[30][29] = 9'b111111111;
assign micromatri[30][30] = 9'b111110111;
assign micromatri[30][31] = 9'b111111111;
assign micromatri[30][32] = 9'b111111111;
assign micromatri[30][33] = 9'b111111111;
assign micromatri[30][34] = 9'b110001101;
assign micromatri[30][35] = 9'b111110111;
assign micromatri[30][36] = 9'b111110111;
assign micromatri[30][37] = 9'b111110111;
assign micromatri[30][38] = 9'b111110111;
assign micromatri[30][39] = 9'b111110111;
assign micromatri[30][40] = 9'b111110111;
assign micromatri[30][41] = 9'b111110111;
assign micromatri[30][42] = 9'b111110011;
assign micromatri[30][43] = 9'b110001101;
assign micromatri[30][44] = 9'b111111111;
assign micromatri[30][45] = 9'b111110111;
assign micromatri[30][46] = 9'b111111111;
assign micromatri[30][47] = 9'b110110110;
assign micromatri[30][48] = 9'b111111111;
assign micromatri[30][49] = 9'b111111111;
assign micromatri[30][50] = 9'b111111111;
assign micromatri[30][51] = 9'b111111111;
assign micromatri[30][52] = 9'b111111111;
assign micromatri[30][53] = 9'b111111111;
assign micromatri[30][54] = 9'b111111111;
assign micromatri[30][55] = 9'b111111111;
assign micromatri[30][56] = 9'b111111111;
assign micromatri[30][57] = 9'b110111111;
assign micromatri[30][58] = 9'b110111111;
assign micromatri[30][59] = 9'b110110010;
assign micromatri[30][60] = 9'b111110111;
assign micromatri[30][61] = 9'b111110111;
assign micromatri[30][62] = 9'b111110111;
assign micromatri[30][63] = 9'b111110111;
assign micromatri[30][64] = 9'b111110111;
assign micromatri[30][65] = 9'b110110010;
assign micromatri[30][66] = 9'b111111111;
assign micromatri[30][67] = 9'b111111111;
assign micromatri[30][68] = 9'b110110110;
assign micromatri[30][69] = 9'b110001110;
assign micromatri[30][70] = 9'b111110111;
assign micromatri[30][71] = 9'b111110111;
assign micromatri[30][72] = 9'b111110111;
assign micromatri[30][73] = 9'b111110111;
assign micromatri[30][74] = 9'b111110111;
assign micromatri[30][75] = 9'b111110111;
assign micromatri[30][76] = 9'b111110111;
assign micromatri[30][77] = 9'b111110111;
assign micromatri[30][78] = 9'b111110111;
assign micromatri[30][79] = 9'b110001101;
assign micromatri[30][80] = 9'b110110111;
assign micromatri[30][81] = 9'b111111111;
assign micromatri[30][82] = 9'b111110111;
assign micromatri[30][83] = 9'b111111111;
assign micromatri[30][84] = 9'b111111111;
assign micromatri[30][85] = 9'b111111111;
assign micromatri[30][86] = 9'b111111111;
assign micromatri[30][87] = 9'b111111111;
assign micromatri[30][88] = 9'b111111111;
assign micromatri[30][89] = 9'b111111111;
assign micromatri[30][90] = 9'b111111111;
assign micromatri[30][91] = 9'b111111111;
assign micromatri[30][92] = 9'b111111111;
assign micromatri[30][93] = 9'b111111111;
assign micromatri[30][94] = 9'b111111111;
assign micromatri[30][95] = 9'b111111111;
assign micromatri[30][96] = 9'b111111111;
assign micromatri[30][97] = 9'b111111111;
assign micromatri[30][98] = 9'b111111111;
assign micromatri[30][99] = 9'b111111111;
assign micromatri[31][0] = 9'b111111111;
assign micromatri[31][1] = 9'b111111111;
assign micromatri[31][2] = 9'b111111111;
assign micromatri[31][3] = 9'b111111111;
assign micromatri[31][4] = 9'b111111111;
assign micromatri[31][5] = 9'b111111111;
assign micromatri[31][6] = 9'b111111111;
assign micromatri[31][7] = 9'b111111111;
assign micromatri[31][8] = 9'b111111111;
assign micromatri[31][9] = 9'b111111111;
assign micromatri[31][10] = 9'b111111111;
assign micromatri[31][11] = 9'b111111111;
assign micromatri[31][12] = 9'b111111111;
assign micromatri[31][13] = 9'b111111111;
assign micromatri[31][14] = 9'b111111111;
assign micromatri[31][15] = 9'b111111111;
assign micromatri[31][16] = 9'b111111111;
assign micromatri[31][17] = 9'b111111111;
assign micromatri[31][18] = 9'b110010001;
assign micromatri[31][19] = 9'b110001101;
assign micromatri[31][20] = 9'b111110111;
assign micromatri[31][21] = 9'b111110111;
assign micromatri[31][22] = 9'b111110111;
assign micromatri[31][23] = 9'b111110111;
assign micromatri[31][24] = 9'b111110111;
assign micromatri[31][25] = 9'b111110010;
assign micromatri[31][26] = 9'b110001101;
assign micromatri[31][27] = 9'b110110010;
assign micromatri[31][28] = 9'b111111111;
assign micromatri[31][29] = 9'b111110111;
assign micromatri[31][30] = 9'b111111111;
assign micromatri[31][31] = 9'b111111111;
assign micromatri[31][32] = 9'b111111111;
assign micromatri[31][33] = 9'b111111111;
assign micromatri[31][34] = 9'b110110110;
assign micromatri[31][35] = 9'b110001101;
assign micromatri[31][36] = 9'b111110111;
assign micromatri[31][37] = 9'b111110111;
assign micromatri[31][38] = 9'b111110111;
assign micromatri[31][39] = 9'b111110111;
assign micromatri[31][40] = 9'b111110111;
assign micromatri[31][41] = 9'b110110011;
assign micromatri[31][42] = 9'b101101101;
assign micromatri[31][43] = 9'b111111111;
assign micromatri[31][44] = 9'b111111111;
assign micromatri[31][45] = 9'b111111111;
assign micromatri[31][46] = 9'b111111111;
assign micromatri[31][47] = 9'b110010110;
assign micromatri[31][48] = 9'b110111111;
assign micromatri[31][49] = 9'b111111111;
assign micromatri[31][50] = 9'b111111111;
assign micromatri[31][51] = 9'b111111111;
assign micromatri[31][52] = 9'b111111111;
assign micromatri[31][53] = 9'b111111111;
assign micromatri[31][54] = 9'b111111111;
assign micromatri[31][55] = 9'b111111111;
assign micromatri[31][56] = 9'b111111111;
assign micromatri[31][57] = 9'b110010110;
assign micromatri[31][58] = 9'b110110110;
assign micromatri[31][59] = 9'b110110010;
assign micromatri[31][60] = 9'b111111111;
assign micromatri[31][61] = 9'b111111111;
assign micromatri[31][62] = 9'b111111111;
assign micromatri[31][63] = 9'b111111111;
assign micromatri[31][64] = 9'b111110111;
assign micromatri[31][65] = 9'b110010001;
assign micromatri[31][66] = 9'b111111111;
assign micromatri[31][67] = 9'b111111111;
assign micromatri[31][68] = 9'b111111111;
assign micromatri[31][69] = 9'b110110110;
assign micromatri[31][70] = 9'b101101101;
assign micromatri[31][71] = 9'b110110011;
assign micromatri[31][72] = 9'b111110111;
assign micromatri[31][73] = 9'b111110111;
assign micromatri[31][74] = 9'b111110111;
assign micromatri[31][75] = 9'b111110111;
assign micromatri[31][76] = 9'b111110011;
assign micromatri[31][77] = 9'b110010010;
assign micromatri[31][78] = 9'b110001101;
assign micromatri[31][79] = 9'b111110111;
assign micromatri[31][80] = 9'b111111111;
assign micromatri[31][81] = 9'b111110111;
assign micromatri[31][82] = 9'b111111111;
assign micromatri[31][83] = 9'b111111111;
assign micromatri[31][84] = 9'b111111111;
assign micromatri[31][85] = 9'b111111111;
assign micromatri[31][86] = 9'b111111111;
assign micromatri[31][87] = 9'b111111111;
assign micromatri[31][88] = 9'b111111111;
assign micromatri[31][89] = 9'b111111111;
assign micromatri[31][90] = 9'b111111111;
assign micromatri[31][91] = 9'b111111111;
assign micromatri[31][92] = 9'b111111111;
assign micromatri[31][93] = 9'b111111111;
assign micromatri[31][94] = 9'b111111111;
assign micromatri[31][95] = 9'b111111111;
assign micromatri[31][96] = 9'b111111111;
assign micromatri[31][97] = 9'b111111111;
assign micromatri[31][98] = 9'b111111111;
assign micromatri[31][99] = 9'b111111111;
assign micromatri[32][0] = 9'b111111111;
assign micromatri[32][1] = 9'b111111111;
assign micromatri[32][2] = 9'b111111111;
assign micromatri[32][3] = 9'b111111111;
assign micromatri[32][4] = 9'b111111111;
assign micromatri[32][5] = 9'b111111111;
assign micromatri[32][6] = 9'b111111111;
assign micromatri[32][7] = 9'b111111111;
assign micromatri[32][8] = 9'b111111111;
assign micromatri[32][9] = 9'b111111111;
assign micromatri[32][10] = 9'b111111111;
assign micromatri[32][11] = 9'b111111111;
assign micromatri[32][12] = 9'b111111111;
assign micromatri[32][13] = 9'b111111111;
assign micromatri[32][14] = 9'b111111111;
assign micromatri[32][15] = 9'b111111111;
assign micromatri[32][16] = 9'b111111111;
assign micromatri[32][17] = 9'b111111111;
assign micromatri[32][18] = 9'b111111111;
assign micromatri[32][19] = 9'b110010001;
assign micromatri[32][20] = 9'b110001101;
assign micromatri[32][21] = 9'b110010001;
assign micromatri[32][22] = 9'b110110010;
assign micromatri[32][23] = 9'b110110010;
assign micromatri[32][24] = 9'b110010001;
assign micromatri[32][25] = 9'b110010010;
assign micromatri[32][26] = 9'b111111111;
assign micromatri[32][27] = 9'b111111111;
assign micromatri[32][28] = 9'b111110111;
assign micromatri[32][29] = 9'b111111111;
assign micromatri[32][30] = 9'b111111111;
assign micromatri[32][31] = 9'b111111111;
assign micromatri[32][32] = 9'b111111111;
assign micromatri[32][33] = 9'b111111111;
assign micromatri[32][34] = 9'b111111111;
assign micromatri[32][35] = 9'b111111111;
assign micromatri[32][36] = 9'b101101101;
assign micromatri[32][37] = 9'b110001110;
assign micromatri[32][38] = 9'b110110010;
assign micromatri[32][39] = 9'b110010010;
assign micromatri[32][40] = 9'b110001110;
assign micromatri[32][41] = 9'b110010001;
assign micromatri[32][42] = 9'b111111111;
assign micromatri[32][43] = 9'b111111111;
assign micromatri[32][44] = 9'b111110111;
assign micromatri[32][45] = 9'b111111111;
assign micromatri[32][46] = 9'b111111111;
assign micromatri[32][47] = 9'b111111111;
assign micromatri[32][48] = 9'b110010001;
assign micromatri[32][49] = 9'b110010010;
assign micromatri[32][50] = 9'b110010110;
assign micromatri[32][51] = 9'b110010010;
assign micromatri[32][52] = 9'b110010110;
assign micromatri[32][53] = 9'b110010110;
assign micromatri[32][54] = 9'b110010110;
assign micromatri[32][55] = 9'b110010110;
assign micromatri[32][56] = 9'b110010110;
assign micromatri[32][57] = 9'b110010110;
assign micromatri[32][58] = 9'b111111111;
assign micromatri[32][59] = 9'b110010001;
assign micromatri[32][60] = 9'b111110010;
assign micromatri[32][61] = 9'b110110010;
assign micromatri[32][62] = 9'b110110010;
assign micromatri[32][63] = 9'b110010001;
assign micromatri[32][64] = 9'b110001101;
assign micromatri[32][65] = 9'b111110010;
assign micromatri[32][66] = 9'b111111111;
assign micromatri[32][67] = 9'b111111111;
assign micromatri[32][68] = 9'b111111111;
assign micromatri[32][69] = 9'b111111111;
assign micromatri[32][70] = 9'b111111111;
assign micromatri[32][71] = 9'b101101101;
assign micromatri[32][72] = 9'b110001101;
assign micromatri[32][73] = 9'b110010010;
assign micromatri[32][74] = 9'b110010010;
assign micromatri[32][75] = 9'b110010010;
assign micromatri[32][76] = 9'b110010010;
assign micromatri[32][77] = 9'b110110010;
assign micromatri[32][78] = 9'b111111111;
assign micromatri[32][79] = 9'b111111111;
assign micromatri[32][80] = 9'b111110111;
assign micromatri[32][81] = 9'b111111111;
assign micromatri[32][82] = 9'b111111111;
assign micromatri[32][83] = 9'b111111111;
assign micromatri[32][84] = 9'b111111111;
assign micromatri[32][85] = 9'b111111111;
assign micromatri[32][86] = 9'b111111111;
assign micromatri[32][87] = 9'b111111111;
assign micromatri[32][88] = 9'b111111111;
assign micromatri[32][89] = 9'b111111111;
assign micromatri[32][90] = 9'b111111111;
assign micromatri[32][91] = 9'b111111111;
assign micromatri[32][92] = 9'b111111111;
assign micromatri[32][93] = 9'b111111111;
assign micromatri[32][94] = 9'b111111111;
assign micromatri[32][95] = 9'b111111111;
assign micromatri[32][96] = 9'b111111111;
assign micromatri[32][97] = 9'b111111111;
assign micromatri[32][98] = 9'b111111111;
assign micromatri[32][99] = 9'b111111111;
assign micromatri[33][0] = 9'b111111111;
assign micromatri[33][1] = 9'b111111111;
assign micromatri[33][2] = 9'b111111111;
assign micromatri[33][3] = 9'b111111111;
assign micromatri[33][4] = 9'b111111111;
assign micromatri[33][5] = 9'b111111111;
assign micromatri[33][6] = 9'b111111111;
assign micromatri[33][7] = 9'b111111111;
assign micromatri[33][8] = 9'b111111111;
assign micromatri[33][9] = 9'b111111111;
assign micromatri[33][10] = 9'b111111111;
assign micromatri[33][11] = 9'b111111111;
assign micromatri[33][12] = 9'b111111111;
assign micromatri[33][13] = 9'b111111111;
assign micromatri[33][14] = 9'b111111111;
assign micromatri[33][15] = 9'b111111111;
assign micromatri[33][16] = 9'b111111111;
assign micromatri[33][17] = 9'b111111111;
assign micromatri[33][18] = 9'b111111111;
assign micromatri[33][19] = 9'b111111111;
assign micromatri[33][20] = 9'b111111111;
assign micromatri[33][21] = 9'b111110111;
assign micromatri[33][22] = 9'b111110111;
assign micromatri[33][23] = 9'b111111111;
assign micromatri[33][24] = 9'b111111111;
assign micromatri[33][25] = 9'b111111111;
assign micromatri[33][26] = 9'b111111111;
assign micromatri[33][27] = 9'b111110111;
assign micromatri[33][28] = 9'b111111111;
assign micromatri[33][29] = 9'b111111111;
assign micromatri[33][30] = 9'b111111111;
assign micromatri[33][31] = 9'b111111111;
assign micromatri[33][32] = 9'b111111111;
assign micromatri[33][33] = 9'b111111111;
assign micromatri[33][34] = 9'b111111111;
assign micromatri[33][35] = 9'b111111111;
assign micromatri[33][36] = 9'b111111111;
assign micromatri[33][37] = 9'b110010010;
assign micromatri[33][38] = 9'b110110010;
assign micromatri[33][39] = 9'b110110111;
assign micromatri[33][40] = 9'b111111111;
assign micromatri[33][41] = 9'b111111111;
assign micromatri[33][42] = 9'b111111111;
assign micromatri[33][43] = 9'b111110111;
assign micromatri[33][44] = 9'b111111111;
assign micromatri[33][45] = 9'b111111111;
assign micromatri[33][46] = 9'b111111111;
assign micromatri[33][47] = 9'b111111111;
assign micromatri[33][48] = 9'b111111111;
assign micromatri[33][49] = 9'b110110110;
assign micromatri[33][50] = 9'b111111111;
assign micromatri[33][51] = 9'b111111111;
assign micromatri[33][52] = 9'b111111111;
assign micromatri[33][53] = 9'b111111111;
assign micromatri[33][54] = 9'b111111111;
assign micromatri[33][55] = 9'b111111111;
assign micromatri[33][56] = 9'b111111111;
assign micromatri[33][57] = 9'b111111111;
assign micromatri[33][58] = 9'b111111111;
assign micromatri[33][59] = 9'b110110110;
assign micromatri[33][60] = 9'b110110110;
assign micromatri[33][61] = 9'b110110010;
assign micromatri[33][62] = 9'b111111111;
assign micromatri[33][63] = 9'b111111111;
assign micromatri[33][64] = 9'b111111111;
assign micromatri[33][65] = 9'b111111111;
assign micromatri[33][66] = 9'b111110111;
assign micromatri[33][67] = 9'b111111111;
assign micromatri[33][68] = 9'b111111111;
assign micromatri[33][69] = 9'b111111111;
assign micromatri[33][70] = 9'b111111111;
assign micromatri[33][71] = 9'b111111111;
assign micromatri[33][72] = 9'b111111111;
assign micromatri[33][73] = 9'b111110111;
assign micromatri[33][74] = 9'b111110111;
assign micromatri[33][75] = 9'b111111111;
assign micromatri[33][76] = 9'b111111111;
assign micromatri[33][77] = 9'b111111111;
assign micromatri[33][78] = 9'b111110111;
assign micromatri[33][79] = 9'b111111111;
assign micromatri[33][80] = 9'b111111111;
assign micromatri[33][81] = 9'b111111111;
assign micromatri[33][82] = 9'b111111111;
assign micromatri[33][83] = 9'b111111111;
assign micromatri[33][84] = 9'b111111111;
assign micromatri[33][85] = 9'b111111111;
assign micromatri[33][86] = 9'b111111111;
assign micromatri[33][87] = 9'b111111111;
assign micromatri[33][88] = 9'b111111111;
assign micromatri[33][89] = 9'b111111111;
assign micromatri[33][90] = 9'b111111111;
assign micromatri[33][91] = 9'b111111111;
assign micromatri[33][92] = 9'b111111111;
assign micromatri[33][93] = 9'b111111111;
assign micromatri[33][94] = 9'b111111111;
assign micromatri[33][95] = 9'b111111111;
assign micromatri[33][96] = 9'b111111111;
assign micromatri[33][97] = 9'b111111111;
assign micromatri[33][98] = 9'b111111111;
assign micromatri[33][99] = 9'b111111111;
assign micromatri[34][0] = 9'b111111111;
assign micromatri[34][1] = 9'b111111111;
assign micromatri[34][2] = 9'b111111111;
assign micromatri[34][3] = 9'b111111111;
assign micromatri[34][4] = 9'b111111111;
assign micromatri[34][5] = 9'b111111111;
assign micromatri[34][6] = 9'b111111111;
assign micromatri[34][7] = 9'b111111111;
assign micromatri[34][8] = 9'b111111111;
assign micromatri[34][9] = 9'b111111111;
assign micromatri[34][10] = 9'b111111111;
assign micromatri[34][11] = 9'b111111111;
assign micromatri[34][12] = 9'b111111111;
assign micromatri[34][13] = 9'b111111111;
assign micromatri[34][14] = 9'b111111111;
assign micromatri[34][15] = 9'b111111111;
assign micromatri[34][16] = 9'b111111111;
assign micromatri[34][17] = 9'b111111111;
assign micromatri[34][18] = 9'b111111111;
assign micromatri[34][19] = 9'b111111111;
assign micromatri[34][20] = 9'b111111111;
assign micromatri[34][21] = 9'b111111111;
assign micromatri[34][22] = 9'b111111111;
assign micromatri[34][23] = 9'b111111111;
assign micromatri[34][24] = 9'b111111111;
assign micromatri[34][25] = 9'b111111111;
assign micromatri[34][26] = 9'b111111111;
assign micromatri[34][27] = 9'b111111111;
assign micromatri[34][28] = 9'b111111111;
assign micromatri[34][29] = 9'b111111111;
assign micromatri[34][30] = 9'b111111111;
assign micromatri[34][31] = 9'b111111111;
assign micromatri[34][32] = 9'b111111111;
assign micromatri[34][33] = 9'b111111111;
assign micromatri[34][34] = 9'b111111111;
assign micromatri[34][35] = 9'b111111111;
assign micromatri[34][36] = 9'b111111111;
assign micromatri[34][37] = 9'b111111111;
assign micromatri[34][38] = 9'b111111111;
assign micromatri[34][39] = 9'b111111111;
assign micromatri[34][40] = 9'b111111111;
assign micromatri[34][41] = 9'b111111111;
assign micromatri[34][42] = 9'b111111111;
assign micromatri[34][43] = 9'b111111111;
assign micromatri[34][44] = 9'b111111111;
assign micromatri[34][45] = 9'b111111111;
assign micromatri[34][46] = 9'b111111111;
assign micromatri[34][47] = 9'b111111111;
assign micromatri[34][48] = 9'b111111111;
assign micromatri[34][49] = 9'b111111111;
assign micromatri[34][50] = 9'b111111111;
assign micromatri[34][51] = 9'b111111111;
assign micromatri[34][52] = 9'b111111111;
assign micromatri[34][53] = 9'b111111111;
assign micromatri[34][54] = 9'b111111111;
assign micromatri[34][55] = 9'b111111111;
assign micromatri[34][56] = 9'b111111111;
assign micromatri[34][57] = 9'b111111111;
assign micromatri[34][58] = 9'b111111111;
assign micromatri[34][59] = 9'b111111111;
assign micromatri[34][60] = 9'b111111111;
assign micromatri[34][61] = 9'b111111111;
assign micromatri[34][62] = 9'b111111111;
assign micromatri[34][63] = 9'b111111111;
assign micromatri[34][64] = 9'b111111111;
assign micromatri[34][65] = 9'b111111111;
assign micromatri[34][66] = 9'b111111111;
assign micromatri[34][67] = 9'b111111111;
assign micromatri[34][68] = 9'b111111111;
assign micromatri[34][69] = 9'b111111111;
assign micromatri[34][70] = 9'b111111111;
assign micromatri[34][71] = 9'b111111111;
assign micromatri[34][72] = 9'b111111111;
assign micromatri[34][73] = 9'b111111111;
assign micromatri[34][74] = 9'b111111111;
assign micromatri[34][75] = 9'b111111111;
assign micromatri[34][76] = 9'b111111111;
assign micromatri[34][77] = 9'b111111111;
assign micromatri[34][78] = 9'b111111111;
assign micromatri[34][79] = 9'b111111111;
assign micromatri[34][80] = 9'b111111111;
assign micromatri[34][81] = 9'b111111111;
assign micromatri[34][82] = 9'b111111111;
assign micromatri[34][83] = 9'b111111111;
assign micromatri[34][84] = 9'b111111111;
assign micromatri[34][85] = 9'b111111111;
assign micromatri[34][86] = 9'b111111111;
assign micromatri[34][87] = 9'b111111111;
assign micromatri[34][88] = 9'b111111111;
assign micromatri[34][89] = 9'b111111111;
assign micromatri[34][90] = 9'b111111111;
assign micromatri[34][91] = 9'b111111111;
assign micromatri[34][92] = 9'b111111111;
assign micromatri[34][93] = 9'b111111111;
assign micromatri[34][94] = 9'b111111111;
assign micromatri[34][95] = 9'b111111111;
assign micromatri[34][96] = 9'b111111111;
assign micromatri[34][97] = 9'b111111111;
assign micromatri[34][98] = 9'b111111111;
assign micromatri[34][99] = 9'b111111111;
assign micromatri[35][0] = 9'b111111111;
assign micromatri[35][1] = 9'b111111111;
assign micromatri[35][2] = 9'b111111111;
assign micromatri[35][3] = 9'b111111111;
assign micromatri[35][4] = 9'b111111111;
assign micromatri[35][5] = 9'b111111111;
assign micromatri[35][6] = 9'b111111111;
assign micromatri[35][7] = 9'b111111111;
assign micromatri[35][8] = 9'b111111111;
assign micromatri[35][9] = 9'b111111111;
assign micromatri[35][10] = 9'b111111111;
assign micromatri[35][11] = 9'b111111111;
assign micromatri[35][12] = 9'b111111111;
assign micromatri[35][13] = 9'b111111111;
assign micromatri[35][14] = 9'b111111111;
assign micromatri[35][15] = 9'b111111111;
assign micromatri[35][16] = 9'b111111111;
assign micromatri[35][17] = 9'b111111111;
assign micromatri[35][18] = 9'b111111111;
assign micromatri[35][19] = 9'b111111111;
assign micromatri[35][20] = 9'b111111111;
assign micromatri[35][21] = 9'b111111111;
assign micromatri[35][22] = 9'b111111111;
assign micromatri[35][23] = 9'b111111111;
assign micromatri[35][24] = 9'b111111111;
assign micromatri[35][25] = 9'b111111111;
assign micromatri[35][26] = 9'b111111111;
assign micromatri[35][27] = 9'b111111111;
assign micromatri[35][28] = 9'b111111111;
assign micromatri[35][29] = 9'b111111111;
assign micromatri[35][30] = 9'b111111111;
assign micromatri[35][31] = 9'b111111111;
assign micromatri[35][32] = 9'b111111111;
assign micromatri[35][33] = 9'b111111111;
assign micromatri[35][34] = 9'b111111111;
assign micromatri[35][35] = 9'b111111111;
assign micromatri[35][36] = 9'b111111111;
assign micromatri[35][37] = 9'b111111111;
assign micromatri[35][38] = 9'b111111111;
assign micromatri[35][39] = 9'b111111111;
assign micromatri[35][40] = 9'b111111111;
assign micromatri[35][41] = 9'b111111111;
assign micromatri[35][42] = 9'b111111111;
assign micromatri[35][43] = 9'b111111111;
assign micromatri[35][44] = 9'b111111111;
assign micromatri[35][45] = 9'b111111111;
assign micromatri[35][46] = 9'b111111111;
assign micromatri[35][47] = 9'b111111111;
assign micromatri[35][48] = 9'b111111111;
assign micromatri[35][49] = 9'b111111111;
assign micromatri[35][50] = 9'b111111111;
assign micromatri[35][51] = 9'b111111111;
assign micromatri[35][52] = 9'b111111111;
assign micromatri[35][53] = 9'b111111111;
assign micromatri[35][54] = 9'b111111111;
assign micromatri[35][55] = 9'b111111111;
assign micromatri[35][56] = 9'b111111111;
assign micromatri[35][57] = 9'b111111111;
assign micromatri[35][58] = 9'b111111111;
assign micromatri[35][59] = 9'b111111111;
assign micromatri[35][60] = 9'b111111111;
assign micromatri[35][61] = 9'b111111111;
assign micromatri[35][62] = 9'b111111111;
assign micromatri[35][63] = 9'b111111111;
assign micromatri[35][64] = 9'b111111111;
assign micromatri[35][65] = 9'b111111111;
assign micromatri[35][66] = 9'b111111111;
assign micromatri[35][67] = 9'b111111111;
assign micromatri[35][68] = 9'b111111111;
assign micromatri[35][69] = 9'b111111111;
assign micromatri[35][70] = 9'b111111111;
assign micromatri[35][71] = 9'b111111111;
assign micromatri[35][72] = 9'b111111111;
assign micromatri[35][73] = 9'b111111111;
assign micromatri[35][74] = 9'b111111111;
assign micromatri[35][75] = 9'b111111111;
assign micromatri[35][76] = 9'b111111111;
assign micromatri[35][77] = 9'b111111111;
assign micromatri[35][78] = 9'b111111111;
assign micromatri[35][79] = 9'b111111111;
assign micromatri[35][80] = 9'b111111111;
assign micromatri[35][81] = 9'b111111111;
assign micromatri[35][82] = 9'b111111111;
assign micromatri[35][83] = 9'b111111111;
assign micromatri[35][84] = 9'b111111111;
assign micromatri[35][85] = 9'b111111111;
assign micromatri[35][86] = 9'b111111111;
assign micromatri[35][87] = 9'b111111111;
assign micromatri[35][88] = 9'b111111111;
assign micromatri[35][89] = 9'b111111111;
assign micromatri[35][90] = 9'b111111111;
assign micromatri[35][91] = 9'b111111111;
assign micromatri[35][92] = 9'b111111111;
assign micromatri[35][93] = 9'b111111111;
assign micromatri[35][94] = 9'b111111111;
assign micromatri[35][95] = 9'b111111111;
assign micromatri[35][96] = 9'b111111111;
assign micromatri[35][97] = 9'b111111111;
assign micromatri[35][98] = 9'b111111111;
assign micromatri[35][99] = 9'b111111111;
assign micromatri[36][0] = 9'b111111111;
assign micromatri[36][1] = 9'b111111111;
assign micromatri[36][2] = 9'b111111111;
assign micromatri[36][3] = 9'b111111111;
assign micromatri[36][4] = 9'b111111111;
assign micromatri[36][5] = 9'b111111111;
assign micromatri[36][6] = 9'b111111111;
assign micromatri[36][7] = 9'b111111111;
assign micromatri[36][8] = 9'b111111111;
assign micromatri[36][9] = 9'b111111111;
assign micromatri[36][10] = 9'b111111111;
assign micromatri[36][11] = 9'b111111111;
assign micromatri[36][12] = 9'b111111111;
assign micromatri[36][13] = 9'b111111111;
assign micromatri[36][14] = 9'b111111111;
assign micromatri[36][15] = 9'b111111111;
assign micromatri[36][16] = 9'b111111111;
assign micromatri[36][17] = 9'b111111111;
assign micromatri[36][18] = 9'b111111111;
assign micromatri[36][19] = 9'b111111111;
assign micromatri[36][20] = 9'b111111111;
assign micromatri[36][21] = 9'b111111111;
assign micromatri[36][22] = 9'b111111111;
assign micromatri[36][23] = 9'b111111111;
assign micromatri[36][24] = 9'b111111111;
assign micromatri[36][25] = 9'b111111111;
assign micromatri[36][26] = 9'b111111111;
assign micromatri[36][27] = 9'b111111111;
assign micromatri[36][28] = 9'b111111111;
assign micromatri[36][29] = 9'b111111111;
assign micromatri[36][30] = 9'b111111111;
assign micromatri[36][31] = 9'b111111111;
assign micromatri[36][32] = 9'b111111111;
assign micromatri[36][33] = 9'b111111111;
assign micromatri[36][34] = 9'b111111111;
assign micromatri[36][35] = 9'b111111111;
assign micromatri[36][36] = 9'b111111111;
assign micromatri[36][37] = 9'b111111111;
assign micromatri[36][38] = 9'b111111111;
assign micromatri[36][39] = 9'b111111111;
assign micromatri[36][40] = 9'b111111111;
assign micromatri[36][41] = 9'b111111111;
assign micromatri[36][42] = 9'b111111111;
assign micromatri[36][43] = 9'b111111111;
assign micromatri[36][44] = 9'b111111111;
assign micromatri[36][45] = 9'b111111111;
assign micromatri[36][46] = 9'b111111111;
assign micromatri[36][47] = 9'b111111111;
assign micromatri[36][48] = 9'b111111111;
assign micromatri[36][49] = 9'b111111111;
assign micromatri[36][50] = 9'b111111111;
assign micromatri[36][51] = 9'b111111111;
assign micromatri[36][52] = 9'b111111111;
assign micromatri[36][53] = 9'b111111111;
assign micromatri[36][54] = 9'b111111111;
assign micromatri[36][55] = 9'b111111111;
assign micromatri[36][56] = 9'b111111111;
assign micromatri[36][57] = 9'b111111111;
assign micromatri[36][58] = 9'b111111111;
assign micromatri[36][59] = 9'b111111111;
assign micromatri[36][60] = 9'b111111111;
assign micromatri[36][61] = 9'b111111111;
assign micromatri[36][62] = 9'b111111111;
assign micromatri[36][63] = 9'b111111111;
assign micromatri[36][64] = 9'b111111111;
assign micromatri[36][65] = 9'b111111111;
assign micromatri[36][66] = 9'b111111111;
assign micromatri[36][67] = 9'b111111111;
assign micromatri[36][68] = 9'b111111111;
assign micromatri[36][69] = 9'b111111111;
assign micromatri[36][70] = 9'b111111111;
assign micromatri[36][71] = 9'b111111111;
assign micromatri[36][72] = 9'b111111111;
assign micromatri[36][73] = 9'b111111111;
assign micromatri[36][74] = 9'b111111111;
assign micromatri[36][75] = 9'b111111111;
assign micromatri[36][76] = 9'b111111111;
assign micromatri[36][77] = 9'b111111111;
assign micromatri[36][78] = 9'b111111111;
assign micromatri[36][79] = 9'b111111111;
assign micromatri[36][80] = 9'b111111111;
assign micromatri[36][81] = 9'b111111111;
assign micromatri[36][82] = 9'b111111111;
assign micromatri[36][83] = 9'b111111111;
assign micromatri[36][84] = 9'b111111111;
assign micromatri[36][85] = 9'b111111111;
assign micromatri[36][86] = 9'b111111111;
assign micromatri[36][87] = 9'b111111111;
assign micromatri[36][88] = 9'b111111111;
assign micromatri[36][89] = 9'b111111111;
assign micromatri[36][90] = 9'b111111111;
assign micromatri[36][91] = 9'b111111111;
assign micromatri[36][92] = 9'b111111111;
assign micromatri[36][93] = 9'b111111111;
assign micromatri[36][94] = 9'b111111111;
assign micromatri[36][95] = 9'b111111111;
assign micromatri[36][96] = 9'b111111111;
assign micromatri[36][97] = 9'b111111111;
assign micromatri[36][98] = 9'b111111111;
assign micromatri[36][99] = 9'b111111111;
assign micromatri[37][0] = 9'b111111111;
assign micromatri[37][1] = 9'b111111111;
assign micromatri[37][2] = 9'b111111111;
assign micromatri[37][3] = 9'b111111111;
assign micromatri[37][4] = 9'b111111111;
assign micromatri[37][5] = 9'b111111111;
assign micromatri[37][6] = 9'b111111111;
assign micromatri[37][7] = 9'b111111111;
assign micromatri[37][8] = 9'b111111111;
assign micromatri[37][9] = 9'b111111111;
assign micromatri[37][10] = 9'b111111111;
assign micromatri[37][11] = 9'b111111111;
assign micromatri[37][12] = 9'b111111111;
assign micromatri[37][13] = 9'b111111111;
assign micromatri[37][14] = 9'b111111111;
assign micromatri[37][15] = 9'b111111111;
assign micromatri[37][16] = 9'b111111111;
assign micromatri[37][17] = 9'b111111111;
assign micromatri[37][18] = 9'b111111111;
assign micromatri[37][19] = 9'b111111111;
assign micromatri[37][20] = 9'b111111111;
assign micromatri[37][21] = 9'b111111111;
assign micromatri[37][22] = 9'b111111111;
assign micromatri[37][23] = 9'b111111111;
assign micromatri[37][24] = 9'b111111111;
assign micromatri[37][25] = 9'b111111111;
assign micromatri[37][26] = 9'b111111111;
assign micromatri[37][27] = 9'b111111111;
assign micromatri[37][28] = 9'b111111111;
assign micromatri[37][29] = 9'b111111111;
assign micromatri[37][30] = 9'b111111111;
assign micromatri[37][31] = 9'b111111111;
assign micromatri[37][32] = 9'b111111111;
assign micromatri[37][33] = 9'b111111111;
assign micromatri[37][34] = 9'b111111111;
assign micromatri[37][35] = 9'b111111111;
assign micromatri[37][36] = 9'b111111111;
assign micromatri[37][37] = 9'b111111111;
assign micromatri[37][38] = 9'b111111111;
assign micromatri[37][39] = 9'b111111111;
assign micromatri[37][40] = 9'b111111111;
assign micromatri[37][41] = 9'b111111111;
assign micromatri[37][42] = 9'b111111111;
assign micromatri[37][43] = 9'b111111111;
assign micromatri[37][44] = 9'b111111111;
assign micromatri[37][45] = 9'b111111111;
assign micromatri[37][46] = 9'b111111111;
assign micromatri[37][47] = 9'b111111111;
assign micromatri[37][48] = 9'b111111111;
assign micromatri[37][49] = 9'b111111111;
assign micromatri[37][50] = 9'b111111111;
assign micromatri[37][51] = 9'b111111111;
assign micromatri[37][52] = 9'b111111111;
assign micromatri[37][53] = 9'b111111111;
assign micromatri[37][54] = 9'b111111111;
assign micromatri[37][55] = 9'b111111111;
assign micromatri[37][56] = 9'b111111111;
assign micromatri[37][57] = 9'b111111111;
assign micromatri[37][58] = 9'b111111111;
assign micromatri[37][59] = 9'b111111111;
assign micromatri[37][60] = 9'b111111111;
assign micromatri[37][61] = 9'b111111111;
assign micromatri[37][62] = 9'b111111111;
assign micromatri[37][63] = 9'b111111111;
assign micromatri[37][64] = 9'b111111111;
assign micromatri[37][65] = 9'b111111111;
assign micromatri[37][66] = 9'b111111111;
assign micromatri[37][67] = 9'b111111111;
assign micromatri[37][68] = 9'b111111111;
assign micromatri[37][69] = 9'b111111111;
assign micromatri[37][70] = 9'b111111111;
assign micromatri[37][71] = 9'b111111111;
assign micromatri[37][72] = 9'b111111111;
assign micromatri[37][73] = 9'b111111111;
assign micromatri[37][74] = 9'b111111111;
assign micromatri[37][75] = 9'b111111111;
assign micromatri[37][76] = 9'b111111111;
assign micromatri[37][77] = 9'b111111111;
assign micromatri[37][78] = 9'b111111111;
assign micromatri[37][79] = 9'b111111111;
assign micromatri[37][80] = 9'b111111111;
assign micromatri[37][81] = 9'b111111111;
assign micromatri[37][82] = 9'b111111111;
assign micromatri[37][83] = 9'b111111111;
assign micromatri[37][84] = 9'b111111111;
assign micromatri[37][85] = 9'b111111111;
assign micromatri[37][86] = 9'b111111111;
assign micromatri[37][87] = 9'b111111111;
assign micromatri[37][88] = 9'b111111111;
assign micromatri[37][89] = 9'b111111111;
assign micromatri[37][90] = 9'b111111111;
assign micromatri[37][91] = 9'b111111111;
assign micromatri[37][92] = 9'b111111111;
assign micromatri[37][93] = 9'b111111111;
assign micromatri[37][94] = 9'b111111111;
assign micromatri[37][95] = 9'b111111111;
assign micromatri[37][96] = 9'b111111111;
assign micromatri[37][97] = 9'b111111111;
assign micromatri[37][98] = 9'b111111111;
assign micromatri[37][99] = 9'b111111111;
assign micromatri[38][0] = 9'b111111111;
assign micromatri[38][1] = 9'b111111111;
assign micromatri[38][2] = 9'b111111111;
assign micromatri[38][3] = 9'b111111111;
assign micromatri[38][4] = 9'b111111111;
assign micromatri[38][5] = 9'b111111111;
assign micromatri[38][6] = 9'b111111111;
assign micromatri[38][7] = 9'b111111111;
assign micromatri[38][8] = 9'b111111111;
assign micromatri[38][9] = 9'b111111111;
assign micromatri[38][10] = 9'b111111111;
assign micromatri[38][11] = 9'b111111111;
assign micromatri[38][12] = 9'b111111111;
assign micromatri[38][13] = 9'b111111111;
assign micromatri[38][14] = 9'b111111111;
assign micromatri[38][15] = 9'b111111111;
assign micromatri[38][16] = 9'b111111111;
assign micromatri[38][17] = 9'b111111111;
assign micromatri[38][18] = 9'b111111111;
assign micromatri[38][19] = 9'b111111111;
assign micromatri[38][20] = 9'b111111111;
assign micromatri[38][21] = 9'b111111111;
assign micromatri[38][22] = 9'b111111111;
assign micromatri[38][23] = 9'b111111111;
assign micromatri[38][24] = 9'b111111111;
assign micromatri[38][25] = 9'b111111111;
assign micromatri[38][26] = 9'b111111111;
assign micromatri[38][27] = 9'b111111111;
assign micromatri[38][28] = 9'b111111111;
assign micromatri[38][29] = 9'b111111111;
assign micromatri[38][30] = 9'b111111111;
assign micromatri[38][31] = 9'b111111111;
assign micromatri[38][32] = 9'b111111111;
assign micromatri[38][33] = 9'b111111111;
assign micromatri[38][34] = 9'b111111111;
assign micromatri[38][35] = 9'b111111111;
assign micromatri[38][36] = 9'b111111111;
assign micromatri[38][37] = 9'b111111111;
assign micromatri[38][38] = 9'b111111111;
assign micromatri[38][39] = 9'b111111111;
assign micromatri[38][40] = 9'b111111111;
assign micromatri[38][41] = 9'b111111111;
assign micromatri[38][42] = 9'b111111111;
assign micromatri[38][43] = 9'b111111111;
assign micromatri[38][44] = 9'b111111111;
assign micromatri[38][45] = 9'b111111111;
assign micromatri[38][46] = 9'b111111111;
assign micromatri[38][47] = 9'b111111111;
assign micromatri[38][48] = 9'b111111111;
assign micromatri[38][49] = 9'b111111111;
assign micromatri[38][50] = 9'b111111111;
assign micromatri[38][51] = 9'b111111111;
assign micromatri[38][52] = 9'b111111111;
assign micromatri[38][53] = 9'b111111111;
assign micromatri[38][54] = 9'b111111111;
assign micromatri[38][55] = 9'b111111111;
assign micromatri[38][56] = 9'b111111111;
assign micromatri[38][57] = 9'b111111111;
assign micromatri[38][58] = 9'b111111111;
assign micromatri[38][59] = 9'b111111111;
assign micromatri[38][60] = 9'b111111111;
assign micromatri[38][61] = 9'b111111111;
assign micromatri[38][62] = 9'b111111111;
assign micromatri[38][63] = 9'b111111111;
assign micromatri[38][64] = 9'b111111111;
assign micromatri[38][65] = 9'b111111111;
assign micromatri[38][66] = 9'b111111111;
assign micromatri[38][67] = 9'b111111111;
assign micromatri[38][68] = 9'b111111111;
assign micromatri[38][69] = 9'b111111111;
assign micromatri[38][70] = 9'b111111111;
assign micromatri[38][71] = 9'b111111111;
assign micromatri[38][72] = 9'b111111111;
assign micromatri[38][73] = 9'b111111111;
assign micromatri[38][74] = 9'b111111111;
assign micromatri[38][75] = 9'b111111111;
assign micromatri[38][76] = 9'b111111111;
assign micromatri[38][77] = 9'b111111111;
assign micromatri[38][78] = 9'b111111111;
assign micromatri[38][79] = 9'b111111111;
assign micromatri[38][80] = 9'b111111111;
assign micromatri[38][81] = 9'b111111111;
assign micromatri[38][82] = 9'b111111111;
assign micromatri[38][83] = 9'b111111111;
assign micromatri[38][84] = 9'b111111111;
assign micromatri[38][85] = 9'b111111111;
assign micromatri[38][86] = 9'b111111111;
assign micromatri[38][87] = 9'b111111111;
assign micromatri[38][88] = 9'b111111111;
assign micromatri[38][89] = 9'b111111111;
assign micromatri[38][90] = 9'b111111111;
assign micromatri[38][91] = 9'b111111111;
assign micromatri[38][92] = 9'b111111111;
assign micromatri[38][93] = 9'b111111111;
assign micromatri[38][94] = 9'b111111111;
assign micromatri[38][95] = 9'b111111111;
assign micromatri[38][96] = 9'b111111111;
assign micromatri[38][97] = 9'b111111111;
assign micromatri[38][98] = 9'b111111111;
assign micromatri[38][99] = 9'b111111111;
assign micromatri[39][0] = 9'b111111111;
assign micromatri[39][1] = 9'b111111111;
assign micromatri[39][2] = 9'b111111111;
assign micromatri[39][3] = 9'b111111111;
assign micromatri[39][4] = 9'b111111111;
assign micromatri[39][5] = 9'b111111111;
assign micromatri[39][6] = 9'b111111111;
assign micromatri[39][7] = 9'b111111111;
assign micromatri[39][8] = 9'b111111111;
assign micromatri[39][9] = 9'b111111111;
assign micromatri[39][10] = 9'b111111111;
assign micromatri[39][11] = 9'b111111111;
assign micromatri[39][12] = 9'b111111111;
assign micromatri[39][13] = 9'b111111111;
assign micromatri[39][14] = 9'b111111111;
assign micromatri[39][15] = 9'b111111111;
assign micromatri[39][16] = 9'b111111111;
assign micromatri[39][17] = 9'b111111111;
assign micromatri[39][18] = 9'b111111111;
assign micromatri[39][19] = 9'b111111111;
assign micromatri[39][20] = 9'b111111111;
assign micromatri[39][21] = 9'b111111111;
assign micromatri[39][22] = 9'b111111111;
assign micromatri[39][23] = 9'b111111111;
assign micromatri[39][24] = 9'b111111111;
assign micromatri[39][25] = 9'b111111111;
assign micromatri[39][26] = 9'b111111111;
assign micromatri[39][27] = 9'b111111111;
assign micromatri[39][28] = 9'b111111111;
assign micromatri[39][29] = 9'b111111111;
assign micromatri[39][30] = 9'b111111111;
assign micromatri[39][31] = 9'b111111111;
assign micromatri[39][32] = 9'b111111111;
assign micromatri[39][33] = 9'b111111111;
assign micromatri[39][34] = 9'b111111111;
assign micromatri[39][35] = 9'b111111111;
assign micromatri[39][36] = 9'b111111111;
assign micromatri[39][37] = 9'b111111111;
assign micromatri[39][38] = 9'b111111111;
assign micromatri[39][39] = 9'b111111111;
assign micromatri[39][40] = 9'b111111111;
assign micromatri[39][41] = 9'b111111111;
assign micromatri[39][42] = 9'b111111111;
assign micromatri[39][43] = 9'b111111111;
assign micromatri[39][44] = 9'b111111111;
assign micromatri[39][45] = 9'b111111111;
assign micromatri[39][46] = 9'b111111111;
assign micromatri[39][47] = 9'b111111111;
assign micromatri[39][48] = 9'b111111111;
assign micromatri[39][49] = 9'b111111111;
assign micromatri[39][50] = 9'b111111111;
assign micromatri[39][51] = 9'b111111111;
assign micromatri[39][52] = 9'b111111111;
assign micromatri[39][53] = 9'b111111111;
assign micromatri[39][54] = 9'b111111111;
assign micromatri[39][55] = 9'b111111111;
assign micromatri[39][56] = 9'b111111111;
assign micromatri[39][57] = 9'b111111111;
assign micromatri[39][58] = 9'b111111111;
assign micromatri[39][59] = 9'b111111111;
assign micromatri[39][60] = 9'b111111111;
assign micromatri[39][61] = 9'b111111111;
assign micromatri[39][62] = 9'b111111111;
assign micromatri[39][63] = 9'b111111111;
assign micromatri[39][64] = 9'b111111111;
assign micromatri[39][65] = 9'b111111111;
assign micromatri[39][66] = 9'b111111111;
assign micromatri[39][67] = 9'b111111111;
assign micromatri[39][68] = 9'b111111111;
assign micromatri[39][69] = 9'b111111111;
assign micromatri[39][70] = 9'b111111111;
assign micromatri[39][71] = 9'b111111111;
assign micromatri[39][72] = 9'b111111111;
assign micromatri[39][73] = 9'b111111111;
assign micromatri[39][74] = 9'b111111111;
assign micromatri[39][75] = 9'b111111111;
assign micromatri[39][76] = 9'b111111111;
assign micromatri[39][77] = 9'b111111111;
assign micromatri[39][78] = 9'b111111111;
assign micromatri[39][79] = 9'b111111111;
assign micromatri[39][80] = 9'b111111111;
assign micromatri[39][81] = 9'b111111111;
assign micromatri[39][82] = 9'b111111111;
assign micromatri[39][83] = 9'b111111111;
assign micromatri[39][84] = 9'b111111111;
assign micromatri[39][85] = 9'b111111111;
assign micromatri[39][86] = 9'b111111111;
assign micromatri[39][87] = 9'b111111111;
assign micromatri[39][88] = 9'b111111111;
assign micromatri[39][89] = 9'b111111111;
assign micromatri[39][90] = 9'b111111111;
assign micromatri[39][91] = 9'b111111111;
assign micromatri[39][92] = 9'b111111111;
assign micromatri[39][93] = 9'b111111111;
assign micromatri[39][94] = 9'b111111111;
assign micromatri[39][95] = 9'b111111111;
assign micromatri[39][96] = 9'b111111111;
assign micromatri[39][97] = 9'b111111111;
assign micromatri[39][98] = 9'b111111111;
assign micromatri[39][99] = 9'b111111111;
assign micromatri[40][0] = 9'b111111111;
assign micromatri[40][1] = 9'b111111111;
assign micromatri[40][2] = 9'b111111111;
assign micromatri[40][3] = 9'b111111111;
assign micromatri[40][4] = 9'b111111111;
assign micromatri[40][5] = 9'b111111111;
assign micromatri[40][6] = 9'b111111111;
assign micromatri[40][7] = 9'b111111111;
assign micromatri[40][8] = 9'b111111111;
assign micromatri[40][9] = 9'b111111111;
assign micromatri[40][10] = 9'b111111111;
assign micromatri[40][11] = 9'b111111111;
assign micromatri[40][12] = 9'b111111111;
assign micromatri[40][13] = 9'b111111111;
assign micromatri[40][14] = 9'b111111111;
assign micromatri[40][15] = 9'b111111111;
assign micromatri[40][16] = 9'b111111111;
assign micromatri[40][17] = 9'b111111111;
assign micromatri[40][18] = 9'b111111111;
assign micromatri[40][19] = 9'b111111111;
assign micromatri[40][20] = 9'b111111111;
assign micromatri[40][21] = 9'b111111111;
assign micromatri[40][22] = 9'b111111111;
assign micromatri[40][23] = 9'b111111111;
assign micromatri[40][24] = 9'b111111111;
assign micromatri[40][25] = 9'b111111111;
assign micromatri[40][26] = 9'b111111111;
assign micromatri[40][27] = 9'b111111111;
assign micromatri[40][28] = 9'b111111111;
assign micromatri[40][29] = 9'b111111111;
assign micromatri[40][30] = 9'b111111111;
assign micromatri[40][31] = 9'b111111111;
assign micromatri[40][32] = 9'b111111111;
assign micromatri[40][33] = 9'b111111111;
assign micromatri[40][34] = 9'b111111111;
assign micromatri[40][35] = 9'b111111111;
assign micromatri[40][36] = 9'b111111111;
assign micromatri[40][37] = 9'b111111111;
assign micromatri[40][38] = 9'b111111111;
assign micromatri[40][39] = 9'b111111111;
assign micromatri[40][40] = 9'b111111111;
assign micromatri[40][41] = 9'b111111111;
assign micromatri[40][42] = 9'b111111111;
assign micromatri[40][43] = 9'b111111111;
assign micromatri[40][44] = 9'b111111111;
assign micromatri[40][45] = 9'b111111111;
assign micromatri[40][46] = 9'b111111111;
assign micromatri[40][47] = 9'b111111111;
assign micromatri[40][48] = 9'b111111111;
assign micromatri[40][49] = 9'b111111111;
assign micromatri[40][50] = 9'b111111111;
assign micromatri[40][51] = 9'b111111111;
assign micromatri[40][52] = 9'b111111111;
assign micromatri[40][53] = 9'b111111111;
assign micromatri[40][54] = 9'b111111111;
assign micromatri[40][55] = 9'b111111111;
assign micromatri[40][56] = 9'b111111111;
assign micromatri[40][57] = 9'b111111111;
assign micromatri[40][58] = 9'b111111111;
assign micromatri[40][59] = 9'b111111111;
assign micromatri[40][60] = 9'b111111111;
assign micromatri[40][61] = 9'b111111111;
assign micromatri[40][62] = 9'b111111111;
assign micromatri[40][63] = 9'b111111111;
assign micromatri[40][64] = 9'b111111111;
assign micromatri[40][65] = 9'b111111111;
assign micromatri[40][66] = 9'b111111111;
assign micromatri[40][67] = 9'b111111111;
assign micromatri[40][68] = 9'b111111111;
assign micromatri[40][69] = 9'b111111111;
assign micromatri[40][70] = 9'b111111111;
assign micromatri[40][71] = 9'b111111111;
assign micromatri[40][72] = 9'b111111111;
assign micromatri[40][73] = 9'b111111111;
assign micromatri[40][74] = 9'b111111111;
assign micromatri[40][75] = 9'b111111111;
assign micromatri[40][76] = 9'b111111111;
assign micromatri[40][77] = 9'b111111111;
assign micromatri[40][78] = 9'b111111111;
assign micromatri[40][79] = 9'b111111111;
assign micromatri[40][80] = 9'b111111111;
assign micromatri[40][81] = 9'b111111111;
assign micromatri[40][82] = 9'b111111111;
assign micromatri[40][83] = 9'b111111111;
assign micromatri[40][84] = 9'b111111111;
assign micromatri[40][85] = 9'b111111111;
assign micromatri[40][86] = 9'b111111111;
assign micromatri[40][87] = 9'b111111111;
assign micromatri[40][88] = 9'b111111111;
assign micromatri[40][89] = 9'b111111111;
assign micromatri[40][90] = 9'b111111111;
assign micromatri[40][91] = 9'b111111111;
assign micromatri[40][92] = 9'b111111111;
assign micromatri[40][93] = 9'b111111111;
assign micromatri[40][94] = 9'b111111111;
assign micromatri[40][95] = 9'b111111111;
assign micromatri[40][96] = 9'b111111111;
assign micromatri[40][97] = 9'b111111111;
assign micromatri[40][98] = 9'b111111111;
assign micromatri[40][99] = 9'b111111111;
assign micromatri[41][0] = 9'b111111111;
assign micromatri[41][1] = 9'b111111111;
assign micromatri[41][2] = 9'b111111111;
assign micromatri[41][3] = 9'b111111111;
assign micromatri[41][4] = 9'b111111111;
assign micromatri[41][5] = 9'b111111111;
assign micromatri[41][6] = 9'b111111111;
assign micromatri[41][7] = 9'b111111111;
assign micromatri[41][8] = 9'b111111111;
assign micromatri[41][9] = 9'b111111111;
assign micromatri[41][10] = 9'b111111111;
assign micromatri[41][11] = 9'b111111111;
assign micromatri[41][12] = 9'b111111111;
assign micromatri[41][13] = 9'b111111111;
assign micromatri[41][14] = 9'b111111111;
assign micromatri[41][15] = 9'b111111111;
assign micromatri[41][16] = 9'b111111111;
assign micromatri[41][17] = 9'b111111111;
assign micromatri[41][18] = 9'b111111111;
assign micromatri[41][19] = 9'b111111111;
assign micromatri[41][20] = 9'b111111111;
assign micromatri[41][21] = 9'b111111111;
assign micromatri[41][22] = 9'b111111111;
assign micromatri[41][23] = 9'b111111111;
assign micromatri[41][24] = 9'b111111111;
assign micromatri[41][25] = 9'b111111111;
assign micromatri[41][26] = 9'b111111111;
assign micromatri[41][27] = 9'b111111111;
assign micromatri[41][28] = 9'b111111111;
assign micromatri[41][29] = 9'b111111111;
assign micromatri[41][30] = 9'b111111111;
assign micromatri[41][31] = 9'b111111111;
assign micromatri[41][32] = 9'b111111111;
assign micromatri[41][33] = 9'b111111111;
assign micromatri[41][34] = 9'b111111111;
assign micromatri[41][35] = 9'b111111111;
assign micromatri[41][36] = 9'b111111111;
assign micromatri[41][37] = 9'b111111111;
assign micromatri[41][38] = 9'b111111111;
assign micromatri[41][39] = 9'b111111111;
assign micromatri[41][40] = 9'b111111111;
assign micromatri[41][41] = 9'b111111111;
assign micromatri[41][42] = 9'b111111111;
assign micromatri[41][43] = 9'b111111111;
assign micromatri[41][44] = 9'b111111111;
assign micromatri[41][45] = 9'b111111111;
assign micromatri[41][46] = 9'b111111111;
assign micromatri[41][47] = 9'b111111111;
assign micromatri[41][48] = 9'b111111111;
assign micromatri[41][49] = 9'b111111111;
assign micromatri[41][50] = 9'b111111111;
assign micromatri[41][51] = 9'b111111111;
assign micromatri[41][52] = 9'b111111111;
assign micromatri[41][53] = 9'b111111111;
assign micromatri[41][54] = 9'b111111111;
assign micromatri[41][55] = 9'b111111111;
assign micromatri[41][56] = 9'b111111111;
assign micromatri[41][57] = 9'b111111111;
assign micromatri[41][58] = 9'b111111111;
assign micromatri[41][59] = 9'b111111111;
assign micromatri[41][60] = 9'b111111111;
assign micromatri[41][61] = 9'b111111111;
assign micromatri[41][62] = 9'b111111111;
assign micromatri[41][63] = 9'b111111111;
assign micromatri[41][64] = 9'b111111111;
assign micromatri[41][65] = 9'b111111111;
assign micromatri[41][66] = 9'b111111111;
assign micromatri[41][67] = 9'b111111111;
assign micromatri[41][68] = 9'b111111111;
assign micromatri[41][69] = 9'b111111111;
assign micromatri[41][70] = 9'b111111111;
assign micromatri[41][71] = 9'b111111111;
assign micromatri[41][72] = 9'b111111111;
assign micromatri[41][73] = 9'b111111111;
assign micromatri[41][74] = 9'b111111111;
assign micromatri[41][75] = 9'b111111111;
assign micromatri[41][76] = 9'b111111111;
assign micromatri[41][77] = 9'b111111111;
assign micromatri[41][78] = 9'b111111111;
assign micromatri[41][79] = 9'b111111111;
assign micromatri[41][80] = 9'b111111111;
assign micromatri[41][81] = 9'b111111111;
assign micromatri[41][82] = 9'b111111111;
assign micromatri[41][83] = 9'b111111111;
assign micromatri[41][84] = 9'b111111111;
assign micromatri[41][85] = 9'b111111111;
assign micromatri[41][86] = 9'b111111111;
assign micromatri[41][87] = 9'b111111111;
assign micromatri[41][88] = 9'b111111111;
assign micromatri[41][89] = 9'b111111111;
assign micromatri[41][90] = 9'b111111111;
assign micromatri[41][91] = 9'b111111111;
assign micromatri[41][92] = 9'b111111111;
assign micromatri[41][93] = 9'b111111111;
assign micromatri[41][94] = 9'b111111111;
assign micromatri[41][95] = 9'b111111111;
assign micromatri[41][96] = 9'b111111111;
assign micromatri[41][97] = 9'b111111111;
assign micromatri[41][98] = 9'b111111111;
assign micromatri[41][99] = 9'b111111111;
assign micromatri[42][0] = 9'b111111111;
assign micromatri[42][1] = 9'b111111111;
assign micromatri[42][2] = 9'b111111111;
assign micromatri[42][3] = 9'b111111111;
assign micromatri[42][4] = 9'b111111111;
assign micromatri[42][5] = 9'b111111111;
assign micromatri[42][6] = 9'b111111111;
assign micromatri[42][7] = 9'b111111111;
assign micromatri[42][8] = 9'b111111111;
assign micromatri[42][9] = 9'b111111111;
assign micromatri[42][10] = 9'b111111111;
assign micromatri[42][11] = 9'b111111111;
assign micromatri[42][12] = 9'b111111111;
assign micromatri[42][13] = 9'b111111111;
assign micromatri[42][14] = 9'b111111111;
assign micromatri[42][15] = 9'b111111111;
assign micromatri[42][16] = 9'b111111111;
assign micromatri[42][17] = 9'b111111111;
assign micromatri[42][18] = 9'b111111111;
assign micromatri[42][19] = 9'b111111111;
assign micromatri[42][20] = 9'b111111111;
assign micromatri[42][21] = 9'b111111111;
assign micromatri[42][22] = 9'b111111111;
assign micromatri[42][23] = 9'b111111111;
assign micromatri[42][24] = 9'b111111111;
assign micromatri[42][25] = 9'b111111111;
assign micromatri[42][26] = 9'b111111111;
assign micromatri[42][27] = 9'b111111111;
assign micromatri[42][28] = 9'b111111111;
assign micromatri[42][29] = 9'b111111111;
assign micromatri[42][30] = 9'b111111111;
assign micromatri[42][31] = 9'b111111111;
assign micromatri[42][32] = 9'b111111111;
assign micromatri[42][33] = 9'b111111111;
assign micromatri[42][34] = 9'b111111111;
assign micromatri[42][35] = 9'b111111111;
assign micromatri[42][36] = 9'b111111111;
assign micromatri[42][37] = 9'b111111111;
assign micromatri[42][38] = 9'b111111111;
assign micromatri[42][39] = 9'b111111111;
assign micromatri[42][40] = 9'b111111111;
assign micromatri[42][41] = 9'b111111111;
assign micromatri[42][42] = 9'b111111111;
assign micromatri[42][43] = 9'b111111111;
assign micromatri[42][44] = 9'b111111111;
assign micromatri[42][45] = 9'b111111111;
assign micromatri[42][46] = 9'b111111111;
assign micromatri[42][47] = 9'b111111111;
assign micromatri[42][48] = 9'b111111111;
assign micromatri[42][49] = 9'b111111111;
assign micromatri[42][50] = 9'b111111111;
assign micromatri[42][51] = 9'b111111111;
assign micromatri[42][52] = 9'b111111111;
assign micromatri[42][53] = 9'b111111111;
assign micromatri[42][54] = 9'b111111111;
assign micromatri[42][55] = 9'b111111111;
assign micromatri[42][56] = 9'b111111111;
assign micromatri[42][57] = 9'b111111111;
assign micromatri[42][58] = 9'b111111111;
assign micromatri[42][59] = 9'b111111111;
assign micromatri[42][60] = 9'b111111111;
assign micromatri[42][61] = 9'b111111111;
assign micromatri[42][62] = 9'b111111111;
assign micromatri[42][63] = 9'b111111111;
assign micromatri[42][64] = 9'b111111111;
assign micromatri[42][65] = 9'b111111111;
assign micromatri[42][66] = 9'b111111111;
assign micromatri[42][67] = 9'b111111111;
assign micromatri[42][68] = 9'b111111111;
assign micromatri[42][69] = 9'b111111111;
assign micromatri[42][70] = 9'b111111111;
assign micromatri[42][71] = 9'b111111111;
assign micromatri[42][72] = 9'b111111111;
assign micromatri[42][73] = 9'b111111111;
assign micromatri[42][74] = 9'b111111111;
assign micromatri[42][75] = 9'b111111111;
assign micromatri[42][76] = 9'b111111111;
assign micromatri[42][77] = 9'b111111111;
assign micromatri[42][78] = 9'b111111111;
assign micromatri[42][79] = 9'b111111111;
assign micromatri[42][80] = 9'b111111111;
assign micromatri[42][81] = 9'b111111111;
assign micromatri[42][82] = 9'b111111111;
assign micromatri[42][83] = 9'b111111111;
assign micromatri[42][84] = 9'b111111111;
assign micromatri[42][85] = 9'b111111111;
assign micromatri[42][86] = 9'b111111111;
assign micromatri[42][87] = 9'b111111111;
assign micromatri[42][88] = 9'b111111111;
assign micromatri[42][89] = 9'b111111111;
assign micromatri[42][90] = 9'b111111111;
assign micromatri[42][91] = 9'b111111111;
assign micromatri[42][92] = 9'b111111111;
assign micromatri[42][93] = 9'b111111111;
assign micromatri[42][94] = 9'b111111111;
assign micromatri[42][95] = 9'b111111111;
assign micromatri[42][96] = 9'b111111111;
assign micromatri[42][97] = 9'b111111111;
assign micromatri[42][98] = 9'b111111111;
assign micromatri[42][99] = 9'b111111111;
assign micromatri[43][0] = 9'b111111111;
assign micromatri[43][1] = 9'b111111111;
assign micromatri[43][2] = 9'b111111111;
assign micromatri[43][3] = 9'b111111111;
assign micromatri[43][4] = 9'b111111111;
assign micromatri[43][5] = 9'b111111111;
assign micromatri[43][6] = 9'b111111111;
assign micromatri[43][7] = 9'b111111111;
assign micromatri[43][8] = 9'b111111111;
assign micromatri[43][9] = 9'b111111111;
assign micromatri[43][10] = 9'b111111111;
assign micromatri[43][11] = 9'b111111111;
assign micromatri[43][12] = 9'b111111111;
assign micromatri[43][13] = 9'b111111111;
assign micromatri[43][14] = 9'b111111111;
assign micromatri[43][15] = 9'b111111111;
assign micromatri[43][16] = 9'b111111111;
assign micromatri[43][17] = 9'b111111111;
assign micromatri[43][18] = 9'b111111111;
assign micromatri[43][19] = 9'b111111111;
assign micromatri[43][20] = 9'b111111111;
assign micromatri[43][21] = 9'b111111111;
assign micromatri[43][22] = 9'b111111111;
assign micromatri[43][23] = 9'b111111111;
assign micromatri[43][24] = 9'b111111111;
assign micromatri[43][25] = 9'b111111111;
assign micromatri[43][26] = 9'b111111111;
assign micromatri[43][27] = 9'b111111111;
assign micromatri[43][28] = 9'b111111111;
assign micromatri[43][29] = 9'b111111111;
assign micromatri[43][30] = 9'b111111111;
assign micromatri[43][31] = 9'b111111111;
assign micromatri[43][32] = 9'b111111111;
assign micromatri[43][33] = 9'b111111111;
assign micromatri[43][34] = 9'b111111111;
assign micromatri[43][35] = 9'b111111111;
assign micromatri[43][36] = 9'b111111111;
assign micromatri[43][37] = 9'b111111111;
assign micromatri[43][38] = 9'b111111111;
assign micromatri[43][39] = 9'b111111111;
assign micromatri[43][40] = 9'b111111111;
assign micromatri[43][41] = 9'b111111111;
assign micromatri[43][42] = 9'b111111111;
assign micromatri[43][43] = 9'b111111111;
assign micromatri[43][44] = 9'b111111111;
assign micromatri[43][45] = 9'b111111111;
assign micromatri[43][46] = 9'b111111111;
assign micromatri[43][47] = 9'b111111111;
assign micromatri[43][48] = 9'b111111111;
assign micromatri[43][49] = 9'b111111111;
assign micromatri[43][50] = 9'b111111111;
assign micromatri[43][51] = 9'b111111111;
assign micromatri[43][52] = 9'b111111111;
assign micromatri[43][53] = 9'b111111111;
assign micromatri[43][54] = 9'b111111111;
assign micromatri[43][55] = 9'b111111111;
assign micromatri[43][56] = 9'b111111111;
assign micromatri[43][57] = 9'b111111111;
assign micromatri[43][58] = 9'b111111111;
assign micromatri[43][59] = 9'b111111111;
assign micromatri[43][60] = 9'b111111111;
assign micromatri[43][61] = 9'b111111111;
assign micromatri[43][62] = 9'b111111111;
assign micromatri[43][63] = 9'b111111111;
assign micromatri[43][64] = 9'b111111111;
assign micromatri[43][65] = 9'b111111111;
assign micromatri[43][66] = 9'b111111111;
assign micromatri[43][67] = 9'b111111111;
assign micromatri[43][68] = 9'b111111111;
assign micromatri[43][69] = 9'b111111111;
assign micromatri[43][70] = 9'b111111111;
assign micromatri[43][71] = 9'b111111111;
assign micromatri[43][72] = 9'b111111111;
assign micromatri[43][73] = 9'b111111111;
assign micromatri[43][74] = 9'b111111111;
assign micromatri[43][75] = 9'b111111111;
assign micromatri[43][76] = 9'b111111111;
assign micromatri[43][77] = 9'b111111111;
assign micromatri[43][78] = 9'b111111111;
assign micromatri[43][79] = 9'b111111111;
assign micromatri[43][80] = 9'b111111111;
assign micromatri[43][81] = 9'b111111111;
assign micromatri[43][82] = 9'b111111111;
assign micromatri[43][83] = 9'b111111111;
assign micromatri[43][84] = 9'b111111111;
assign micromatri[43][85] = 9'b111111111;
assign micromatri[43][86] = 9'b111111111;
assign micromatri[43][87] = 9'b111111111;
assign micromatri[43][88] = 9'b111111111;
assign micromatri[43][89] = 9'b111111111;
assign micromatri[43][90] = 9'b111111111;
assign micromatri[43][91] = 9'b111111111;
assign micromatri[43][92] = 9'b111111111;
assign micromatri[43][93] = 9'b111111111;
assign micromatri[43][94] = 9'b111111111;
assign micromatri[43][95] = 9'b111111111;
assign micromatri[43][96] = 9'b111111111;
assign micromatri[43][97] = 9'b111111111;
assign micromatri[43][98] = 9'b111111111;
assign micromatri[43][99] = 9'b111111111;
assign micromatri[44][0] = 9'b111111111;
assign micromatri[44][1] = 9'b111111111;
assign micromatri[44][2] = 9'b111111111;
assign micromatri[44][3] = 9'b111111111;
assign micromatri[44][4] = 9'b111111111;
assign micromatri[44][5] = 9'b111111111;
assign micromatri[44][6] = 9'b111111111;
assign micromatri[44][7] = 9'b111111111;
assign micromatri[44][8] = 9'b111111111;
assign micromatri[44][9] = 9'b111111111;
assign micromatri[44][10] = 9'b111111111;
assign micromatri[44][11] = 9'b111111111;
assign micromatri[44][12] = 9'b111111111;
assign micromatri[44][13] = 9'b111111111;
assign micromatri[44][14] = 9'b111111111;
assign micromatri[44][15] = 9'b111111111;
assign micromatri[44][16] = 9'b111111111;
assign micromatri[44][17] = 9'b111111111;
assign micromatri[44][18] = 9'b111111111;
assign micromatri[44][19] = 9'b111111111;
assign micromatri[44][20] = 9'b111111111;
assign micromatri[44][21] = 9'b111111111;
assign micromatri[44][22] = 9'b111111111;
assign micromatri[44][23] = 9'b111111111;
assign micromatri[44][24] = 9'b111111111;
assign micromatri[44][25] = 9'b111111111;
assign micromatri[44][26] = 9'b111111111;
assign micromatri[44][27] = 9'b111111111;
assign micromatri[44][28] = 9'b111111111;
assign micromatri[44][29] = 9'b111111111;
assign micromatri[44][30] = 9'b111111111;
assign micromatri[44][31] = 9'b111111111;
assign micromatri[44][32] = 9'b111111111;
assign micromatri[44][33] = 9'b111111111;
assign micromatri[44][34] = 9'b111111111;
assign micromatri[44][35] = 9'b111111111;
assign micromatri[44][36] = 9'b111111111;
assign micromatri[44][37] = 9'b111111111;
assign micromatri[44][38] = 9'b111111111;
assign micromatri[44][39] = 9'b111111111;
assign micromatri[44][40] = 9'b111111111;
assign micromatri[44][41] = 9'b111111111;
assign micromatri[44][42] = 9'b111111111;
assign micromatri[44][43] = 9'b111111111;
assign micromatri[44][44] = 9'b111111111;
assign micromatri[44][45] = 9'b111111111;
assign micromatri[44][46] = 9'b111111111;
assign micromatri[44][47] = 9'b111111111;
assign micromatri[44][48] = 9'b111111111;
assign micromatri[44][49] = 9'b111111111;
assign micromatri[44][50] = 9'b111111111;
assign micromatri[44][51] = 9'b111111111;
assign micromatri[44][52] = 9'b111111111;
assign micromatri[44][53] = 9'b111111111;
assign micromatri[44][54] = 9'b111111111;
assign micromatri[44][55] = 9'b111111111;
assign micromatri[44][56] = 9'b111111111;
assign micromatri[44][57] = 9'b111111111;
assign micromatri[44][58] = 9'b111111111;
assign micromatri[44][59] = 9'b111111111;
assign micromatri[44][60] = 9'b111111111;
assign micromatri[44][61] = 9'b111111111;
assign micromatri[44][62] = 9'b111111111;
assign micromatri[44][63] = 9'b111111111;
assign micromatri[44][64] = 9'b111111111;
assign micromatri[44][65] = 9'b111111111;
assign micromatri[44][66] = 9'b111111111;
assign micromatri[44][67] = 9'b111111111;
assign micromatri[44][68] = 9'b111111111;
assign micromatri[44][69] = 9'b111111111;
assign micromatri[44][70] = 9'b111111111;
assign micromatri[44][71] = 9'b111111111;
assign micromatri[44][72] = 9'b111111111;
assign micromatri[44][73] = 9'b111111111;
assign micromatri[44][74] = 9'b111111111;
assign micromatri[44][75] = 9'b111111111;
assign micromatri[44][76] = 9'b111111111;
assign micromatri[44][77] = 9'b111111111;
assign micromatri[44][78] = 9'b111111111;
assign micromatri[44][79] = 9'b111111111;
assign micromatri[44][80] = 9'b111111111;
assign micromatri[44][81] = 9'b111111111;
assign micromatri[44][82] = 9'b111111111;
assign micromatri[44][83] = 9'b111111111;
assign micromatri[44][84] = 9'b111111111;
assign micromatri[44][85] = 9'b111111111;
assign micromatri[44][86] = 9'b111111111;
assign micromatri[44][87] = 9'b111111111;
assign micromatri[44][88] = 9'b111111111;
assign micromatri[44][89] = 9'b111111111;
assign micromatri[44][90] = 9'b111111111;
assign micromatri[44][91] = 9'b111111111;
assign micromatri[44][92] = 9'b111111111;
assign micromatri[44][93] = 9'b111111111;
assign micromatri[44][94] = 9'b111111111;
assign micromatri[44][95] = 9'b111111111;
assign micromatri[44][96] = 9'b111111111;
assign micromatri[44][97] = 9'b111111111;
assign micromatri[44][98] = 9'b111111111;
assign micromatri[44][99] = 9'b111111111;
assign micromatri[45][0] = 9'b111111111;
assign micromatri[45][1] = 9'b111111111;
assign micromatri[45][2] = 9'b111111111;
assign micromatri[45][3] = 9'b111111111;
assign micromatri[45][4] = 9'b111111111;
assign micromatri[45][5] = 9'b111111111;
assign micromatri[45][6] = 9'b111111111;
assign micromatri[45][7] = 9'b111111111;
assign micromatri[45][8] = 9'b111111111;
assign micromatri[45][9] = 9'b111111111;
assign micromatri[45][10] = 9'b111111111;
assign micromatri[45][11] = 9'b111111111;
assign micromatri[45][12] = 9'b111111111;
assign micromatri[45][13] = 9'b111111111;
assign micromatri[45][14] = 9'b111111111;
assign micromatri[45][15] = 9'b111111111;
assign micromatri[45][16] = 9'b111111111;
assign micromatri[45][17] = 9'b111111111;
assign micromatri[45][18] = 9'b111111111;
assign micromatri[45][19] = 9'b111111111;
assign micromatri[45][20] = 9'b111111111;
assign micromatri[45][21] = 9'b111111111;
assign micromatri[45][22] = 9'b111111111;
assign micromatri[45][23] = 9'b111111111;
assign micromatri[45][24] = 9'b111111111;
assign micromatri[45][25] = 9'b111111111;
assign micromatri[45][26] = 9'b111111111;
assign micromatri[45][27] = 9'b111111111;
assign micromatri[45][28] = 9'b111111111;
assign micromatri[45][29] = 9'b111111111;
assign micromatri[45][30] = 9'b111111111;
assign micromatri[45][31] = 9'b111111111;
assign micromatri[45][32] = 9'b111111111;
assign micromatri[45][33] = 9'b111111111;
assign micromatri[45][34] = 9'b111111111;
assign micromatri[45][35] = 9'b111111111;
assign micromatri[45][36] = 9'b111111111;
assign micromatri[45][37] = 9'b111111111;
assign micromatri[45][38] = 9'b111111111;
assign micromatri[45][39] = 9'b111111111;
assign micromatri[45][40] = 9'b111111111;
assign micromatri[45][41] = 9'b111111111;
assign micromatri[45][42] = 9'b111111111;
assign micromatri[45][43] = 9'b111111111;
assign micromatri[45][44] = 9'b111111111;
assign micromatri[45][45] = 9'b111111111;
assign micromatri[45][46] = 9'b111111111;
assign micromatri[45][47] = 9'b111111111;
assign micromatri[45][48] = 9'b111111111;
assign micromatri[45][49] = 9'b111111111;
assign micromatri[45][50] = 9'b111111111;
assign micromatri[45][51] = 9'b111111111;
assign micromatri[45][52] = 9'b111111111;
assign micromatri[45][53] = 9'b111111111;
assign micromatri[45][54] = 9'b111111111;
assign micromatri[45][55] = 9'b111111111;
assign micromatri[45][56] = 9'b111111111;
assign micromatri[45][57] = 9'b111111111;
assign micromatri[45][58] = 9'b111111111;
assign micromatri[45][59] = 9'b111111111;
assign micromatri[45][60] = 9'b111111111;
assign micromatri[45][61] = 9'b111111111;
assign micromatri[45][62] = 9'b111111111;
assign micromatri[45][63] = 9'b111111111;
assign micromatri[45][64] = 9'b111111111;
assign micromatri[45][65] = 9'b111111111;
assign micromatri[45][66] = 9'b111111111;
assign micromatri[45][67] = 9'b111111111;
assign micromatri[45][68] = 9'b111111111;
assign micromatri[45][69] = 9'b111111111;
assign micromatri[45][70] = 9'b111111111;
assign micromatri[45][71] = 9'b111111111;
assign micromatri[45][72] = 9'b111111111;
assign micromatri[45][73] = 9'b111111111;
assign micromatri[45][74] = 9'b111111111;
assign micromatri[45][75] = 9'b111111111;
assign micromatri[45][76] = 9'b111111111;
assign micromatri[45][77] = 9'b111111111;
assign micromatri[45][78] = 9'b111111111;
assign micromatri[45][79] = 9'b111111111;
assign micromatri[45][80] = 9'b111111111;
assign micromatri[45][81] = 9'b111111111;
assign micromatri[45][82] = 9'b111111111;
assign micromatri[45][83] = 9'b111111111;
assign micromatri[45][84] = 9'b111111111;
assign micromatri[45][85] = 9'b111111111;
assign micromatri[45][86] = 9'b111111111;
assign micromatri[45][87] = 9'b111111111;
assign micromatri[45][88] = 9'b111111111;
assign micromatri[45][89] = 9'b111111111;
assign micromatri[45][90] = 9'b111111111;
assign micromatri[45][91] = 9'b111111111;
assign micromatri[45][92] = 9'b111111111;
assign micromatri[45][93] = 9'b111111111;
assign micromatri[45][94] = 9'b111111111;
assign micromatri[45][95] = 9'b111111111;
assign micromatri[45][96] = 9'b111111111;
assign micromatri[45][97] = 9'b111111111;
assign micromatri[45][98] = 9'b111111111;
assign micromatri[45][99] = 9'b111111111;
assign micromatri[46][0] = 9'b111111111;
assign micromatri[46][1] = 9'b111111111;
assign micromatri[46][2] = 9'b111111111;
assign micromatri[46][3] = 9'b111111111;
assign micromatri[46][4] = 9'b111111111;
assign micromatri[46][5] = 9'b111111111;
assign micromatri[46][6] = 9'b111111111;
assign micromatri[46][7] = 9'b111111111;
assign micromatri[46][8] = 9'b111111111;
assign micromatri[46][9] = 9'b111111111;
assign micromatri[46][10] = 9'b111111111;
assign micromatri[46][11] = 9'b111111111;
assign micromatri[46][12] = 9'b111111111;
assign micromatri[46][13] = 9'b111111111;
assign micromatri[46][14] = 9'b111111111;
assign micromatri[46][15] = 9'b111111111;
assign micromatri[46][16] = 9'b111111111;
assign micromatri[46][17] = 9'b111111111;
assign micromatri[46][18] = 9'b111111111;
assign micromatri[46][19] = 9'b111111111;
assign micromatri[46][20] = 9'b111111111;
assign micromatri[46][21] = 9'b111111111;
assign micromatri[46][22] = 9'b111111111;
assign micromatri[46][23] = 9'b111111111;
assign micromatri[46][24] = 9'b111111111;
assign micromatri[46][25] = 9'b111111111;
assign micromatri[46][26] = 9'b111111111;
assign micromatri[46][27] = 9'b111111111;
assign micromatri[46][28] = 9'b111111111;
assign micromatri[46][29] = 9'b111111111;
assign micromatri[46][30] = 9'b111111111;
assign micromatri[46][31] = 9'b111111111;
assign micromatri[46][32] = 9'b111111111;
assign micromatri[46][33] = 9'b111111111;
assign micromatri[46][34] = 9'b111111111;
assign micromatri[46][35] = 9'b111111111;
assign micromatri[46][36] = 9'b111111111;
assign micromatri[46][37] = 9'b111111111;
assign micromatri[46][38] = 9'b111111111;
assign micromatri[46][39] = 9'b111111111;
assign micromatri[46][40] = 9'b111111111;
assign micromatri[46][41] = 9'b111111111;
assign micromatri[46][42] = 9'b111111111;
assign micromatri[46][43] = 9'b111111111;
assign micromatri[46][44] = 9'b111111111;
assign micromatri[46][45] = 9'b111111111;
assign micromatri[46][46] = 9'b111111111;
assign micromatri[46][47] = 9'b111111111;
assign micromatri[46][48] = 9'b111111111;
assign micromatri[46][49] = 9'b111111111;
assign micromatri[46][50] = 9'b111111111;
assign micromatri[46][51] = 9'b111111111;
assign micromatri[46][52] = 9'b111111111;
assign micromatri[46][53] = 9'b111111111;
assign micromatri[46][54] = 9'b111111111;
assign micromatri[46][55] = 9'b111111111;
assign micromatri[46][56] = 9'b111111111;
assign micromatri[46][57] = 9'b111111111;
assign micromatri[46][58] = 9'b111111111;
assign micromatri[46][59] = 9'b111111111;
assign micromatri[46][60] = 9'b111111111;
assign micromatri[46][61] = 9'b111111111;
assign micromatri[46][62] = 9'b111111111;
assign micromatri[46][63] = 9'b111111111;
assign micromatri[46][64] = 9'b111111111;
assign micromatri[46][65] = 9'b111111111;
assign micromatri[46][66] = 9'b111111111;
assign micromatri[46][67] = 9'b111111111;
assign micromatri[46][68] = 9'b111111111;
assign micromatri[46][69] = 9'b111111111;
assign micromatri[46][70] = 9'b111111111;
assign micromatri[46][71] = 9'b111111111;
assign micromatri[46][72] = 9'b111111111;
assign micromatri[46][73] = 9'b111111111;
assign micromatri[46][74] = 9'b111111111;
assign micromatri[46][75] = 9'b111111111;
assign micromatri[46][76] = 9'b111111111;
assign micromatri[46][77] = 9'b111111111;
assign micromatri[46][78] = 9'b111111111;
assign micromatri[46][79] = 9'b111111111;
assign micromatri[46][80] = 9'b111111111;
assign micromatri[46][81] = 9'b111111111;
assign micromatri[46][82] = 9'b111111111;
assign micromatri[46][83] = 9'b111111111;
assign micromatri[46][84] = 9'b111111111;
assign micromatri[46][85] = 9'b111111111;
assign micromatri[46][86] = 9'b111111111;
assign micromatri[46][87] = 9'b111111111;
assign micromatri[46][88] = 9'b111111111;
assign micromatri[46][89] = 9'b111111111;
assign micromatri[46][90] = 9'b111111111;
assign micromatri[46][91] = 9'b111111111;
assign micromatri[46][92] = 9'b111111111;
assign micromatri[46][93] = 9'b111111111;
assign micromatri[46][94] = 9'b111111111;
assign micromatri[46][95] = 9'b111111111;
assign micromatri[46][96] = 9'b111111111;
assign micromatri[46][97] = 9'b111111111;
assign micromatri[46][98] = 9'b111111111;
assign micromatri[46][99] = 9'b111111111;
assign micromatri[47][0] = 9'b111111111;
assign micromatri[47][1] = 9'b111111111;
assign micromatri[47][2] = 9'b111111111;
assign micromatri[47][3] = 9'b111111111;
assign micromatri[47][4] = 9'b111111111;
assign micromatri[47][5] = 9'b111111111;
assign micromatri[47][6] = 9'b111111111;
assign micromatri[47][7] = 9'b111111111;
assign micromatri[47][8] = 9'b111111111;
assign micromatri[47][9] = 9'b111111111;
assign micromatri[47][10] = 9'b111111111;
assign micromatri[47][11] = 9'b111111111;
assign micromatri[47][12] = 9'b111111111;
assign micromatri[47][13] = 9'b111111111;
assign micromatri[47][14] = 9'b111111111;
assign micromatri[47][15] = 9'b111111111;
assign micromatri[47][16] = 9'b111111111;
assign micromatri[47][17] = 9'b111111111;
assign micromatri[47][18] = 9'b111111111;
assign micromatri[47][19] = 9'b111111111;
assign micromatri[47][20] = 9'b111111111;
assign micromatri[47][21] = 9'b111111111;
assign micromatri[47][22] = 9'b111111111;
assign micromatri[47][23] = 9'b111111111;
assign micromatri[47][24] = 9'b111111111;
assign micromatri[47][25] = 9'b111111111;
assign micromatri[47][26] = 9'b111111111;
assign micromatri[47][27] = 9'b111111111;
assign micromatri[47][28] = 9'b111111111;
assign micromatri[47][29] = 9'b111111111;
assign micromatri[47][30] = 9'b111111111;
assign micromatri[47][31] = 9'b111111111;
assign micromatri[47][32] = 9'b111111111;
assign micromatri[47][33] = 9'b111111111;
assign micromatri[47][34] = 9'b111111111;
assign micromatri[47][35] = 9'b111111111;
assign micromatri[47][36] = 9'b111111111;
assign micromatri[47][37] = 9'b111111111;
assign micromatri[47][38] = 9'b111111111;
assign micromatri[47][39] = 9'b111111111;
assign micromatri[47][40] = 9'b111111111;
assign micromatri[47][41] = 9'b111111111;
assign micromatri[47][42] = 9'b111111111;
assign micromatri[47][43] = 9'b111111111;
assign micromatri[47][44] = 9'b111111111;
assign micromatri[47][45] = 9'b111111111;
assign micromatri[47][46] = 9'b111111111;
assign micromatri[47][47] = 9'b111111111;
assign micromatri[47][48] = 9'b111111111;
assign micromatri[47][49] = 9'b111111111;
assign micromatri[47][50] = 9'b111111111;
assign micromatri[47][51] = 9'b111111111;
assign micromatri[47][52] = 9'b111111111;
assign micromatri[47][53] = 9'b111111111;
assign micromatri[47][54] = 9'b111111111;
assign micromatri[47][55] = 9'b111111111;
assign micromatri[47][56] = 9'b111111111;
assign micromatri[47][57] = 9'b111111111;
assign micromatri[47][58] = 9'b111111111;
assign micromatri[47][59] = 9'b111111111;
assign micromatri[47][60] = 9'b111111111;
assign micromatri[47][61] = 9'b111111111;
assign micromatri[47][62] = 9'b111111111;
assign micromatri[47][63] = 9'b111111111;
assign micromatri[47][64] = 9'b111111111;
assign micromatri[47][65] = 9'b111111111;
assign micromatri[47][66] = 9'b111111111;
assign micromatri[47][67] = 9'b111111111;
assign micromatri[47][68] = 9'b111111111;
assign micromatri[47][69] = 9'b111111111;
assign micromatri[47][70] = 9'b111111111;
assign micromatri[47][71] = 9'b111111111;
assign micromatri[47][72] = 9'b111111111;
assign micromatri[47][73] = 9'b111111111;
assign micromatri[47][74] = 9'b111111111;
assign micromatri[47][75] = 9'b111111111;
assign micromatri[47][76] = 9'b111111111;
assign micromatri[47][77] = 9'b111111111;
assign micromatri[47][78] = 9'b111111111;
assign micromatri[47][79] = 9'b111111111;
assign micromatri[47][80] = 9'b111111111;
assign micromatri[47][81] = 9'b111111111;
assign micromatri[47][82] = 9'b111111111;
assign micromatri[47][83] = 9'b111111111;
assign micromatri[47][84] = 9'b111111111;
assign micromatri[47][85] = 9'b111111111;
assign micromatri[47][86] = 9'b111111111;
assign micromatri[47][87] = 9'b111111111;
assign micromatri[47][88] = 9'b111111111;
assign micromatri[47][89] = 9'b111111111;
assign micromatri[47][90] = 9'b111111111;
assign micromatri[47][91] = 9'b111111111;
assign micromatri[47][92] = 9'b111111111;
assign micromatri[47][93] = 9'b111111111;
assign micromatri[47][94] = 9'b111111111;
assign micromatri[47][95] = 9'b111111111;
assign micromatri[47][96] = 9'b111111111;
assign micromatri[47][97] = 9'b111111111;
assign micromatri[47][98] = 9'b111111111;
assign micromatri[47][99] = 9'b111111111;
assign micromatri[48][0] = 9'b111111111;
assign micromatri[48][1] = 9'b111111111;
assign micromatri[48][2] = 9'b111111111;
assign micromatri[48][3] = 9'b111111111;
assign micromatri[48][4] = 9'b111111111;
assign micromatri[48][5] = 9'b111111111;
assign micromatri[48][6] = 9'b111111111;
assign micromatri[48][7] = 9'b111111111;
assign micromatri[48][8] = 9'b111111111;
assign micromatri[48][9] = 9'b111111111;
assign micromatri[48][10] = 9'b111111111;
assign micromatri[48][11] = 9'b111111111;
assign micromatri[48][12] = 9'b111111111;
assign micromatri[48][13] = 9'b111111111;
assign micromatri[48][14] = 9'b111111111;
assign micromatri[48][15] = 9'b111111111;
assign micromatri[48][16] = 9'b111111111;
assign micromatri[48][17] = 9'b111111111;
assign micromatri[48][18] = 9'b111111111;
assign micromatri[48][19] = 9'b111111111;
assign micromatri[48][20] = 9'b111111111;
assign micromatri[48][21] = 9'b111111111;
assign micromatri[48][22] = 9'b111111111;
assign micromatri[48][23] = 9'b111111111;
assign micromatri[48][24] = 9'b111111111;
assign micromatri[48][25] = 9'b111111111;
assign micromatri[48][26] = 9'b111111111;
assign micromatri[48][27] = 9'b111111111;
assign micromatri[48][28] = 9'b111111111;
assign micromatri[48][29] = 9'b111111111;
assign micromatri[48][30] = 9'b111111111;
assign micromatri[48][31] = 9'b111111111;
assign micromatri[48][32] = 9'b111111111;
assign micromatri[48][33] = 9'b111111111;
assign micromatri[48][34] = 9'b111111111;
assign micromatri[48][35] = 9'b111111111;
assign micromatri[48][36] = 9'b111111111;
assign micromatri[48][37] = 9'b111111111;
assign micromatri[48][38] = 9'b111111111;
assign micromatri[48][39] = 9'b111111111;
assign micromatri[48][40] = 9'b111111111;
assign micromatri[48][41] = 9'b111111111;
assign micromatri[48][42] = 9'b111111111;
assign micromatri[48][43] = 9'b111111111;
assign micromatri[48][44] = 9'b111111111;
assign micromatri[48][45] = 9'b111111111;
assign micromatri[48][46] = 9'b111111111;
assign micromatri[48][47] = 9'b111111111;
assign micromatri[48][48] = 9'b111111111;
assign micromatri[48][49] = 9'b111111111;
assign micromatri[48][50] = 9'b111111111;
assign micromatri[48][51] = 9'b111111111;
assign micromatri[48][52] = 9'b111111111;
assign micromatri[48][53] = 9'b111111111;
assign micromatri[48][54] = 9'b111111111;
assign micromatri[48][55] = 9'b111111111;
assign micromatri[48][56] = 9'b111111111;
assign micromatri[48][57] = 9'b111111111;
assign micromatri[48][58] = 9'b111111111;
assign micromatri[48][59] = 9'b111111111;
assign micromatri[48][60] = 9'b111111111;
assign micromatri[48][61] = 9'b111111111;
assign micromatri[48][62] = 9'b111111111;
assign micromatri[48][63] = 9'b111111111;
assign micromatri[48][64] = 9'b111111111;
assign micromatri[48][65] = 9'b111111111;
assign micromatri[48][66] = 9'b111111111;
assign micromatri[48][67] = 9'b111111111;
assign micromatri[48][68] = 9'b111111111;
assign micromatri[48][69] = 9'b111111111;
assign micromatri[48][70] = 9'b111111111;
assign micromatri[48][71] = 9'b111111111;
assign micromatri[48][72] = 9'b111111111;
assign micromatri[48][73] = 9'b111111111;
assign micromatri[48][74] = 9'b111111111;
assign micromatri[48][75] = 9'b111111111;
assign micromatri[48][76] = 9'b111111111;
assign micromatri[48][77] = 9'b111111111;
assign micromatri[48][78] = 9'b111111111;
assign micromatri[48][79] = 9'b111111111;
assign micromatri[48][80] = 9'b111111111;
assign micromatri[48][81] = 9'b111111111;
assign micromatri[48][82] = 9'b111111111;
assign micromatri[48][83] = 9'b111111111;
assign micromatri[48][84] = 9'b111111111;
assign micromatri[48][85] = 9'b111111111;
assign micromatri[48][86] = 9'b111111111;
assign micromatri[48][87] = 9'b111111111;
assign micromatri[48][88] = 9'b111111111;
assign micromatri[48][89] = 9'b111111111;
assign micromatri[48][90] = 9'b111111111;
assign micromatri[48][91] = 9'b111111111;
assign micromatri[48][92] = 9'b111111111;
assign micromatri[48][93] = 9'b111111111;
assign micromatri[48][94] = 9'b111111111;
assign micromatri[48][95] = 9'b111111111;
assign micromatri[48][96] = 9'b111111111;
assign micromatri[48][97] = 9'b111111111;
assign micromatri[48][98] = 9'b111111111;
assign micromatri[48][99] = 9'b111111111;
assign micromatri[49][0] = 9'b111111111;
assign micromatri[49][1] = 9'b111111111;
assign micromatri[49][2] = 9'b111111111;
assign micromatri[49][3] = 9'b111111111;
assign micromatri[49][4] = 9'b111111111;
assign micromatri[49][5] = 9'b111111111;
assign micromatri[49][6] = 9'b111111111;
assign micromatri[49][7] = 9'b111111111;
assign micromatri[49][8] = 9'b111111111;
assign micromatri[49][9] = 9'b111111111;
assign micromatri[49][10] = 9'b111111111;
assign micromatri[49][11] = 9'b111111111;
assign micromatri[49][12] = 9'b111111111;
assign micromatri[49][13] = 9'b111111111;
assign micromatri[49][14] = 9'b111111111;
assign micromatri[49][15] = 9'b111111111;
assign micromatri[49][16] = 9'b111111111;
assign micromatri[49][17] = 9'b111111111;
assign micromatri[49][18] = 9'b111111111;
assign micromatri[49][19] = 9'b111111111;
assign micromatri[49][20] = 9'b111111111;
assign micromatri[49][21] = 9'b111111111;
assign micromatri[49][22] = 9'b111111111;
assign micromatri[49][23] = 9'b111111111;
assign micromatri[49][24] = 9'b111111111;
assign micromatri[49][25] = 9'b111111111;
assign micromatri[49][26] = 9'b111111111;
assign micromatri[49][27] = 9'b111111111;
assign micromatri[49][28] = 9'b111111111;
assign micromatri[49][29] = 9'b111111111;
assign micromatri[49][30] = 9'b111111111;
assign micromatri[49][31] = 9'b111111111;
assign micromatri[49][32] = 9'b111111111;
assign micromatri[49][33] = 9'b111111111;
assign micromatri[49][34] = 9'b111111111;
assign micromatri[49][35] = 9'b111111111;
assign micromatri[49][36] = 9'b111111111;
assign micromatri[49][37] = 9'b111111111;
assign micromatri[49][38] = 9'b111111111;
assign micromatri[49][39] = 9'b111111111;
assign micromatri[49][40] = 9'b111111111;
assign micromatri[49][41] = 9'b111111111;
assign micromatri[49][42] = 9'b111111111;
assign micromatri[49][43] = 9'b111111111;
assign micromatri[49][44] = 9'b111111111;
assign micromatri[49][45] = 9'b111111111;
assign micromatri[49][46] = 9'b111111111;
assign micromatri[49][47] = 9'b111111111;
assign micromatri[49][48] = 9'b111111111;
assign micromatri[49][49] = 9'b111111111;
assign micromatri[49][50] = 9'b111111111;
assign micromatri[49][51] = 9'b111111111;
assign micromatri[49][52] = 9'b111111111;
assign micromatri[49][53] = 9'b111111111;
assign micromatri[49][54] = 9'b111111111;
assign micromatri[49][55] = 9'b111111111;
assign micromatri[49][56] = 9'b111111111;
assign micromatri[49][57] = 9'b111111111;
assign micromatri[49][58] = 9'b111111111;
assign micromatri[49][59] = 9'b111111111;
assign micromatri[49][60] = 9'b111111111;
assign micromatri[49][61] = 9'b111111111;
assign micromatri[49][62] = 9'b111111111;
assign micromatri[49][63] = 9'b111111111;
assign micromatri[49][64] = 9'b111111111;
assign micromatri[49][65] = 9'b111111111;
assign micromatri[49][66] = 9'b111111111;
assign micromatri[49][67] = 9'b111111111;
assign micromatri[49][68] = 9'b111111111;
assign micromatri[49][69] = 9'b111111111;
assign micromatri[49][70] = 9'b111111111;
assign micromatri[49][71] = 9'b111111111;
assign micromatri[49][72] = 9'b111111111;
assign micromatri[49][73] = 9'b111111111;
assign micromatri[49][74] = 9'b111111111;
assign micromatri[49][75] = 9'b111111111;
assign micromatri[49][76] = 9'b111111111;
assign micromatri[49][77] = 9'b111111111;
assign micromatri[49][78] = 9'b111111111;
assign micromatri[49][79] = 9'b111111111;
assign micromatri[49][80] = 9'b111111111;
assign micromatri[49][81] = 9'b111111111;
assign micromatri[49][82] = 9'b111111111;
assign micromatri[49][83] = 9'b111111111;
assign micromatri[49][84] = 9'b111111111;
assign micromatri[49][85] = 9'b111111111;
assign micromatri[49][86] = 9'b111111111;
assign micromatri[49][87] = 9'b111111111;
assign micromatri[49][88] = 9'b111111111;
assign micromatri[49][89] = 9'b111111111;
assign micromatri[49][90] = 9'b111111111;
assign micromatri[49][91] = 9'b111111111;
assign micromatri[49][92] = 9'b111111111;
assign micromatri[49][93] = 9'b111111111;
assign micromatri[49][94] = 9'b111111111;
assign micromatri[49][95] = 9'b111111111;
assign micromatri[49][96] = 9'b111111111;
assign micromatri[49][97] = 9'b111111111;
assign micromatri[49][98] = 9'b111111111;
assign micromatri[49][99] = 9'b111111111;
//Total de Lineas = 5000
endmodule



