`timescale 1ns / 1ps
module seleccion_alonzo (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (F[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= F[vcount- posy][hcount- posx][7:5];
				green <= F[vcount- posy][hcount- posx][4:2];
            blue 	<= F[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 64;
parameter RESOLUCION_Y = 64;
wire [8:0] F[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign F[5][29] = 9'b111111111;
assign F[5][30] = 9'b111111111;
assign F[5][31] = 9'b111111111;
assign F[5][32] = 9'b111111111;
assign F[5][33] = 9'b111111111;
assign F[5][34] = 9'b111111111;
assign F[6][27] = 9'b111111111;
assign F[6][28] = 9'b111111111;
assign F[6][29] = 9'b111111111;
assign F[6][30] = 9'b111111111;
assign F[6][31] = 9'b111111111;
assign F[6][32] = 9'b111111111;
assign F[6][33] = 9'b111111111;
assign F[6][34] = 9'b111111111;
assign F[6][35] = 9'b111111111;
assign F[6][36] = 9'b111111111;
assign F[7][26] = 9'b111111111;
assign F[7][27] = 9'b111111111;
assign F[7][28] = 9'b111111111;
assign F[7][29] = 9'b110010010;
assign F[7][30] = 9'b101101110;
assign F[7][31] = 9'b101101110;
assign F[7][32] = 9'b101101110;
assign F[7][33] = 9'b101101110;
assign F[7][34] = 9'b110010011;
assign F[7][35] = 9'b111111111;
assign F[7][36] = 9'b111111111;
assign F[7][37] = 9'b111111111;
assign F[8][25] = 9'b111111111;
assign F[8][26] = 9'b111111111;
assign F[8][27] = 9'b111111110;
assign F[8][28] = 9'b101101001;
assign F[8][29] = 9'b100100001;
assign F[8][30] = 9'b101101010;
assign F[8][31] = 9'b101101010;
assign F[8][32] = 9'b101101110;
assign F[8][33] = 9'b101101010;
assign F[8][34] = 9'b100100001;
assign F[8][35] = 9'b110001101;
assign F[8][36] = 9'b111111111;
assign F[8][37] = 9'b111111111;
assign F[8][38] = 9'b111111111;
assign F[9][25] = 9'b111111111;
assign F[9][26] = 9'b111111111;
assign F[9][27] = 9'b101110001;
assign F[9][28] = 9'b110011100;
assign F[9][29] = 9'b101001001;
assign F[9][30] = 9'b100100001;
assign F[9][31] = 9'b100100001;
assign F[9][32] = 9'b100100001;
assign F[9][33] = 9'b100100001;
assign F[9][34] = 9'b101101101;
assign F[9][35] = 9'b110011100;
assign F[9][36] = 9'b101110001;
assign F[9][37] = 9'b111111111;
assign F[9][38] = 9'b111111111;
assign F[10][24] = 9'b111111111;
assign F[10][25] = 9'b111111111;
assign F[10][26] = 9'b101110110;
assign F[10][27] = 9'b100101110;
assign F[10][28] = 9'b101110101;
assign F[10][29] = 9'b101101101;
assign F[10][30] = 9'b101000110;
assign F[10][31] = 9'b101000101;
assign F[10][32] = 9'b101000101;
assign F[10][33] = 9'b101000101;
assign F[10][34] = 9'b101101101;
assign F[10][35] = 9'b101010001;
assign F[10][36] = 9'b100101110;
assign F[10][37] = 9'b110011111;
assign F[10][38] = 9'b111111111;
assign F[10][39] = 9'b111111111;
assign F[11][24] = 9'b111111111;
assign F[11][25] = 9'b111111111;
assign F[11][26] = 9'b101110001;
assign F[11][27] = 9'b101110001;
assign F[11][28] = 9'b110011100;
assign F[11][29] = 9'b110010000;
assign F[11][30] = 9'b101101101;
assign F[11][31] = 9'b101101101;
assign F[11][32] = 9'b101101101;
assign F[11][33] = 9'b101101101;
assign F[11][34] = 9'b110010000;
assign F[11][35] = 9'b110010101;
assign F[11][36] = 9'b101010001;
assign F[11][37] = 9'b101110101;
assign F[11][38] = 9'b111111111;
assign F[11][39] = 9'b111111111;
assign F[12][24] = 9'b111111111;
assign F[12][25] = 9'b110010010;
assign F[12][26] = 9'b100000000;
assign F[12][27] = 9'b100000001;
assign F[12][28] = 9'b100100000;
assign F[12][29] = 9'b100100100;
assign F[12][30] = 9'b101001001;
assign F[12][31] = 9'b101110010;
assign F[12][32] = 9'b110011110;
assign F[12][33] = 9'b101101101;
assign F[12][34] = 9'b100100100;
assign F[12][35] = 9'b100100000;
assign F[12][36] = 9'b100000001;
assign F[12][37] = 9'b100000000;
assign F[12][38] = 9'b111111111;
assign F[12][39] = 9'b111111111;
assign F[13][24] = 9'b111111111;
assign F[13][25] = 9'b110001110;
assign F[13][26] = 9'b100000000;
assign F[13][27] = 9'b100000000;
assign F[13][28] = 9'b100000000;
assign F[13][29] = 9'b100000000;
assign F[13][30] = 9'b100100101;
assign F[13][31] = 9'b101110011;
assign F[13][32] = 9'b101110111;
assign F[13][33] = 9'b101001010;
assign F[13][34] = 9'b100000001;
assign F[13][35] = 9'b100000000;
assign F[13][36] = 9'b100000000;
assign F[13][37] = 9'b100000000;
assign F[13][38] = 9'b111111111;
assign F[13][39] = 9'b111111111;
assign F[14][24] = 9'b111111111;
assign F[14][25] = 9'b110010010;
assign F[14][26] = 9'b100000000;
assign F[14][27] = 9'b100100000;
assign F[14][28] = 9'b100100000;
assign F[14][29] = 9'b100000000;
assign F[14][30] = 9'b100100101;
assign F[14][31] = 9'b101110011;
assign F[14][32] = 9'b101110111;
assign F[14][33] = 9'b101001001;
assign F[14][34] = 9'b100000001;
assign F[14][35] = 9'b100000000;
assign F[14][36] = 9'b100000000;
assign F[14][37] = 9'b100000000;
assign F[14][38] = 9'b111111111;
assign F[14][39] = 9'b111111111;
assign F[15][24] = 9'b111111111;
assign F[15][25] = 9'b110010010;
assign F[15][26] = 9'b100000000;
assign F[15][27] = 9'b100100000;
assign F[15][28] = 9'b100100000;
assign F[15][29] = 9'b100000000;
assign F[15][30] = 9'b100100101;
assign F[15][31] = 9'b101110011;
assign F[15][32] = 9'b101110111;
assign F[15][33] = 9'b101001001;
assign F[15][34] = 9'b100000001;
assign F[15][35] = 9'b100000000;
assign F[15][36] = 9'b100000000;
assign F[15][37] = 9'b100000000;
assign F[15][38] = 9'b111111111;
assign F[15][39] = 9'b111111111;
assign F[16][24] = 9'b111111111;
assign F[16][25] = 9'b110010010;
assign F[16][26] = 9'b100000000;
assign F[16][27] = 9'b100100000;
assign F[16][28] = 9'b100000000;
assign F[16][29] = 9'b100000000;
assign F[16][30] = 9'b100100101;
assign F[16][31] = 9'b101110011;
assign F[16][32] = 9'b101110111;
assign F[16][33] = 9'b101001001;
assign F[16][34] = 9'b100000001;
assign F[16][35] = 9'b100000000;
assign F[16][36] = 9'b100000000;
assign F[16][37] = 9'b100000000;
assign F[16][38] = 9'b111111111;
assign F[16][39] = 9'b111111111;
assign F[17][24] = 9'b111111111;
assign F[17][25] = 9'b111111111;
assign F[17][26] = 9'b101001001;
assign F[17][27] = 9'b100000000;
assign F[17][28] = 9'b100100000;
assign F[17][29] = 9'b100000000;
assign F[17][30] = 9'b100100101;
assign F[17][31] = 9'b101110011;
assign F[17][32] = 9'b110011111;
assign F[17][33] = 9'b101001001;
assign F[17][34] = 9'b100000000;
assign F[17][35] = 9'b100000000;
assign F[17][36] = 9'b100000000;
assign F[17][37] = 9'b101000101;
assign F[17][38] = 9'b111111111;
assign F[17][39] = 9'b111111111;
assign F[18][24] = 9'b111111111;
assign F[18][25] = 9'b111111111;
assign F[18][26] = 9'b110111111;
assign F[18][27] = 9'b100001001;
assign F[18][28] = 9'b101110001;
assign F[18][29] = 9'b110110100;
assign F[18][30] = 9'b110010100;
assign F[18][31] = 9'b101101100;
assign F[18][32] = 9'b101110000;
assign F[18][33] = 9'b110111100;
assign F[18][34] = 9'b110110100;
assign F[18][35] = 9'b110010000;
assign F[18][36] = 9'b100101101;
assign F[18][37] = 9'b101110010;
assign F[18][38] = 9'b111111111;
assign F[18][39] = 9'b111111111;
assign F[19][23] = 9'b111111111;
assign F[19][24] = 9'b111111111;
assign F[19][25] = 9'b111111111;
assign F[19][26] = 9'b110011111;
assign F[19][27] = 9'b100101110;
assign F[19][28] = 9'b101110101;
assign F[19][29] = 9'b110011101;
assign F[19][30] = 9'b110011101;
assign F[19][31] = 9'b101010001;
assign F[19][32] = 9'b101110001;
assign F[19][33] = 9'b110011101;
assign F[19][34] = 9'b110011101;
assign F[19][35] = 9'b101110101;
assign F[19][36] = 9'b100101110;
assign F[19][37] = 9'b101110011;
assign F[19][38] = 9'b111111111;
assign F[19][39] = 9'b111111111;
assign F[19][40] = 9'b111111111;
assign F[20][22] = 9'b111111111;
assign F[20][23] = 9'b111111111;
assign F[20][24] = 9'b111111111;
assign F[20][25] = 9'b100101000;
assign F[20][26] = 9'b100001001;
assign F[20][27] = 9'b101010001;
assign F[20][28] = 9'b100101101;
assign F[20][29] = 9'b100001001;
assign F[20][30] = 9'b100001001;
assign F[20][31] = 9'b100001001;
assign F[20][32] = 9'b100001001;
assign F[20][33] = 9'b100001001;
assign F[20][34] = 9'b100001001;
assign F[20][35] = 9'b101010001;
assign F[20][36] = 9'b100001001;
assign F[20][37] = 9'b100000100;
assign F[20][38] = 9'b101001101;
assign F[20][39] = 9'b111111111;
assign F[20][40] = 9'b111111111;
assign F[20][41] = 9'b111111111;
assign F[21][21] = 9'b111111111;
assign F[21][22] = 9'b111111111;
assign F[21][23] = 9'b110111111;
assign F[21][24] = 9'b100001001;
assign F[21][25] = 9'b100000100;
assign F[21][26] = 9'b101001100;
assign F[21][27] = 9'b100101100;
assign F[21][28] = 9'b100001000;
assign F[21][29] = 9'b100001000;
assign F[21][30] = 9'b100001000;
assign F[21][31] = 9'b100001000;
assign F[21][32] = 9'b100001000;
assign F[21][33] = 9'b100001000;
assign F[21][34] = 9'b100001000;
assign F[21][35] = 9'b100001000;
assign F[21][36] = 9'b101001100;
assign F[21][37] = 9'b100000100;
assign F[21][38] = 9'b100001000;
assign F[21][39] = 9'b100101101;
assign F[21][40] = 9'b111111111;
assign F[21][41] = 9'b111111111;
assign F[22][21] = 9'b111111111;
assign F[22][22] = 9'b111111111;
assign F[22][23] = 9'b100101101;
assign F[22][24] = 9'b100000100;
assign F[22][25] = 9'b100101000;
assign F[22][26] = 9'b100101100;
assign F[22][27] = 9'b101001101;
assign F[22][28] = 9'b101110001;
assign F[22][29] = 9'b101110001;
assign F[22][30] = 9'b100001000;
assign F[22][31] = 9'b100001000;
assign F[22][32] = 9'b100001000;
assign F[22][33] = 9'b100101101;
assign F[22][34] = 9'b101001101;
assign F[22][35] = 9'b100101101;
assign F[22][36] = 9'b100101100;
assign F[22][37] = 9'b101001100;
assign F[22][38] = 9'b100001000;
assign F[22][39] = 9'b100001000;
assign F[22][40] = 9'b101110001;
assign F[22][41] = 9'b111111111;
assign F[22][42] = 9'b111111111;
assign F[23][20] = 9'b111111111;
assign F[23][21] = 9'b111111111;
assign F[23][22] = 9'b110010110;
assign F[23][23] = 9'b100001000;
assign F[23][24] = 9'b100001000;
assign F[23][25] = 9'b100000100;
assign F[23][26] = 9'b100001000;
assign F[23][27] = 9'b110010110;
assign F[23][28] = 9'b111111111;
assign F[23][29] = 9'b110011110;
assign F[23][30] = 9'b100001000;
assign F[23][31] = 9'b100001000;
assign F[23][32] = 9'b100001000;
assign F[23][33] = 9'b101110001;
assign F[23][34] = 9'b110010110;
assign F[23][35] = 9'b110010110;
assign F[23][36] = 9'b100001001;
assign F[23][37] = 9'b100000100;
assign F[23][38] = 9'b100000100;
assign F[23][39] = 9'b100001000;
assign F[23][40] = 9'b100001000;
assign F[23][41] = 9'b111111111;
assign F[23][42] = 9'b111111111;
assign F[24][20] = 9'b111111111;
assign F[24][21] = 9'b111111111;
assign F[24][22] = 9'b100101001;
assign F[24][23] = 9'b100101001;
assign F[24][24] = 9'b100001000;
assign F[24][25] = 9'b100000100;
assign F[24][26] = 9'b100001000;
assign F[24][27] = 9'b101001101;
assign F[24][28] = 9'b101110001;
assign F[24][29] = 9'b101001101;
assign F[24][30] = 9'b100001000;
assign F[24][31] = 9'b100001000;
assign F[24][32] = 9'b100001000;
assign F[24][33] = 9'b101110001;
assign F[24][34] = 9'b110111111;
assign F[24][35] = 9'b110111111;
assign F[24][36] = 9'b100101101;
assign F[24][37] = 9'b100000100;
assign F[24][38] = 9'b100000100;
assign F[24][39] = 9'b100101101;
assign F[24][40] = 9'b100001000;
assign F[24][41] = 9'b101001101;
assign F[24][42] = 9'b111111111;
assign F[24][43] = 9'b111111111;
assign F[25][20] = 9'b111111111;
assign F[25][21] = 9'b110111111;
assign F[25][22] = 9'b100001000;
assign F[25][23] = 9'b101110001;
assign F[25][24] = 9'b100000100;
assign F[25][25] = 9'b100000100;
assign F[25][26] = 9'b100001000;
assign F[25][27] = 9'b101001101;
assign F[25][28] = 9'b110010110;
assign F[25][29] = 9'b101010001;
assign F[25][30] = 9'b100001000;
assign F[25][31] = 9'b100001000;
assign F[25][32] = 9'b100001000;
assign F[25][33] = 9'b100101001;
assign F[25][34] = 9'b100101101;
assign F[25][35] = 9'b100101001;
assign F[25][36] = 9'b100001000;
assign F[25][37] = 9'b100001000;
assign F[25][38] = 9'b100000100;
assign F[25][39] = 9'b101110001;
assign F[25][40] = 9'b100101101;
assign F[25][41] = 9'b100001000;
assign F[25][42] = 9'b111111111;
assign F[25][43] = 9'b111111111;
assign F[26][19] = 9'b111111111;
assign F[26][20] = 9'b111111111;
assign F[26][21] = 9'b101001101;
assign F[26][22] = 9'b101001101;
assign F[26][23] = 9'b101110001;
assign F[26][24] = 9'b100000000;
assign F[26][25] = 9'b100001000;
assign F[26][26] = 9'b100001000;
assign F[26][27] = 9'b100101101;
assign F[26][28] = 9'b100101101;
assign F[26][29] = 9'b100101101;
assign F[26][30] = 9'b100101101;
assign F[26][31] = 9'b100101001;
assign F[26][32] = 9'b100101001;
assign F[26][33] = 9'b100101101;
assign F[26][34] = 9'b100101101;
assign F[26][35] = 9'b100101101;
assign F[26][36] = 9'b100101001;
assign F[26][37] = 9'b100001000;
assign F[26][38] = 9'b100000100;
assign F[26][39] = 9'b101001101;
assign F[26][40] = 9'b101110001;
assign F[26][41] = 9'b100000100;
assign F[26][42] = 9'b101110010;
assign F[26][43] = 9'b111111111;
assign F[27][19] = 9'b111111111;
assign F[27][20] = 9'b111111111;
assign F[27][21] = 9'b100101101;
assign F[27][22] = 9'b101110001;
assign F[27][23] = 9'b100101101;
assign F[27][24] = 9'b100000100;
assign F[27][25] = 9'b100000100;
assign F[27][26] = 9'b100101101;
assign F[27][27] = 9'b101110001;
assign F[27][28] = 9'b101110001;
assign F[27][29] = 9'b101110001;
assign F[27][30] = 9'b101110001;
assign F[27][31] = 9'b101110001;
assign F[27][32] = 9'b101110001;
assign F[27][33] = 9'b101110001;
assign F[27][34] = 9'b101110001;
assign F[27][35] = 9'b101110001;
assign F[27][36] = 9'b101001101;
assign F[27][37] = 9'b100001000;
assign F[27][38] = 9'b100000100;
assign F[27][39] = 9'b100001000;
assign F[27][40] = 9'b101110001;
assign F[27][41] = 9'b100001000;
assign F[27][42] = 9'b101001101;
assign F[27][43] = 9'b111111111;
assign F[28][19] = 9'b111111111;
assign F[28][20] = 9'b111111111;
assign F[28][21] = 9'b100101101;
assign F[28][22] = 9'b100101001;
assign F[28][23] = 9'b100000100;
assign F[28][24] = 9'b100000100;
assign F[28][25] = 9'b100001000;
assign F[28][26] = 9'b100001000;
assign F[28][27] = 9'b100001000;
assign F[28][28] = 9'b100001000;
assign F[28][29] = 9'b100001000;
assign F[28][30] = 9'b100001000;
assign F[28][31] = 9'b100001000;
assign F[28][32] = 9'b100001000;
assign F[28][33] = 9'b100001000;
assign F[28][34] = 9'b100001000;
assign F[28][35] = 9'b100001000;
assign F[28][36] = 9'b100001000;
assign F[28][37] = 9'b100001001;
assign F[28][38] = 9'b100000100;
assign F[28][39] = 9'b100000100;
assign F[28][40] = 9'b101010001;
assign F[28][41] = 9'b100101101;
assign F[28][42] = 9'b101110001;
assign F[28][43] = 9'b111111111;
assign F[28][44] = 9'b111111111;
assign F[29][18] = 9'b111111111;
assign F[29][19] = 9'b111111111;
assign F[29][20] = 9'b111111111;
assign F[29][21] = 9'b110111111;
assign F[29][22] = 9'b110010110;
assign F[29][23] = 9'b110010001;
assign F[29][24] = 9'b100000100;
assign F[29][25] = 9'b100001000;
assign F[29][26] = 9'b100101101;
assign F[29][27] = 9'b101010001;
assign F[29][28] = 9'b101010001;
assign F[29][29] = 9'b101001101;
assign F[29][30] = 9'b101001101;
assign F[29][31] = 9'b101001101;
assign F[29][32] = 9'b101001101;
assign F[29][33] = 9'b101001101;
assign F[29][34] = 9'b101001101;
assign F[29][35] = 9'b101010001;
assign F[29][36] = 9'b100101101;
assign F[29][37] = 9'b100001000;
assign F[29][38] = 9'b100000100;
assign F[29][39] = 9'b101101101;
assign F[29][40] = 9'b111111111;
assign F[29][41] = 9'b111111111;
assign F[29][42] = 9'b111111111;
assign F[29][43] = 9'b111111111;
assign F[29][44] = 9'b111111111;
assign F[30][18] = 9'b111111111;
assign F[30][19] = 9'b111111111;
assign F[30][20] = 9'b111111111;
assign F[30][21] = 9'b111111111;
assign F[30][22] = 9'b111111111;
assign F[30][23] = 9'b111111111;
assign F[30][24] = 9'b110111111;
assign F[30][25] = 9'b100001000;
assign F[30][26] = 9'b100101101;
assign F[30][27] = 9'b101110001;
assign F[30][28] = 9'b101110001;
assign F[30][29] = 9'b101110001;
assign F[30][30] = 9'b101110001;
assign F[30][31] = 9'b101110001;
assign F[30][32] = 9'b101110001;
assign F[30][33] = 9'b101110001;
assign F[30][34] = 9'b101110001;
assign F[30][35] = 9'b101110001;
assign F[30][36] = 9'b101001101;
assign F[30][37] = 9'b100001000;
assign F[30][38] = 9'b100101101;
assign F[30][39] = 9'b111111111;
assign F[30][40] = 9'b111111111;
assign F[30][41] = 9'b111111111;
assign F[30][42] = 9'b111111111;
assign F[30][43] = 9'b111111111;
assign F[30][44] = 9'b111111111;
assign F[31][18] = 9'b111111111;
assign F[31][19] = 9'b111111111;
assign F[31][20] = 9'b111111111;
assign F[31][21] = 9'b111111111;
assign F[31][22] = 9'b111111111;
assign F[31][23] = 9'b111111111;
assign F[31][24] = 9'b111111111;
assign F[31][25] = 9'b100101001;
assign F[31][26] = 9'b100001000;
assign F[31][27] = 9'b100001000;
assign F[31][28] = 9'b100001000;
assign F[31][29] = 9'b100001000;
assign F[31][30] = 9'b100001000;
assign F[31][31] = 9'b100001000;
assign F[31][32] = 9'b100001000;
assign F[31][33] = 9'b100001000;
assign F[31][34] = 9'b100001000;
assign F[31][35] = 9'b100001000;
assign F[31][36] = 9'b100001000;
assign F[31][37] = 9'b100001000;
assign F[31][38] = 9'b101001101;
assign F[31][39] = 9'b111111111;
assign F[31][40] = 9'b111111111;
assign F[31][41] = 9'b111111111;
assign F[31][42] = 9'b111111111;
assign F[31][43] = 9'b111111111;
assign F[31][44] = 9'b111111111;
assign F[32][18] = 9'b111111111;
assign F[32][19] = 9'b111111111;
assign F[32][20] = 9'b111111111;
assign F[32][21] = 9'b111111111;
assign F[32][22] = 9'b111111111;
assign F[32][23] = 9'b111111111;
assign F[32][24] = 9'b111111111;
assign F[32][25] = 9'b100001001;
assign F[32][26] = 9'b100001000;
assign F[32][27] = 9'b100001000;
assign F[32][28] = 9'b100001000;
assign F[32][29] = 9'b100001001;
assign F[32][30] = 9'b100001001;
assign F[32][31] = 9'b100001000;
assign F[32][32] = 9'b100001000;
assign F[32][33] = 9'b100001000;
assign F[32][34] = 9'b100001000;
assign F[32][35] = 9'b100001000;
assign F[32][36] = 9'b100001000;
assign F[32][37] = 9'b100001000;
assign F[32][38] = 9'b100101101;
assign F[32][39] = 9'b111111111;
assign F[32][40] = 9'b111111111;
assign F[32][41] = 9'b111111111;
assign F[32][42] = 9'b111111111;
assign F[32][43] = 9'b111111111;
assign F[32][44] = 9'b111111111;
assign F[33][18] = 9'b111111111;
assign F[33][19] = 9'b111111111;
assign F[33][20] = 9'b111111111;
assign F[33][21] = 9'b111111111;
assign F[33][22] = 9'b111111111;
assign F[33][23] = 9'b111111111;
assign F[33][24] = 9'b101101101;
assign F[33][25] = 9'b100000100;
assign F[33][26] = 9'b100000100;
assign F[33][27] = 9'b100000100;
assign F[33][28] = 9'b100000100;
assign F[33][29] = 9'b100000100;
assign F[33][30] = 9'b100000100;
assign F[33][31] = 9'b100000100;
assign F[33][32] = 9'b100000100;
assign F[33][33] = 9'b100000100;
assign F[33][34] = 9'b100000100;
assign F[33][35] = 9'b100000100;
assign F[33][36] = 9'b100000100;
assign F[33][37] = 9'b100000100;
assign F[33][38] = 9'b100000100;
assign F[33][39] = 9'b110010110;
assign F[33][40] = 9'b111111111;
assign F[33][41] = 9'b111111111;
assign F[33][42] = 9'b111111111;
assign F[33][43] = 9'b111111111;
assign F[33][44] = 9'b111111111;
assign F[34][18] = 9'b111111111;
assign F[34][19] = 9'b111111111;
assign F[34][20] = 9'b111111111;
assign F[34][21] = 9'b111111111;
assign F[34][22] = 9'b111111111;
assign F[34][23] = 9'b111111111;
assign F[34][24] = 9'b101110001;
assign F[34][25] = 9'b100000100;
assign F[34][26] = 9'b100000100;
assign F[34][27] = 9'b100001000;
assign F[34][28] = 9'b100101000;
assign F[34][29] = 9'b111101000;
assign F[34][30] = 9'b111101000;
assign F[34][31] = 9'b100001000;
assign F[34][32] = 9'b100101001;
assign F[34][33] = 9'b101001101;
assign F[34][34] = 9'b101001101;
assign F[34][35] = 9'b101001101;
assign F[34][36] = 9'b100101101;
assign F[34][37] = 9'b100101101;
assign F[34][38] = 9'b100001000;
assign F[34][39] = 9'b110010110;
assign F[34][40] = 9'b111111111;
assign F[34][41] = 9'b111111111;
assign F[34][42] = 9'b111111111;
assign F[34][43] = 9'b111111111;
assign F[34][44] = 9'b111111111;
assign F[35][19] = 9'b111111111;
assign F[35][20] = 9'b111111111;
assign F[35][22] = 9'b111111111;
assign F[35][23] = 9'b111111111;
assign F[35][24] = 9'b101101101;
assign F[35][25] = 9'b100000000;
assign F[35][26] = 9'b100000100;
assign F[35][27] = 9'b100000100;
assign F[35][28] = 9'b100000100;
assign F[35][29] = 9'b101100100;
assign F[35][30] = 9'b101000100;
assign F[35][31] = 9'b100000100;
assign F[35][32] = 9'b100000100;
assign F[35][33] = 9'b100000100;
assign F[35][34] = 9'b100000100;
assign F[35][35] = 9'b100000100;
assign F[35][36] = 9'b100000100;
assign F[35][37] = 9'b100000100;
assign F[35][38] = 9'b100000100;
assign F[35][39] = 9'b110010110;
assign F[35][40] = 9'b111111111;
assign F[35][42] = 9'b111111111;
assign F[35][43] = 9'b111111111;
assign F[36][23] = 9'b111111111;
assign F[36][24] = 9'b101110001;
assign F[36][25] = 9'b100000100;
assign F[36][26] = 9'b100001000;
assign F[36][27] = 9'b100001000;
assign F[36][28] = 9'b100001000;
assign F[36][29] = 9'b100001000;
assign F[36][30] = 9'b100001000;
assign F[36][31] = 9'b100000100;
assign F[36][32] = 9'b100001000;
assign F[36][33] = 9'b100001000;
assign F[36][34] = 9'b100001000;
assign F[36][35] = 9'b100001000;
assign F[36][36] = 9'b100101001;
assign F[36][37] = 9'b100101001;
assign F[36][38] = 9'b100000100;
assign F[36][39] = 9'b110111110;
assign F[36][40] = 9'b111111111;
assign F[37][23] = 9'b111111111;
assign F[37][24] = 9'b101110001;
assign F[37][25] = 9'b100001000;
assign F[37][26] = 9'b100001000;
assign F[37][27] = 9'b100001000;
assign F[37][28] = 9'b100001000;
assign F[37][29] = 9'b100001000;
assign F[37][30] = 9'b100001000;
assign F[37][31] = 9'b100001000;
assign F[37][32] = 9'b100001000;
assign F[37][33] = 9'b100001000;
assign F[37][34] = 9'b100001000;
assign F[37][35] = 9'b100001000;
assign F[37][36] = 9'b101001101;
assign F[37][37] = 9'b101110001;
assign F[37][38] = 9'b100001000;
assign F[37][39] = 9'b110111111;
assign F[37][40] = 9'b111111111;
assign F[38][23] = 9'b111111111;
assign F[38][24] = 9'b101110001;
assign F[38][25] = 9'b100001000;
assign F[38][26] = 9'b100001000;
assign F[38][27] = 9'b100001000;
assign F[38][28] = 9'b100001000;
assign F[38][29] = 9'b100001000;
assign F[38][30] = 9'b100001000;
assign F[38][31] = 9'b100001000;
assign F[38][32] = 9'b100001000;
assign F[38][33] = 9'b100001000;
assign F[38][34] = 9'b100001000;
assign F[38][35] = 9'b100001000;
assign F[38][36] = 9'b101001101;
assign F[38][37] = 9'b101010001;
assign F[38][38] = 9'b100001000;
assign F[38][39] = 9'b110111111;
assign F[38][40] = 9'b111111111;
assign F[39][23] = 9'b111111111;
assign F[39][24] = 9'b101110001;
assign F[39][25] = 9'b100001000;
assign F[39][26] = 9'b100001000;
assign F[39][27] = 9'b100001000;
assign F[39][28] = 9'b100001000;
assign F[39][29] = 9'b100001000;
assign F[39][30] = 9'b100001000;
assign F[39][31] = 9'b101110001;
assign F[39][32] = 9'b101001101;
assign F[39][33] = 9'b100001000;
assign F[39][34] = 9'b100001000;
assign F[39][35] = 9'b100001000;
assign F[39][36] = 9'b101001101;
assign F[39][37] = 9'b101110001;
assign F[39][38] = 9'b100001000;
assign F[39][39] = 9'b110111111;
assign F[39][40] = 9'b111111111;
assign F[40][23] = 9'b111111111;
assign F[40][24] = 9'b101110001;
assign F[40][25] = 9'b100001000;
assign F[40][26] = 9'b100001000;
assign F[40][27] = 9'b100001000;
assign F[40][28] = 9'b100001000;
assign F[40][29] = 9'b100001000;
assign F[40][30] = 9'b100001000;
assign F[40][31] = 9'b101110001;
assign F[40][32] = 9'b101001101;
assign F[40][33] = 9'b100001000;
assign F[40][34] = 9'b100001000;
assign F[40][35] = 9'b100001000;
assign F[40][36] = 9'b100001001;
assign F[40][37] = 9'b101001101;
assign F[40][38] = 9'b100001000;
assign F[40][39] = 9'b110111111;
assign F[40][40] = 9'b111111111;
assign F[41][23] = 9'b111111111;
assign F[41][24] = 9'b101110001;
assign F[41][25] = 9'b100001000;
assign F[41][26] = 9'b100001000;
assign F[41][27] = 9'b100001000;
assign F[41][28] = 9'b100001000;
assign F[41][29] = 9'b100001000;
assign F[41][30] = 9'b100001000;
assign F[41][31] = 9'b101110001;
assign F[41][32] = 9'b101001101;
assign F[41][33] = 9'b100001000;
assign F[41][34] = 9'b100001000;
assign F[41][35] = 9'b100001000;
assign F[41][36] = 9'b100101101;
assign F[41][37] = 9'b100101001;
assign F[41][38] = 9'b100001000;
assign F[41][39] = 9'b110111111;
assign F[41][40] = 9'b111111111;
assign F[42][23] = 9'b111111111;
assign F[42][24] = 9'b101110001;
assign F[42][25] = 9'b100001000;
assign F[42][26] = 9'b100001000;
assign F[42][27] = 9'b100001000;
assign F[42][28] = 9'b100001000;
assign F[42][29] = 9'b100001000;
assign F[42][30] = 9'b100001000;
assign F[42][31] = 9'b101110001;
assign F[42][32] = 9'b101001101;
assign F[42][33] = 9'b100001000;
assign F[42][34] = 9'b100001000;
assign F[42][35] = 9'b100001000;
assign F[42][36] = 9'b101001101;
assign F[42][37] = 9'b101110001;
assign F[42][38] = 9'b100001000;
assign F[42][39] = 9'b110111111;
assign F[42][40] = 9'b111111111;
assign F[43][23] = 9'b111111111;
assign F[43][24] = 9'b101110001;
assign F[43][25] = 9'b100001000;
assign F[43][26] = 9'b100001000;
assign F[43][27] = 9'b100001000;
assign F[43][28] = 9'b100001000;
assign F[43][29] = 9'b100001000;
assign F[43][30] = 9'b100001000;
assign F[43][31] = 9'b101110001;
assign F[43][32] = 9'b101001101;
assign F[43][33] = 9'b100001000;
assign F[43][34] = 9'b100001000;
assign F[43][35] = 9'b100001000;
assign F[43][36] = 9'b101001101;
assign F[43][37] = 9'b101010001;
assign F[43][38] = 9'b100001000;
assign F[43][39] = 9'b110111111;
assign F[43][40] = 9'b111111111;
assign F[44][23] = 9'b111111111;
assign F[44][24] = 9'b101110001;
assign F[44][25] = 9'b100001000;
assign F[44][26] = 9'b100001000;
assign F[44][27] = 9'b100001000;
assign F[44][28] = 9'b100001000;
assign F[44][29] = 9'b100001000;
assign F[44][30] = 9'b100001000;
assign F[44][31] = 9'b101110001;
assign F[44][32] = 9'b101001101;
assign F[44][33] = 9'b100001000;
assign F[44][34] = 9'b100001000;
assign F[44][35] = 9'b100001000;
assign F[44][36] = 9'b101001101;
assign F[44][37] = 9'b101010001;
assign F[44][38] = 9'b100001000;
assign F[44][39] = 9'b110111111;
assign F[44][40] = 9'b111111111;
assign F[45][23] = 9'b111111111;
assign F[45][24] = 9'b101110001;
assign F[45][25] = 9'b100001000;
assign F[45][26] = 9'b100001000;
assign F[45][27] = 9'b100001000;
assign F[45][28] = 9'b100001000;
assign F[45][29] = 9'b100001000;
assign F[45][30] = 9'b100001000;
assign F[45][31] = 9'b101110001;
assign F[45][32] = 9'b101001101;
assign F[45][33] = 9'b100001000;
assign F[45][34] = 9'b100001000;
assign F[45][35] = 9'b100001000;
assign F[45][36] = 9'b100101001;
assign F[45][37] = 9'b100001001;
assign F[45][38] = 9'b100001000;
assign F[45][39] = 9'b110111111;
assign F[45][40] = 9'b111111111;
assign F[46][23] = 9'b111111111;
assign F[46][24] = 9'b101101101;
assign F[46][25] = 9'b100000000;
assign F[46][26] = 9'b100000000;
assign F[46][27] = 9'b100000000;
assign F[46][28] = 9'b100000000;
assign F[46][29] = 9'b100000000;
assign F[46][30] = 9'b100000000;
assign F[46][31] = 9'b101001101;
assign F[46][32] = 9'b100101000;
assign F[46][33] = 9'b100000000;
assign F[46][34] = 9'b100000000;
assign F[46][35] = 9'b100000000;
assign F[46][36] = 9'b100000000;
assign F[46][37] = 9'b100000000;
assign F[46][38] = 9'b100000000;
assign F[46][39] = 9'b110010010;
assign F[46][40] = 9'b111111111;
assign F[47][23] = 9'b111111111;
assign F[47][24] = 9'b110010001;
assign F[47][25] = 9'b100000000;
assign F[47][26] = 9'b100000000;
assign F[47][27] = 9'b100000000;
assign F[47][28] = 9'b100000000;
assign F[47][29] = 9'b100000000;
assign F[47][30] = 9'b100000000;
assign F[47][31] = 9'b110010001;
assign F[47][32] = 9'b101101101;
assign F[47][33] = 9'b100000000;
assign F[47][34] = 9'b100000000;
assign F[47][35] = 9'b100000000;
assign F[47][36] = 9'b100000000;
assign F[47][37] = 9'b100000000;
assign F[47][38] = 9'b100000000;
assign F[47][39] = 9'b111111111;
assign F[47][40] = 9'b111111111;
assign F[48][23] = 9'b111111111;
assign F[48][24] = 9'b111111111;
assign F[48][25] = 9'b100000000;
assign F[48][26] = 9'b100000000;
assign F[48][27] = 9'b100000000;
assign F[48][28] = 9'b100000000;
assign F[48][29] = 9'b100000000;
assign F[48][30] = 9'b100000000;
assign F[48][31] = 9'b111111111;
assign F[48][32] = 9'b110010001;
assign F[48][33] = 9'b100000000;
assign F[48][34] = 9'b100000000;
assign F[48][35] = 9'b100000000;
assign F[48][36] = 9'b100000000;
assign F[48][37] = 9'b100000000;
assign F[48][38] = 9'b100100100;
assign F[48][39] = 9'b111111111;
assign F[48][40] = 9'b111111111;
assign F[49][23] = 9'b111111111;
assign F[49][24] = 9'b101001001;
assign F[49][25] = 9'b100000000;
assign F[49][26] = 9'b100000000;
assign F[49][27] = 9'b100000000;
assign F[49][28] = 9'b100000000;
assign F[49][29] = 9'b100000000;
assign F[49][30] = 9'b100000000;
assign F[49][31] = 9'b101001001;
assign F[49][32] = 9'b100100100;
assign F[49][33] = 9'b100000000;
assign F[49][34] = 9'b100000000;
assign F[49][35] = 9'b100000000;
assign F[49][36] = 9'b100000000;
assign F[49][37] = 9'b100000000;
assign F[49][38] = 9'b100000000;
assign F[49][39] = 9'b110010001;
assign F[49][40] = 9'b111111111;
assign F[50][23] = 9'b111111111;
assign F[50][24] = 9'b101101101;
assign F[50][25] = 9'b100100100;
assign F[50][26] = 9'b100100100;
assign F[50][27] = 9'b100100100;
assign F[50][28] = 9'b100100100;
assign F[50][29] = 9'b100100100;
assign F[50][30] = 9'b100100100;
assign F[50][31] = 9'b101101101;
assign F[50][32] = 9'b101001001;
assign F[50][33] = 9'b100100100;
assign F[50][34] = 9'b100100100;
assign F[50][35] = 9'b100100100;
assign F[50][36] = 9'b100100100;
assign F[50][37] = 9'b100100100;
assign F[50][38] = 9'b100100100;
assign F[50][39] = 9'b110110110;
assign F[50][40] = 9'b111111111;
assign F[51][23] = 9'b111111111;
assign F[51][24] = 9'b111111111;
assign F[51][25] = 9'b111111111;
assign F[51][26] = 9'b111111111;
assign F[51][27] = 9'b111111111;
assign F[51][28] = 9'b111111111;
assign F[51][29] = 9'b111111111;
assign F[51][30] = 9'b111111111;
assign F[51][31] = 9'b111111111;
assign F[51][32] = 9'b111111111;
assign F[51][33] = 9'b111111111;
assign F[51][34] = 9'b111111111;
assign F[51][35] = 9'b111111111;
assign F[51][36] = 9'b111111111;
assign F[51][37] = 9'b111111111;
assign F[51][38] = 9'b111111111;
assign F[51][39] = 9'b111111111;
assign F[51][40] = 9'b111111111;
assign F[52][23] = 9'b111111111;
assign F[52][24] = 9'b111111111;
assign F[52][25] = 9'b111111111;
assign F[52][26] = 9'b111111111;
assign F[52][27] = 9'b111111111;
assign F[52][28] = 9'b111111111;
assign F[52][29] = 9'b111111111;
assign F[52][30] = 9'b111111111;
assign F[52][31] = 9'b111111111;
assign F[52][32] = 9'b111111111;
assign F[52][33] = 9'b111111111;
assign F[52][34] = 9'b111111111;
assign F[52][35] = 9'b111111111;
assign F[52][36] = 9'b111111111;
assign F[52][37] = 9'b111111111;
assign F[52][38] = 9'b111111111;
assign F[52][39] = 9'b111111111;
assign F[52][40] = 9'b111111111;
assign F[53][23] = 9'b111111111;
assign F[53][24] = 9'b111110010;
assign F[53][25] = 9'b111101001;
assign F[53][26] = 9'b111101001;
assign F[53][27] = 9'b111101001;
assign F[53][28] = 9'b111111111;
assign F[53][29] = 9'b111111111;
assign F[53][30] = 9'b101101101;
assign F[53][31] = 9'b101101101;
assign F[53][32] = 9'b111111111;
assign F[53][33] = 9'b110010001;
assign F[53][34] = 9'b110010001;
assign F[53][35] = 9'b111111111;
assign F[53][36] = 9'b111111111;
assign F[53][37] = 9'b101101101;
assign F[53][38] = 9'b101101101;
assign F[53][39] = 9'b101101101;
assign F[53][40] = 9'b111111111;
assign F[53][41] = 9'b111111111;
assign F[54][23] = 9'b111111111;
assign F[54][24] = 9'b111110101;
assign F[54][25] = 9'b111101100;
assign F[54][26] = 9'b111101100;
assign F[54][27] = 9'b111101100;
assign F[54][28] = 9'b111111110;
assign F[54][29] = 9'b101001101;
assign F[54][30] = 9'b101101101;
assign F[54][31] = 9'b101101101;
assign F[54][32] = 9'b101101101;
assign F[54][33] = 9'b101101101;
assign F[54][34] = 9'b101101101;
assign F[54][35] = 9'b111111111;
assign F[54][36] = 9'b110010001;
assign F[54][37] = 9'b100100100;
assign F[54][38] = 9'b111111111;
assign F[54][39] = 9'b100100100;
assign F[54][40] = 9'b111111111;
assign F[54][41] = 9'b111111111;
assign F[55][23] = 9'b111111111;
assign F[55][24] = 9'b111110001;
assign F[55][25] = 9'b111101000;
assign F[55][26] = 9'b111101000;
assign F[55][27] = 9'b111101000;
assign F[55][28] = 9'b111111110;
assign F[55][29] = 9'b100101000;
assign F[55][30] = 9'b101001001;
assign F[55][31] = 9'b101001001;
assign F[55][32] = 9'b101001001;
assign F[55][33] = 9'b101101101;
assign F[55][34] = 9'b101001001;
assign F[55][35] = 9'b111111111;
assign F[55][36] = 9'b110010001;
assign F[55][37] = 9'b100100100;
assign F[55][38] = 9'b111111111;
assign F[55][39] = 9'b100100100;
assign F[55][40] = 9'b111111111;
assign F[55][41] = 9'b111111111;
assign F[56][23] = 9'b111111111;
assign F[56][24] = 9'b111110110;
assign F[56][25] = 9'b111101101;
assign F[56][26] = 9'b111101101;
assign F[56][27] = 9'b111101101;
assign F[56][28] = 9'b111111111;
assign F[56][29] = 9'b110010010;
assign F[56][30] = 9'b111111111;
assign F[56][31] = 9'b111111111;
assign F[56][32] = 9'b110110110;
assign F[56][33] = 9'b111111111;
assign F[56][34] = 9'b101101101;
assign F[56][35] = 9'b110010001;
assign F[56][36] = 9'b111111111;
assign F[56][37] = 9'b110010010;
assign F[56][38] = 9'b110010001;
assign F[56][39] = 9'b110110110;
assign F[56][40] = 9'b111111111;
assign F[56][41] = 9'b111111111;
assign F[57][23] = 9'b111111111;
assign F[57][24] = 9'b111111111;
assign F[57][25] = 9'b111111111;
assign F[57][26] = 9'b111111111;
assign F[57][27] = 9'b111111111;
assign F[57][28] = 9'b111111111;
assign F[57][29] = 9'b111111111;
assign F[57][30] = 9'b111111111;
assign F[57][31] = 9'b111111111;
assign F[57][32] = 9'b111111111;
assign F[57][33] = 9'b111111111;
assign F[57][34] = 9'b111111111;
assign F[57][35] = 9'b111111111;
assign F[57][36] = 9'b111111111;
assign F[57][37] = 9'b111111111;
assign F[57][38] = 9'b111111111;
assign F[57][39] = 9'b111111111;
assign F[57][40] = 9'b111111111;
//Total de Lineas = 1013
endmodule

