`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:25:57 02/07/2023 
// Design Name: 
// Module Name:    menuprincipal 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module menuprincipal(input [4:0]a,b, output [5:0]out);

sumador_de_5bits suma_0 (a,b,out);

endmodule
