`timescale 1ns / 1ps
module estado_alonso (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (F[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= F[vcount- posy][hcount- posx][7:5];
				green <= F[vcount- posy][hcount- posx][4:2];
            blue 	<= F[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 100;
parameter RESOLUCION_Y = 50;
wire [8:0] F[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign F[3][47] = 9'b100111101;
assign F[3][48] = 9'b100111101;
assign F[3][49] = 9'b100111101;
assign F[3][50] = 9'b100111101;
assign F[3][51] = 9'b100111101;
assign F[3][52] = 9'b100111101;
assign F[3][53] = 9'b100111101;
assign F[3][54] = 9'b100111101;
assign F[3][55] = 9'b100111101;
assign F[3][56] = 9'b100111101;
assign F[4][45] = 9'b100111101;
assign F[4][46] = 9'b100111101;
assign F[4][47] = 9'b100111101;
assign F[4][48] = 9'b100111101;
assign F[4][49] = 9'b100111101;
assign F[4][50] = 9'b100111101;
assign F[4][51] = 9'b100111101;
assign F[4][52] = 9'b100111101;
assign F[4][53] = 9'b100111101;
assign F[4][54] = 9'b100111101;
assign F[4][55] = 9'b100111101;
assign F[4][56] = 9'b100111101;
assign F[4][57] = 9'b100111101;
assign F[4][58] = 9'b100111101;
assign F[5][44] = 9'b100111101;
assign F[5][45] = 9'b100111101;
assign F[5][46] = 9'b100111101;
assign F[5][47] = 9'b100111101;
assign F[5][48] = 9'b100111101;
assign F[5][49] = 9'b100111101;
assign F[5][50] = 9'b100111101;
assign F[5][51] = 9'b100111101;
assign F[5][52] = 9'b100111101;
assign F[5][53] = 9'b100011101;
assign F[5][54] = 9'b100011101;
assign F[5][55] = 9'b100011101;
assign F[5][56] = 9'b100011101;
assign F[5][57] = 9'b100011101;
assign F[5][58] = 9'b100111101;
assign F[5][59] = 9'b100110101;
assign F[6][43] = 9'b100111101;
assign F[6][44] = 9'b100111101;
assign F[6][45] = 9'b100111101;
assign F[6][46] = 9'b100111101;
assign F[6][47] = 9'b100111101;
assign F[6][48] = 9'b100111101;
assign F[6][49] = 9'b100111101;
assign F[6][50] = 9'b100111101;
assign F[6][51] = 9'b100111101;
assign F[6][52] = 9'b101011101;
assign F[6][53] = 9'b101111110;
assign F[6][54] = 9'b101111110;
assign F[6][55] = 9'b101111110;
assign F[6][56] = 9'b101111110;
assign F[6][57] = 9'b101111110;
assign F[6][58] = 9'b100111101;
assign F[6][59] = 9'b100111101;
assign F[6][60] = 9'b100111101;
assign F[7][43] = 9'b100111101;
assign F[7][44] = 9'b100111101;
assign F[7][45] = 9'b100111101;
assign F[7][46] = 9'b100111101;
assign F[7][47] = 9'b100111101;
assign F[7][48] = 9'b100111101;
assign F[7][49] = 9'b100111101;
assign F[7][50] = 9'b100111101;
assign F[7][51] = 9'b100011101;
assign F[7][52] = 9'b101111110;
assign F[7][53] = 9'b111111111;
assign F[7][54] = 9'b111111111;
assign F[7][55] = 9'b111111111;
assign F[7][56] = 9'b111111111;
assign F[7][57] = 9'b111111111;
assign F[7][58] = 9'b100111101;
assign F[7][59] = 9'b100111101;
assign F[7][60] = 9'b100111101;
assign F[8][41] = 9'b100111101;
assign F[8][42] = 9'b100111101;
assign F[8][43] = 9'b100111101;
assign F[8][44] = 9'b100111101;
assign F[8][45] = 9'b100111101;
assign F[8][46] = 9'b100111101;
assign F[8][47] = 9'b100111101;
assign F[8][48] = 9'b100111101;
assign F[8][49] = 9'b100111101;
assign F[8][50] = 9'b100111101;
assign F[8][51] = 9'b100011101;
assign F[8][52] = 9'b101111110;
assign F[8][53] = 9'b111111111;
assign F[8][54] = 9'b111111111;
assign F[8][55] = 9'b111111111;
assign F[8][56] = 9'b111111111;
assign F[8][57] = 9'b111111111;
assign F[8][58] = 9'b100111101;
assign F[8][59] = 9'b100111101;
assign F[8][60] = 9'b100111101;
assign F[8][61] = 9'b100111101;
assign F[9][41] = 9'b100111101;
assign F[9][42] = 9'b100111101;
assign F[9][43] = 9'b100111101;
assign F[9][44] = 9'b100111101;
assign F[9][45] = 9'b100111101;
assign F[9][46] = 9'b100111101;
assign F[9][47] = 9'b100111101;
assign F[9][48] = 9'b100111101;
assign F[9][49] = 9'b100111101;
assign F[9][50] = 9'b100111101;
assign F[9][51] = 9'b100111101;
assign F[9][52] = 9'b101011101;
assign F[9][53] = 9'b110011111;
assign F[9][54] = 9'b110011111;
assign F[9][55] = 9'b110011111;
assign F[9][56] = 9'b110011111;
assign F[9][57] = 9'b110011110;
assign F[9][58] = 9'b100111101;
assign F[9][59] = 9'b100111101;
assign F[9][60] = 9'b100111101;
assign F[9][61] = 9'b100111101;
assign F[9][62] = 9'b100111101;
assign F[10][41] = 9'b100111101;
assign F[10][42] = 9'b100111101;
assign F[10][43] = 9'b100111101;
assign F[10][44] = 9'b100111101;
assign F[10][45] = 9'b100111101;
assign F[10][46] = 9'b100111101;
assign F[10][47] = 9'b100111101;
assign F[10][48] = 9'b100111101;
assign F[10][49] = 9'b100111101;
assign F[10][50] = 9'b100111101;
assign F[10][51] = 9'b100111101;
assign F[10][52] = 9'b100111101;
assign F[10][53] = 9'b100011101;
assign F[10][54] = 9'b100011101;
assign F[10][55] = 9'b100011101;
assign F[10][56] = 9'b100111101;
assign F[10][57] = 9'b100111101;
assign F[10][58] = 9'b100111101;
assign F[10][59] = 9'b100111101;
assign F[10][60] = 9'b100111101;
assign F[10][61] = 9'b100111101;
assign F[10][62] = 9'b100111101;
assign F[11][41] = 9'b100111101;
assign F[11][42] = 9'b100111101;
assign F[11][43] = 9'b100111101;
assign F[11][44] = 9'b100111101;
assign F[11][45] = 9'b100111101;
assign F[11][46] = 9'b100111101;
assign F[11][47] = 9'b100111101;
assign F[11][48] = 9'b100111101;
assign F[11][49] = 9'b100111101;
assign F[11][50] = 9'b100111101;
assign F[11][51] = 9'b100111101;
assign F[11][52] = 9'b100110001;
assign F[11][53] = 9'b101101101;
assign F[11][54] = 9'b101111110;
assign F[11][55] = 9'b101011101;
assign F[11][56] = 9'b100111101;
assign F[11][57] = 9'b100111101;
assign F[11][58] = 9'b100111101;
assign F[11][59] = 9'b100111101;
assign F[11][60] = 9'b100111101;
assign F[11][61] = 9'b100111101;
assign F[12][41] = 9'b100111101;
assign F[12][42] = 9'b100111101;
assign F[12][43] = 9'b100111101;
assign F[12][44] = 9'b100111101;
assign F[12][45] = 9'b100111101;
assign F[12][46] = 9'b100111101;
assign F[12][47] = 9'b100111101;
assign F[12][48] = 9'b100111101;
assign F[12][49] = 9'b100111101;
assign F[12][50] = 9'b100111101;
assign F[12][51] = 9'b100111101;
assign F[12][52] = 9'b101001101;
assign F[12][53] = 9'b110000100;
assign F[12][54] = 9'b111111111;
assign F[12][55] = 9'b101011110;
assign F[12][56] = 9'b100011101;
assign F[12][57] = 9'b100111101;
assign F[12][58] = 9'b100111101;
assign F[12][59] = 9'b100111101;
assign F[12][60] = 9'b100111101;
assign F[12][61] = 9'b100111101;
assign F[12][62] = 9'b100111101;
assign F[13][41] = 9'b100111101;
assign F[13][42] = 9'b100111101;
assign F[13][43] = 9'b100111101;
assign F[13][44] = 9'b100111101;
assign F[13][45] = 9'b100111101;
assign F[13][46] = 9'b100111101;
assign F[13][47] = 9'b100111101;
assign F[13][48] = 9'b100111101;
assign F[13][49] = 9'b100111101;
assign F[13][50] = 9'b100111101;
assign F[13][51] = 9'b100111101;
assign F[13][52] = 9'b100111101;
assign F[13][53] = 9'b100110001;
assign F[13][54] = 9'b110000100;
assign F[13][55] = 9'b110000000;
assign F[13][56] = 9'b110001001;
assign F[13][57] = 9'b110111111;
assign F[13][58] = 9'b100111101;
assign F[13][59] = 9'b100111101;
assign F[13][60] = 9'b100111101;
assign F[13][61] = 9'b100111101;
assign F[13][62] = 9'b100111101;
assign F[13][63] = 9'b100111101;
assign F[14][41] = 9'b100111101;
assign F[14][42] = 9'b100111101;
assign F[14][43] = 9'b100110001;
assign F[14][44] = 9'b100110001;
assign F[14][45] = 9'b100110001;
assign F[14][46] = 9'b100111101;
assign F[14][47] = 9'b100111101;
assign F[14][48] = 9'b100111101;
assign F[14][49] = 9'b100111101;
assign F[14][50] = 9'b100111101;
assign F[14][51] = 9'b100111101;
assign F[14][52] = 9'b100111101;
assign F[14][53] = 9'b100111101;
assign F[14][54] = 9'b101001100;
assign F[14][55] = 9'b101101000;
assign F[14][56] = 9'b101101101;
assign F[14][57] = 9'b110011110;
assign F[14][58] = 9'b100111101;
assign F[14][59] = 9'b100111101;
assign F[14][60] = 9'b100111101;
assign F[14][61] = 9'b100111101;
assign F[14][62] = 9'b100111101;
assign F[14][63] = 9'b100111101;
assign F[14][64] = 9'b100111101;
assign F[14][65] = 9'b100111101;
assign F[15][41] = 9'b100111101;
assign F[15][42] = 9'b100111101;
assign F[15][43] = 9'b100100000;
assign F[15][44] = 9'b100100000;
assign F[15][45] = 9'b100101100;
assign F[15][46] = 9'b100111101;
assign F[15][47] = 9'b100011101;
assign F[15][48] = 9'b100111101;
assign F[15][49] = 9'b100111101;
assign F[15][50] = 9'b100111101;
assign F[15][51] = 9'b100111101;
assign F[15][52] = 9'b100111101;
assign F[15][53] = 9'b100111101;
assign F[15][54] = 9'b100111101;
assign F[15][55] = 9'b100011101;
assign F[15][56] = 9'b100011101;
assign F[15][57] = 9'b100011101;
assign F[15][58] = 9'b100011101;
assign F[15][59] = 9'b100011101;
assign F[15][60] = 9'b100011101;
assign F[15][61] = 9'b100011101;
assign F[15][62] = 9'b100011101;
assign F[15][63] = 9'b100111101;
assign F[15][64] = 9'b100111101;
assign F[15][65] = 9'b100111110;
assign F[15][66] = 9'b100111101;
assign F[16][41] = 9'b100110001;
assign F[16][42] = 9'b100101000;
assign F[16][43] = 9'b100100000;
assign F[16][44] = 9'b100100000;
assign F[16][45] = 9'b100100100;
assign F[16][46] = 9'b100101100;
assign F[16][47] = 9'b110010001;
assign F[16][48] = 9'b101010101;
assign F[16][49] = 9'b100111101;
assign F[16][50] = 9'b100111101;
assign F[16][51] = 9'b100111101;
assign F[16][52] = 9'b100111101;
assign F[16][53] = 9'b100111101;
assign F[16][54] = 9'b100111101;
assign F[16][55] = 9'b101010101;
assign F[16][56] = 9'b110010001;
assign F[16][57] = 9'b110010001;
assign F[16][58] = 9'b110010001;
assign F[16][59] = 9'b110010001;
assign F[16][60] = 9'b110010001;
assign F[16][61] = 9'b110010001;
assign F[16][62] = 9'b101101101;
assign F[16][63] = 9'b101101000;
assign F[16][64] = 9'b101101000;
assign F[16][65] = 9'b101101000;
assign F[16][66] = 9'b101001000;
assign F[17][41] = 9'b100101000;
assign F[17][42] = 9'b100100000;
assign F[17][43] = 9'b100100000;
assign F[17][44] = 9'b100100000;
assign F[17][45] = 9'b100100000;
assign F[17][46] = 9'b101000000;
assign F[17][47] = 9'b111101101;
assign F[17][48] = 9'b101010001;
assign F[17][49] = 9'b100011101;
assign F[17][50] = 9'b100110101;
assign F[17][51] = 9'b100110101;
assign F[17][52] = 9'b100110101;
assign F[17][53] = 9'b100110101;
assign F[17][54] = 9'b100011101;
assign F[17][55] = 9'b101110001;
assign F[17][56] = 9'b111101101;
assign F[17][57] = 9'b111101101;
assign F[17][58] = 9'b111101101;
assign F[17][59] = 9'b111101101;
assign F[17][60] = 9'b111101101;
assign F[17][61] = 9'b111101101;
assign F[17][62] = 9'b110100100;
assign F[17][63] = 9'b110000000;
assign F[17][64] = 9'b110000000;
assign F[17][65] = 9'b110100000;
assign F[17][66] = 9'b110000000;
assign F[18][40] = 9'b100100000;
assign F[18][41] = 9'b100100000;
assign F[18][42] = 9'b100100000;
assign F[18][43] = 9'b100100000;
assign F[18][44] = 9'b100100000;
assign F[18][45] = 9'b100100000;
assign F[18][46] = 9'b100000000;
assign F[18][47] = 9'b100000000;
assign F[18][48] = 9'b100000000;
assign F[18][49] = 9'b100000100;
assign F[18][50] = 9'b100000100;
assign F[18][51] = 9'b100000100;
assign F[18][52] = 9'b100000100;
assign F[18][53] = 9'b100000100;
assign F[18][54] = 9'b100000100;
assign F[18][55] = 9'b100000000;
assign F[18][56] = 9'b100000000;
assign F[18][57] = 9'b100100000;
assign F[18][58] = 9'b100100000;
assign F[18][59] = 9'b100100000;
assign F[18][60] = 9'b100100000;
assign F[18][61] = 9'b100000000;
assign F[18][62] = 9'b101100000;
assign F[18][63] = 9'b110100100;
assign F[18][64] = 9'b110000100;
assign F[18][65] = 9'b110100100;
assign F[18][66] = 9'b110000100;
assign F[19][39] = 9'b100100100;
assign F[19][40] = 9'b100100000;
assign F[19][41] = 9'b101000100;
assign F[19][42] = 9'b101101000;
assign F[19][43] = 9'b101101000;
assign F[19][44] = 9'b101000100;
assign F[19][45] = 9'b100100000;
assign F[19][46] = 9'b100100000;
assign F[19][47] = 9'b101000100;
assign F[19][48] = 9'b101000100;
assign F[19][49] = 9'b101000100;
assign F[19][50] = 9'b100000000;
assign F[19][51] = 9'b100000000;
assign F[19][52] = 9'b100000000;
assign F[19][53] = 9'b100000000;
assign F[19][54] = 9'b100000000;
assign F[19][55] = 9'b101000100;
assign F[19][56] = 9'b101000100;
assign F[19][57] = 9'b100000000;
assign F[19][58] = 9'b100000000;
assign F[19][59] = 9'b100000000;
assign F[19][60] = 9'b100000000;
assign F[19][61] = 9'b100000000;
assign F[19][62] = 9'b101000100;
assign F[19][63] = 9'b110000100;
assign F[19][64] = 9'b101100100;
assign F[19][65] = 9'b110000100;
assign F[20][38] = 9'b100100100;
assign F[20][39] = 9'b100100000;
assign F[20][40] = 9'b100100000;
assign F[20][41] = 9'b101101000;
assign F[20][42] = 9'b111110001;
assign F[20][43] = 9'b111110001;
assign F[20][44] = 9'b101000100;
assign F[20][45] = 9'b100100000;
assign F[20][46] = 9'b101000100;
assign F[20][47] = 9'b111110001;
assign F[20][48] = 9'b111110001;
assign F[20][49] = 9'b110001101;
assign F[20][50] = 9'b100000000;
assign F[20][51] = 9'b100000000;
assign F[20][52] = 9'b100000000;
assign F[20][53] = 9'b100000000;
assign F[20][54] = 9'b100000000;
assign F[20][55] = 9'b110001101;
assign F[20][56] = 9'b110001101;
assign F[20][57] = 9'b100000000;
assign F[20][58] = 9'b100000000;
assign F[20][59] = 9'b100000000;
assign F[20][60] = 9'b100000000;
assign F[20][61] = 9'b100000000;
assign F[21][38] = 9'b100100100;
assign F[21][39] = 9'b100100000;
assign F[21][40] = 9'b100100000;
assign F[21][41] = 9'b101101000;
assign F[21][42] = 9'b111110001;
assign F[21][43] = 9'b111110001;
assign F[21][44] = 9'b110101101;
assign F[21][45] = 9'b101101000;
assign F[21][46] = 9'b100100000;
assign F[21][47] = 9'b111101101;
assign F[21][48] = 9'b111110001;
assign F[21][49] = 9'b110001101;
assign F[21][50] = 9'b100000000;
assign F[21][51] = 9'b100000000;
assign F[21][52] = 9'b100000000;
assign F[21][53] = 9'b100000000;
assign F[21][54] = 9'b100000000;
assign F[21][55] = 9'b110001001;
assign F[21][56] = 9'b110001001;
assign F[21][57] = 9'b100000000;
assign F[21][58] = 9'b100000000;
assign F[21][59] = 9'b100000000;
assign F[21][60] = 9'b100000000;
assign F[21][61] = 9'b100000000;
assign F[22][38] = 9'b100100100;
assign F[22][39] = 9'b100100000;
assign F[22][40] = 9'b100100000;
assign F[22][41] = 9'b101101000;
assign F[22][42] = 9'b111110001;
assign F[22][43] = 9'b111110001;
assign F[22][44] = 9'b111110001;
assign F[22][45] = 9'b110001001;
assign F[22][46] = 9'b100100000;
assign F[22][47] = 9'b111101101;
assign F[22][48] = 9'b111110001;
assign F[22][49] = 9'b110001101;
assign F[22][50] = 9'b100100000;
assign F[22][51] = 9'b100100000;
assign F[22][52] = 9'b100100100;
assign F[22][53] = 9'b100100100;
assign F[22][54] = 9'b100100000;
assign F[22][55] = 9'b110001101;
assign F[22][56] = 9'b110001101;
assign F[22][57] = 9'b100100000;
assign F[22][58] = 9'b100100100;
assign F[22][59] = 9'b100100100;
assign F[22][60] = 9'b100100100;
assign F[22][61] = 9'b100100100;
assign F[23][38] = 9'b100100100;
assign F[23][39] = 9'b100100000;
assign F[23][40] = 9'b100100000;
assign F[23][41] = 9'b100100000;
assign F[23][42] = 9'b101000100;
assign F[23][43] = 9'b111110001;
assign F[23][44] = 9'b111110001;
assign F[23][45] = 9'b110001000;
assign F[23][46] = 9'b100100000;
assign F[23][47] = 9'b111101101;
assign F[23][48] = 9'b111110001;
assign F[23][49] = 9'b111110001;
assign F[23][50] = 9'b111101101;
assign F[23][51] = 9'b111101101;
assign F[23][52] = 9'b111101101;
assign F[23][53] = 9'b111101101;
assign F[23][54] = 9'b111101101;
assign F[23][55] = 9'b111110001;
assign F[23][56] = 9'b111101101;
assign F[23][57] = 9'b110101101;
assign F[23][58] = 9'b111101101;
assign F[23][59] = 9'b111101101;
assign F[23][60] = 9'b111110001;
assign F[23][61] = 9'b111110001;
assign F[24][38] = 9'b100100100;
assign F[24][39] = 9'b100100000;
assign F[24][40] = 9'b100100000;
assign F[24][41] = 9'b100100000;
assign F[24][42] = 9'b101000100;
assign F[24][43] = 9'b110001000;
assign F[24][44] = 9'b111101101;
assign F[24][45] = 9'b110001001;
assign F[24][46] = 9'b100100000;
assign F[24][47] = 9'b111101101;
assign F[24][48] = 9'b111110001;
assign F[24][49] = 9'b111110001;
assign F[24][50] = 9'b111110001;
assign F[24][51] = 9'b111110001;
assign F[24][52] = 9'b111110001;
assign F[24][53] = 9'b111110001;
assign F[24][54] = 9'b111110001;
assign F[24][55] = 9'b111110001;
assign F[24][56] = 9'b111110001;
assign F[24][57] = 9'b111101101;
assign F[24][58] = 9'b111110001;
assign F[24][59] = 9'b111110001;
assign F[24][60] = 9'b111110001;
assign F[24][61] = 9'b111110001;
assign F[25][38] = 9'b100100100;
assign F[25][39] = 9'b100100000;
assign F[25][40] = 9'b100100000;
assign F[25][41] = 9'b100100000;
assign F[25][42] = 9'b100100000;
assign F[25][43] = 9'b100100000;
assign F[25][44] = 9'b110001101;
assign F[25][45] = 9'b110001001;
assign F[25][46] = 9'b100100000;
assign F[25][47] = 9'b111101101;
assign F[25][48] = 9'b111110001;
assign F[25][49] = 9'b111110001;
assign F[25][50] = 9'b111110001;
assign F[25][51] = 9'b111110001;
assign F[25][52] = 9'b111110001;
assign F[25][53] = 9'b111110001;
assign F[25][54] = 9'b111110001;
assign F[25][55] = 9'b111110001;
assign F[25][56] = 9'b111110001;
assign F[25][57] = 9'b111101101;
assign F[25][58] = 9'b111110001;
assign F[25][59] = 9'b111110001;
assign F[25][60] = 9'b111110001;
assign F[25][61] = 9'b111110001;
assign F[26][38] = 9'b100100100;
assign F[26][39] = 9'b100100000;
assign F[26][40] = 9'b100100000;
assign F[26][41] = 9'b100100000;
assign F[26][42] = 9'b100100000;
assign F[26][43] = 9'b100100000;
assign F[26][44] = 9'b110001101;
assign F[26][45] = 9'b110101101;
assign F[26][46] = 9'b101101000;
assign F[26][47] = 9'b111110001;
assign F[26][48] = 9'b111110001;
assign F[26][49] = 9'b111110001;
assign F[26][50] = 9'b111110001;
assign F[26][51] = 9'b111110001;
assign F[26][52] = 9'b111110001;
assign F[26][53] = 9'b111110001;
assign F[26][54] = 9'b111110001;
assign F[26][55] = 9'b101001000;
assign F[26][56] = 9'b100100000;
assign F[26][57] = 9'b100100000;
assign F[26][58] = 9'b110101101;
assign F[26][59] = 9'b111110001;
assign F[26][60] = 9'b111110001;
assign F[26][61] = 9'b111110001;
assign F[27][39] = 9'b100100100;
assign F[27][40] = 9'b100100000;
assign F[27][41] = 9'b100100000;
assign F[27][42] = 9'b100100000;
assign F[27][43] = 9'b100100000;
assign F[27][44] = 9'b110001101;
assign F[27][45] = 9'b111101101;
assign F[27][46] = 9'b110001000;
assign F[27][47] = 9'b110101101;
assign F[27][48] = 9'b111110001;
assign F[27][49] = 9'b111110001;
assign F[27][50] = 9'b111110001;
assign F[27][51] = 9'b111110001;
assign F[27][52] = 9'b111110001;
assign F[27][53] = 9'b111110001;
assign F[27][54] = 9'b111110001;
assign F[27][55] = 9'b101000100;
assign F[27][56] = 9'b100000000;
assign F[27][57] = 9'b100000000;
assign F[27][58] = 9'b110101101;
assign F[27][59] = 9'b111110001;
assign F[27][60] = 9'b111110001;
assign F[27][61] = 9'b111110001;
assign F[28][40] = 9'b100100000;
assign F[28][41] = 9'b100100000;
assign F[28][42] = 9'b100100000;
assign F[28][43] = 9'b100100000;
assign F[28][44] = 9'b110001101;
assign F[28][45] = 9'b111101101;
assign F[28][46] = 9'b110001000;
assign F[28][47] = 9'b110001000;
assign F[28][48] = 9'b110101101;
assign F[28][49] = 9'b111110001;
assign F[28][50] = 9'b111110001;
assign F[28][51] = 9'b111110001;
assign F[28][52] = 9'b111110001;
assign F[28][53] = 9'b111110001;
assign F[28][54] = 9'b111110001;
assign F[28][55] = 9'b111110001;
assign F[28][56] = 9'b111110001;
assign F[28][57] = 9'b111110001;
assign F[28][58] = 9'b111110001;
assign F[28][59] = 9'b111110001;
assign F[28][60] = 9'b111110001;
assign F[28][61] = 9'b111110001;
assign F[29][40] = 9'b100100100;
assign F[29][41] = 9'b100100000;
assign F[29][42] = 9'b100100000;
assign F[29][43] = 9'b100100000;
assign F[29][44] = 9'b110001101;
assign F[29][45] = 9'b110101101;
assign F[29][46] = 9'b110001000;
assign F[29][47] = 9'b110001000;
assign F[29][48] = 9'b110001000;
assign F[29][49] = 9'b110101101;
assign F[29][50] = 9'b111110001;
assign F[29][51] = 9'b111110001;
assign F[29][52] = 9'b110101101;
assign F[29][53] = 9'b110001101;
assign F[29][54] = 9'b110101101;
assign F[29][55] = 9'b110101101;
assign F[29][56] = 9'b110101101;
assign F[29][57] = 9'b110101101;
assign F[29][58] = 9'b110101101;
assign F[29][59] = 9'b110001101;
assign F[29][60] = 9'b110101101;
assign F[29][61] = 9'b111110001;
assign F[30][41] = 9'b100100100;
assign F[30][42] = 9'b100100000;
assign F[30][43] = 9'b100100000;
assign F[30][44] = 9'b110001101;
assign F[30][45] = 9'b111101101;
assign F[30][46] = 9'b110001000;
assign F[30][47] = 9'b110001000;
assign F[30][48] = 9'b110001000;
assign F[30][49] = 9'b110001000;
assign F[30][50] = 9'b111110001;
assign F[30][51] = 9'b111110001;
assign F[30][52] = 9'b110101101;
assign F[30][53] = 9'b101101000;
assign F[30][54] = 9'b110001000;
assign F[30][55] = 9'b110001000;
assign F[30][56] = 9'b110001000;
assign F[30][57] = 9'b110001000;
assign F[30][58] = 9'b110001000;
assign F[30][59] = 9'b110001000;
assign F[30][60] = 9'b110001000;
assign F[30][61] = 9'b111110001;
assign F[31][42] = 9'b100100100;
assign F[31][43] = 9'b100100000;
assign F[31][44] = 9'b110001101;
assign F[31][45] = 9'b111110001;
assign F[31][46] = 9'b110101101;
assign F[31][47] = 9'b110001000;
assign F[31][48] = 9'b110001000;
assign F[31][49] = 9'b110001000;
assign F[31][50] = 9'b110001000;
assign F[31][51] = 9'b111110001;
assign F[31][52] = 9'b110101101;
assign F[31][53] = 9'b101101000;
assign F[31][54] = 9'b100000000;
assign F[31][55] = 9'b100000000;
assign F[31][56] = 9'b100000000;
assign F[31][57] = 9'b100000000;
assign F[31][58] = 9'b100000000;
assign F[31][59] = 9'b101000100;
assign F[31][60] = 9'b110001001;
assign F[31][61] = 9'b111110001;
assign F[32][43] = 9'b100100000;
assign F[32][44] = 9'b110001101;
assign F[32][45] = 9'b111110001;
assign F[32][46] = 9'b111110001;
assign F[32][47] = 9'b110001001;
assign F[32][48] = 9'b110001000;
assign F[32][49] = 9'b110001000;
assign F[32][50] = 9'b110001000;
assign F[32][51] = 9'b110101101;
assign F[32][52] = 9'b110101101;
assign F[32][53] = 9'b101101000;
assign F[32][54] = 9'b100100000;
assign F[32][55] = 9'b100000000;
assign F[32][56] = 9'b100000000;
assign F[32][57] = 9'b100000000;
assign F[32][58] = 9'b100100000;
assign F[32][59] = 9'b101000100;
assign F[32][60] = 9'b110001000;
assign F[32][61] = 9'b111101101;
assign F[32][62] = 9'b110001101;
assign F[33][43] = 9'b100100000;
assign F[33][44] = 9'b110001101;
assign F[33][45] = 9'b111110001;
assign F[33][46] = 9'b111110001;
assign F[33][47] = 9'b111110001;
assign F[33][48] = 9'b110001101;
assign F[33][49] = 9'b101101000;
assign F[33][50] = 9'b110001000;
assign F[33][51] = 9'b110001000;
assign F[33][52] = 9'b110001000;
assign F[33][53] = 9'b110001000;
assign F[33][54] = 9'b111110001;
assign F[33][55] = 9'b110001101;
assign F[33][56] = 9'b110001000;
assign F[33][57] = 9'b110001000;
assign F[33][58] = 9'b111110001;
assign F[33][59] = 9'b110101101;
assign F[33][60] = 9'b110001000;
assign F[33][61] = 9'b110001000;
assign F[34][43] = 9'b100100000;
assign F[34][44] = 9'b110101101;
assign F[34][45] = 9'b111110001;
assign F[34][46] = 9'b111110001;
assign F[34][47] = 9'b111110001;
assign F[34][48] = 9'b110101101;
assign F[34][49] = 9'b110001101;
assign F[34][50] = 9'b110001000;
assign F[34][51] = 9'b110001000;
assign F[34][52] = 9'b110001000;
assign F[34][53] = 9'b110001000;
assign F[34][54] = 9'b111110001;
assign F[34][55] = 9'b110101101;
assign F[34][56] = 9'b110101101;
assign F[34][57] = 9'b110101101;
assign F[34][58] = 9'b111110001;
assign F[34][59] = 9'b110101101;
assign F[34][60] = 9'b110001000;
assign F[34][61] = 9'b110001000;
assign F[35][44] = 9'b111110001;
assign F[35][45] = 9'b111110001;
assign F[35][46] = 9'b111110001;
assign F[35][47] = 9'b111110001;
assign F[35][48] = 9'b111110001;
assign F[35][49] = 9'b111101101;
assign F[35][50] = 9'b110001000;
assign F[35][51] = 9'b110001000;
assign F[35][52] = 9'b110001000;
assign F[35][53] = 9'b110001000;
assign F[35][54] = 9'b111101101;
assign F[35][55] = 9'b111110001;
assign F[35][56] = 9'b111110001;
assign F[35][57] = 9'b111110001;
assign F[35][58] = 9'b111110001;
assign F[35][59] = 9'b110001101;
assign F[35][60] = 9'b110001000;
assign F[35][61] = 9'b110001000;
assign F[36][44] = 9'b111110001;
assign F[36][45] = 9'b111110001;
assign F[36][46] = 9'b111110001;
assign F[36][47] = 9'b111110001;
assign F[36][48] = 9'b111110001;
assign F[36][49] = 9'b111110001;
assign F[36][50] = 9'b111101101;
assign F[36][51] = 9'b110001000;
assign F[36][52] = 9'b110001000;
assign F[36][53] = 9'b110001000;
assign F[36][54] = 9'b110001000;
assign F[36][55] = 9'b110001000;
assign F[36][56] = 9'b110001000;
assign F[36][57] = 9'b110001000;
assign F[36][58] = 9'b110001000;
assign F[36][59] = 9'b110001000;
assign F[36][60] = 9'b110001000;
assign F[37][44] = 9'b111110001;
assign F[37][45] = 9'b111110001;
assign F[37][46] = 9'b111110001;
assign F[37][47] = 9'b111110001;
assign F[37][48] = 9'b111110001;
assign F[37][49] = 9'b111110001;
assign F[37][50] = 9'b111110001;
assign F[37][51] = 9'b110001101;
assign F[37][52] = 9'b110001000;
assign F[37][53] = 9'b110001000;
assign F[37][54] = 9'b110001000;
assign F[37][55] = 9'b110001000;
assign F[37][56] = 9'b110001000;
assign F[37][57] = 9'b110001000;
assign F[37][58] = 9'b101101000;
assign F[37][59] = 9'b110001000;
assign F[37][60] = 9'b101101000;
assign F[38][44] = 9'b111110001;
assign F[38][45] = 9'b111110001;
assign F[38][46] = 9'b111110001;
assign F[38][47] = 9'b111110001;
assign F[38][48] = 9'b111110001;
assign F[38][49] = 9'b111110001;
assign F[38][50] = 9'b111110001;
assign F[38][51] = 9'b111110001;
assign F[38][52] = 9'b111110001;
assign F[38][53] = 9'b111110001;
assign F[38][54] = 9'b111110001;
assign F[38][55] = 9'b111110001;
assign F[38][56] = 9'b111110001;
assign F[38][57] = 9'b111110001;
assign F[39][43] = 9'b100110001;
assign F[39][44] = 9'b101010001;
assign F[39][45] = 9'b101010001;
assign F[39][46] = 9'b101010001;
assign F[39][47] = 9'b101010001;
assign F[39][48] = 9'b101110001;
assign F[39][49] = 9'b110001101;
assign F[39][50] = 9'b111101101;
assign F[39][51] = 9'b111101101;
assign F[39][52] = 9'b111101101;
assign F[39][53] = 9'b110101101;
assign F[39][54] = 9'b101010001;
assign F[39][55] = 9'b101010001;
assign F[39][56] = 9'b101010001;
assign F[39][57] = 9'b101010001;
assign F[39][58] = 9'b100110101;
assign F[39][59] = 9'b100110001;
assign F[40][43] = 9'b100110101;
assign F[40][44] = 9'b100010101;
assign F[40][45] = 9'b100010001;
assign F[40][46] = 9'b100010101;
assign F[40][47] = 9'b100010101;
assign F[40][48] = 9'b100110001;
assign F[40][49] = 9'b101001101;
assign F[40][50] = 9'b110001001;
assign F[40][51] = 9'b110001001;
assign F[40][52] = 9'b110001001;
assign F[40][53] = 9'b110001101;
assign F[40][54] = 9'b100010001;
assign F[40][55] = 9'b100010101;
assign F[40][56] = 9'b100010101;
assign F[40][57] = 9'b100010101;
assign F[40][58] = 9'b100111101;
assign F[40][59] = 9'b100110001;
assign F[41][37] = 9'b100001111;
assign F[41][38] = 9'b100010010;
assign F[41][39] = 9'b100110001;
assign F[41][40] = 9'b100110001;
assign F[41][41] = 9'b100110001;
assign F[41][42] = 9'b100110001;
assign F[41][43] = 9'b100110001;
assign F[41][44] = 9'b100110001;
assign F[41][45] = 9'b100110001;
assign F[41][46] = 9'b100110001;
assign F[41][47] = 9'b100110001;
assign F[41][48] = 9'b100110001;
assign F[41][49] = 9'b100110001;
assign F[41][50] = 9'b100110001;
assign F[41][51] = 9'b100110001;
assign F[41][52] = 9'b100110001;
assign F[41][53] = 9'b100110001;
assign F[41][54] = 9'b100110001;
assign F[41][55] = 9'b100110001;
assign F[41][56] = 9'b100110001;
assign F[41][57] = 9'b100110001;
assign F[41][58] = 9'b100110001;
assign F[41][59] = 9'b100110001;
assign F[41][60] = 9'b100110001;
assign F[41][61] = 9'b100110001;
assign F[41][62] = 9'b100110101;
assign F[41][63] = 9'b100010001;
assign F[41][64] = 9'b100001111;
assign F[42][37] = 9'b100001111;
assign F[42][38] = 9'b100010011;
assign F[42][39] = 9'b100110101;
assign F[42][40] = 9'b100110101;
assign F[42][41] = 9'b100110101;
assign F[42][42] = 9'b100110101;
assign F[42][43] = 9'b100110001;
assign F[42][44] = 9'b100110001;
assign F[42][45] = 9'b100110001;
assign F[42][46] = 9'b100110001;
assign F[42][47] = 9'b100110001;
assign F[42][48] = 9'b100110001;
assign F[42][49] = 9'b100110001;
assign F[42][50] = 9'b100110001;
assign F[42][51] = 9'b100110001;
assign F[42][52] = 9'b100110001;
assign F[42][53] = 9'b100110001;
assign F[42][54] = 9'b100110001;
assign F[42][55] = 9'b100110001;
assign F[42][56] = 9'b100110001;
assign F[42][57] = 9'b100110001;
assign F[42][58] = 9'b100110001;
assign F[42][59] = 9'b100110101;
assign F[42][60] = 9'b100110101;
assign F[42][61] = 9'b100110101;
assign F[42][62] = 9'b100110101;
assign F[42][63] = 9'b100010001;
assign F[42][64] = 9'b100001111;
assign F[43][37] = 9'b100001111;
assign F[43][38] = 9'b100010010;
assign F[43][39] = 9'b100110101;
assign F[43][40] = 9'b100110001;
assign F[43][41] = 9'b100110001;
assign F[43][42] = 9'b100110001;
assign F[43][43] = 9'b100110001;
assign F[43][44] = 9'b100110001;
assign F[43][45] = 9'b100110001;
assign F[43][46] = 9'b100110001;
assign F[43][47] = 9'b100110001;
assign F[43][48] = 9'b100110001;
assign F[43][49] = 9'b100110001;
assign F[43][50] = 9'b100110001;
assign F[43][51] = 9'b100110001;
assign F[43][52] = 9'b100110001;
assign F[43][53] = 9'b100110001;
assign F[43][54] = 9'b100110001;
assign F[43][55] = 9'b100110001;
assign F[43][56] = 9'b100110001;
assign F[43][57] = 9'b100110001;
assign F[43][58] = 9'b100110101;
assign F[43][59] = 9'b100110101;
assign F[43][60] = 9'b100110001;
assign F[43][61] = 9'b100110001;
assign F[43][62] = 9'b100110101;
assign F[43][63] = 9'b100010001;
assign F[43][64] = 9'b100001111;
assign F[44][37] = 9'b100001111;
assign F[44][38] = 9'b100010011;
assign F[44][39] = 9'b100110101;
assign F[44][40] = 9'b100110101;
assign F[44][41] = 9'b100110101;
assign F[44][42] = 9'b100110101;
assign F[44][43] = 9'b100110101;
assign F[44][44] = 9'b100110101;
assign F[44][45] = 9'b100110101;
assign F[44][46] = 9'b100110101;
assign F[44][47] = 9'b100110101;
assign F[44][48] = 9'b100110101;
assign F[44][49] = 9'b100110101;
assign F[44][50] = 9'b100110101;
assign F[44][51] = 9'b100110101;
assign F[44][52] = 9'b100110101;
assign F[44][53] = 9'b100110101;
assign F[44][54] = 9'b100110101;
assign F[44][55] = 9'b100110101;
assign F[44][56] = 9'b100110101;
assign F[44][57] = 9'b100110101;
assign F[44][58] = 9'b100110001;
assign F[44][59] = 9'b100110001;
assign F[44][60] = 9'b100110101;
assign F[44][61] = 9'b100110101;
assign F[44][62] = 9'b100110101;
assign F[44][63] = 9'b100010001;
assign F[44][64] = 9'b100001111;
assign F[45][37] = 9'b100001111;
assign F[45][38] = 9'b100010010;
assign F[45][39] = 9'b100110101;
assign F[45][40] = 9'b100110001;
assign F[45][41] = 9'b100110001;
assign F[45][42] = 9'b100110001;
assign F[45][43] = 9'b100110001;
assign F[45][44] = 9'b100110001;
assign F[45][45] = 9'b100110001;
assign F[45][46] = 9'b100110001;
assign F[45][47] = 9'b100110001;
assign F[45][48] = 9'b100110001;
assign F[45][49] = 9'b100110001;
assign F[45][50] = 9'b100110001;
assign F[45][51] = 9'b100110001;
assign F[45][52] = 9'b100110001;
assign F[45][53] = 9'b100110001;
assign F[45][54] = 9'b100110001;
assign F[45][55] = 9'b100110001;
assign F[45][56] = 9'b100110101;
assign F[45][57] = 9'b100110001;
assign F[45][59] = 9'b100110001;
assign F[45][60] = 9'b100110101;
assign F[45][61] = 9'b100110001;
assign F[45][62] = 9'b100110101;
assign F[45][63] = 9'b100010001;
assign F[45][64] = 9'b100001111;
//Total de Lineas = 937
endmodule






