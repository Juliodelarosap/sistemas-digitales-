`timescale 1ns / 1ps
module prueba_1 (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (micromat[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= micromat[vcount- posy][hcount- posx][7:5];
				green <= micromat[vcount- posy][hcount- posx][4:2];
            blue 	<= micromat[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 100;
parameter RESOLUCION_Y = 100;
wire [8:0] micromat[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign micromat[0][0] = 9'b111111111;
assign micromat[0][1] = 9'b111111111;
assign micromat[0][2] = 9'b111111111;
assign micromat[0][3] = 9'b111111111;
assign micromat[0][4] = 9'b111111111;
assign micromat[0][5] = 9'b111111111;
assign micromat[0][6] = 9'b111111111;
assign micromat[0][7] = 9'b111111111;
assign micromat[0][8] = 9'b111111111;
assign micromat[0][9] = 9'b111111111;
assign micromat[0][10] = 9'b111111111;
assign micromat[0][11] = 9'b111111111;
assign micromat[0][12] = 9'b111111111;
assign micromat[0][13] = 9'b111111111;
assign micromat[0][14] = 9'b111111111;
assign micromat[0][15] = 9'b111111111;
assign micromat[0][16] = 9'b111111111;
assign micromat[0][17] = 9'b111111111;
assign micromat[0][18] = 9'b111111111;
assign micromat[0][19] = 9'b111111111;
assign micromat[0][20] = 9'b111111111;
assign micromat[0][21] = 9'b111111111;
assign micromat[0][22] = 9'b111111111;
assign micromat[0][23] = 9'b111111111;
assign micromat[0][24] = 9'b111111111;
assign micromat[0][25] = 9'b111111111;
assign micromat[0][26] = 9'b111111111;
assign micromat[0][27] = 9'b111111111;
assign micromat[0][28] = 9'b111111111;
assign micromat[0][29] = 9'b111111111;
assign micromat[0][30] = 9'b111111111;
assign micromat[0][31] = 9'b111111111;
assign micromat[0][32] = 9'b111111111;
assign micromat[0][33] = 9'b111111111;
assign micromat[0][34] = 9'b111111111;
assign micromat[0][35] = 9'b111111111;
assign micromat[0][36] = 9'b111111111;
assign micromat[0][37] = 9'b111111111;
assign micromat[0][38] = 9'b111111111;
assign micromat[0][39] = 9'b111111111;
assign micromat[0][40] = 9'b111111111;
assign micromat[0][41] = 9'b111111111;
assign micromat[0][42] = 9'b111111111;
assign micromat[0][43] = 9'b111111111;
assign micromat[0][44] = 9'b111111111;
assign micromat[0][45] = 9'b111111111;
assign micromat[0][46] = 9'b111111111;
assign micromat[0][47] = 9'b111111111;
assign micromat[0][48] = 9'b111111111;
assign micromat[0][49] = 9'b111111111;
assign micromat[0][50] = 9'b111111111;
assign micromat[0][51] = 9'b111111111;
assign micromat[0][52] = 9'b111111111;
assign micromat[0][53] = 9'b111111111;
assign micromat[0][54] = 9'b111111111;
assign micromat[0][55] = 9'b111111111;
assign micromat[0][56] = 9'b111111111;
assign micromat[0][57] = 9'b111111111;
assign micromat[0][58] = 9'b111111111;
assign micromat[0][59] = 9'b111111111;
assign micromat[0][60] = 9'b111111111;
assign micromat[0][61] = 9'b111111111;
assign micromat[0][62] = 9'b111111111;
assign micromat[0][63] = 9'b111111111;
assign micromat[0][64] = 9'b111111111;
assign micromat[0][65] = 9'b111111111;
assign micromat[0][66] = 9'b111111111;
assign micromat[0][67] = 9'b111111111;
assign micromat[0][68] = 9'b111111111;
assign micromat[0][69] = 9'b111111111;
assign micromat[0][70] = 9'b111111111;
assign micromat[0][71] = 9'b111111111;
assign micromat[0][72] = 9'b111111111;
assign micromat[0][73] = 9'b111111111;
assign micromat[0][74] = 9'b111111111;
assign micromat[0][75] = 9'b111111111;
assign micromat[0][76] = 9'b111111111;
assign micromat[0][77] = 9'b111111111;
assign micromat[0][78] = 9'b111111111;
assign micromat[0][79] = 9'b111111111;
assign micromat[0][80] = 9'b111111111;
assign micromat[0][81] = 9'b111111111;
assign micromat[0][82] = 9'b111111111;
assign micromat[0][83] = 9'b111111111;
assign micromat[0][84] = 9'b111111111;
assign micromat[0][85] = 9'b111111111;
assign micromat[0][86] = 9'b111111111;
assign micromat[0][87] = 9'b111111111;
assign micromat[0][88] = 9'b111111111;
assign micromat[0][89] = 9'b111111111;
assign micromat[0][90] = 9'b111111111;
assign micromat[0][91] = 9'b111111111;
assign micromat[0][92] = 9'b111111111;
assign micromat[0][93] = 9'b111111111;
assign micromat[0][94] = 9'b111111111;
assign micromat[0][95] = 9'b111111111;
assign micromat[0][96] = 9'b111111111;
assign micromat[0][97] = 9'b111111111;
assign micromat[0][98] = 9'b111111111;
assign micromat[0][99] = 9'b111111111;
assign micromat[1][0] = 9'b111111111;
assign micromat[1][1] = 9'b111111111;
assign micromat[1][2] = 9'b111111111;
assign micromat[1][3] = 9'b111111111;
assign micromat[1][4] = 9'b111111111;
assign micromat[1][5] = 9'b111111111;
assign micromat[1][6] = 9'b111111111;
assign micromat[1][7] = 9'b111111111;
assign micromat[1][8] = 9'b111111111;
assign micromat[1][9] = 9'b111111111;
assign micromat[1][10] = 9'b111111111;
assign micromat[1][11] = 9'b111111111;
assign micromat[1][12] = 9'b111111111;
assign micromat[1][13] = 9'b111111111;
assign micromat[1][14] = 9'b111111111;
assign micromat[1][15] = 9'b111111111;
assign micromat[1][16] = 9'b111111111;
assign micromat[1][17] = 9'b111111111;
assign micromat[1][18] = 9'b111111111;
assign micromat[1][19] = 9'b111111111;
assign micromat[1][20] = 9'b111111111;
assign micromat[1][21] = 9'b111111111;
assign micromat[1][22] = 9'b111111111;
assign micromat[1][23] = 9'b111111111;
assign micromat[1][24] = 9'b111111111;
assign micromat[1][25] = 9'b111111111;
assign micromat[1][26] = 9'b111111111;
assign micromat[1][27] = 9'b111111111;
assign micromat[1][28] = 9'b111111111;
assign micromat[1][29] = 9'b111111111;
assign micromat[1][30] = 9'b111111111;
assign micromat[1][31] = 9'b111111111;
assign micromat[1][32] = 9'b111111111;
assign micromat[1][33] = 9'b111111111;
assign micromat[1][34] = 9'b111111111;
assign micromat[1][35] = 9'b111111111;
assign micromat[1][36] = 9'b111111111;
assign micromat[1][37] = 9'b111111111;
assign micromat[1][38] = 9'b111111111;
assign micromat[1][39] = 9'b111111111;
assign micromat[1][40] = 9'b111111111;
assign micromat[1][41] = 9'b111111111;
assign micromat[1][42] = 9'b111111111;
assign micromat[1][43] = 9'b111111111;
assign micromat[1][44] = 9'b111111111;
assign micromat[1][45] = 9'b111111111;
assign micromat[1][46] = 9'b111111111;
assign micromat[1][47] = 9'b111111111;
assign micromat[1][48] = 9'b111111111;
assign micromat[1][49] = 9'b111111111;
assign micromat[1][50] = 9'b111111111;
assign micromat[1][51] = 9'b111111111;
assign micromat[1][52] = 9'b111111111;
assign micromat[1][53] = 9'b111111111;
assign micromat[1][54] = 9'b111111111;
assign micromat[1][55] = 9'b111111111;
assign micromat[1][56] = 9'b111111111;
assign micromat[1][57] = 9'b111111111;
assign micromat[1][58] = 9'b111111111;
assign micromat[1][59] = 9'b111111111;
assign micromat[1][60] = 9'b111111111;
assign micromat[1][61] = 9'b111111111;
assign micromat[1][62] = 9'b111111111;
assign micromat[1][63] = 9'b111111111;
assign micromat[1][64] = 9'b111111111;
assign micromat[1][65] = 9'b111111111;
assign micromat[1][66] = 9'b111111111;
assign micromat[1][67] = 9'b111111111;
assign micromat[1][68] = 9'b111111111;
assign micromat[1][69] = 9'b111111111;
assign micromat[1][70] = 9'b111111111;
assign micromat[1][71] = 9'b111111111;
assign micromat[1][72] = 9'b111111111;
assign micromat[1][73] = 9'b111111111;
assign micromat[1][74] = 9'b111111111;
assign micromat[1][75] = 9'b111111111;
assign micromat[1][76] = 9'b111111111;
assign micromat[1][77] = 9'b111111111;
assign micromat[1][78] = 9'b111111111;
assign micromat[1][79] = 9'b111111111;
assign micromat[1][80] = 9'b111111111;
assign micromat[1][81] = 9'b111111111;
assign micromat[1][82] = 9'b111111111;
assign micromat[1][83] = 9'b111111111;
assign micromat[1][84] = 9'b111111111;
assign micromat[1][85] = 9'b111111111;
assign micromat[1][86] = 9'b111111111;
assign micromat[1][87] = 9'b111111111;
assign micromat[1][88] = 9'b111111111;
assign micromat[1][89] = 9'b111111111;
assign micromat[1][90] = 9'b111111111;
assign micromat[1][91] = 9'b111111111;
assign micromat[1][92] = 9'b111111111;
assign micromat[1][93] = 9'b111111111;
assign micromat[1][94] = 9'b111111111;
assign micromat[1][95] = 9'b111111111;
assign micromat[1][96] = 9'b111111111;
assign micromat[1][97] = 9'b111111111;
assign micromat[1][98] = 9'b111111111;
assign micromat[1][99] = 9'b111111111;
assign micromat[2][0] = 9'b111111111;
assign micromat[2][1] = 9'b111111111;
assign micromat[2][2] = 9'b111111111;
assign micromat[2][3] = 9'b111111111;
assign micromat[2][4] = 9'b111111111;
assign micromat[2][5] = 9'b111111111;
assign micromat[2][6] = 9'b111111111;
assign micromat[2][7] = 9'b111111111;
assign micromat[2][8] = 9'b111111111;
assign micromat[2][9] = 9'b111111111;
assign micromat[2][10] = 9'b111111111;
assign micromat[2][11] = 9'b111111111;
assign micromat[2][12] = 9'b111111111;
assign micromat[2][13] = 9'b111111111;
assign micromat[2][14] = 9'b111111111;
assign micromat[2][15] = 9'b111111111;
assign micromat[2][16] = 9'b111111111;
assign micromat[2][17] = 9'b111111111;
assign micromat[2][18] = 9'b111111111;
assign micromat[2][19] = 9'b111111111;
assign micromat[2][20] = 9'b111111111;
assign micromat[2][21] = 9'b111111111;
assign micromat[2][22] = 9'b111111111;
assign micromat[2][23] = 9'b111111111;
assign micromat[2][24] = 9'b111111111;
assign micromat[2][25] = 9'b111111111;
assign micromat[2][26] = 9'b111111111;
assign micromat[2][27] = 9'b111111111;
assign micromat[2][28] = 9'b111111111;
assign micromat[2][29] = 9'b111111111;
assign micromat[2][30] = 9'b111111111;
assign micromat[2][31] = 9'b111111111;
assign micromat[2][32] = 9'b111111111;
assign micromat[2][33] = 9'b111111111;
assign micromat[2][34] = 9'b111111111;
assign micromat[2][35] = 9'b111111111;
assign micromat[2][36] = 9'b111111111;
assign micromat[2][37] = 9'b111111111;
assign micromat[2][38] = 9'b111111111;
assign micromat[2][39] = 9'b111111111;
assign micromat[2][40] = 9'b111111111;
assign micromat[2][41] = 9'b111111111;
assign micromat[2][42] = 9'b111111111;
assign micromat[2][43] = 9'b111111111;
assign micromat[2][44] = 9'b111111111;
assign micromat[2][45] = 9'b111111111;
assign micromat[2][46] = 9'b111111111;
assign micromat[2][47] = 9'b111111111;
assign micromat[2][48] = 9'b111111111;
assign micromat[2][49] = 9'b111111111;
assign micromat[2][50] = 9'b111111111;
assign micromat[2][51] = 9'b111111111;
assign micromat[2][52] = 9'b111111111;
assign micromat[2][53] = 9'b111111111;
assign micromat[2][54] = 9'b111111111;
assign micromat[2][55] = 9'b111111111;
assign micromat[2][56] = 9'b111111111;
assign micromat[2][57] = 9'b111111111;
assign micromat[2][58] = 9'b111111111;
assign micromat[2][59] = 9'b111111111;
assign micromat[2][60] = 9'b111111111;
assign micromat[2][61] = 9'b111111111;
assign micromat[2][62] = 9'b111111111;
assign micromat[2][63] = 9'b111111111;
assign micromat[2][64] = 9'b111111111;
assign micromat[2][65] = 9'b111111111;
assign micromat[2][66] = 9'b111111111;
assign micromat[2][67] = 9'b111111111;
assign micromat[2][68] = 9'b111111111;
assign micromat[2][69] = 9'b111111111;
assign micromat[2][70] = 9'b111111111;
assign micromat[2][71] = 9'b111111111;
assign micromat[2][72] = 9'b111111111;
assign micromat[2][73] = 9'b111111111;
assign micromat[2][74] = 9'b111111111;
assign micromat[2][75] = 9'b111111111;
assign micromat[2][76] = 9'b111111111;
assign micromat[2][77] = 9'b111111111;
assign micromat[2][78] = 9'b111111111;
assign micromat[2][79] = 9'b111111111;
assign micromat[2][80] = 9'b111111111;
assign micromat[2][81] = 9'b111111111;
assign micromat[2][82] = 9'b111111111;
assign micromat[2][83] = 9'b111111111;
assign micromat[2][84] = 9'b111111111;
assign micromat[2][85] = 9'b111111111;
assign micromat[2][86] = 9'b111111111;
assign micromat[2][87] = 9'b111111111;
assign micromat[2][88] = 9'b111111111;
assign micromat[2][89] = 9'b111111111;
assign micromat[2][90] = 9'b111111111;
assign micromat[2][91] = 9'b111111111;
assign micromat[2][92] = 9'b111111111;
assign micromat[2][93] = 9'b111111111;
assign micromat[2][94] = 9'b111111111;
assign micromat[2][95] = 9'b111111111;
assign micromat[2][96] = 9'b111111111;
assign micromat[2][97] = 9'b111111111;
assign micromat[2][98] = 9'b111111111;
assign micromat[2][99] = 9'b111111111;
assign micromat[3][0] = 9'b111111111;
assign micromat[3][1] = 9'b111111111;
assign micromat[3][2] = 9'b111111111;
assign micromat[3][3] = 9'b111111111;
assign micromat[3][4] = 9'b111111111;
assign micromat[3][5] = 9'b111111111;
assign micromat[3][6] = 9'b111111111;
assign micromat[3][7] = 9'b111111111;
assign micromat[3][8] = 9'b111111111;
assign micromat[3][9] = 9'b111111111;
assign micromat[3][10] = 9'b111111111;
assign micromat[3][11] = 9'b111111111;
assign micromat[3][12] = 9'b111111111;
assign micromat[3][13] = 9'b111111111;
assign micromat[3][14] = 9'b111111111;
assign micromat[3][15] = 9'b111111111;
assign micromat[3][16] = 9'b111111111;
assign micromat[3][17] = 9'b111111111;
assign micromat[3][18] = 9'b111111111;
assign micromat[3][19] = 9'b111111111;
assign micromat[3][20] = 9'b111111111;
assign micromat[3][21] = 9'b111111111;
assign micromat[3][22] = 9'b111111111;
assign micromat[3][23] = 9'b111111111;
assign micromat[3][24] = 9'b111111111;
assign micromat[3][25] = 9'b111111111;
assign micromat[3][26] = 9'b111111111;
assign micromat[3][27] = 9'b111111111;
assign micromat[3][28] = 9'b111111111;
assign micromat[3][29] = 9'b111111111;
assign micromat[3][30] = 9'b111111111;
assign micromat[3][31] = 9'b111111111;
assign micromat[3][32] = 9'b111111111;
assign micromat[3][33] = 9'b111111111;
assign micromat[3][34] = 9'b111111111;
assign micromat[3][35] = 9'b111111111;
assign micromat[3][36] = 9'b111111111;
assign micromat[3][37] = 9'b111111111;
assign micromat[3][38] = 9'b111111111;
assign micromat[3][39] = 9'b111111111;
assign micromat[3][40] = 9'b111111111;
assign micromat[3][41] = 9'b111111111;
assign micromat[3][42] = 9'b111111111;
assign micromat[3][43] = 9'b111111111;
assign micromat[3][44] = 9'b111111111;
assign micromat[3][45] = 9'b111111111;
assign micromat[3][46] = 9'b111111111;
assign micromat[3][47] = 9'b111111111;
assign micromat[3][48] = 9'b111111111;
assign micromat[3][49] = 9'b111111111;
assign micromat[3][50] = 9'b111111111;
assign micromat[3][51] = 9'b111111111;
assign micromat[3][52] = 9'b111111111;
assign micromat[3][53] = 9'b111111111;
assign micromat[3][54] = 9'b111111111;
assign micromat[3][55] = 9'b111111111;
assign micromat[3][56] = 9'b111111111;
assign micromat[3][57] = 9'b111111111;
assign micromat[3][58] = 9'b111111111;
assign micromat[3][59] = 9'b111111111;
assign micromat[3][60] = 9'b111111111;
assign micromat[3][61] = 9'b111111111;
assign micromat[3][62] = 9'b111111111;
assign micromat[3][63] = 9'b111111111;
assign micromat[3][64] = 9'b111111111;
assign micromat[3][65] = 9'b111111111;
assign micromat[3][66] = 9'b111111111;
assign micromat[3][67] = 9'b111111111;
assign micromat[3][68] = 9'b111111111;
assign micromat[3][69] = 9'b111111111;
assign micromat[3][70] = 9'b111111111;
assign micromat[3][71] = 9'b111111111;
assign micromat[3][72] = 9'b111111111;
assign micromat[3][73] = 9'b111111111;
assign micromat[3][74] = 9'b111111111;
assign micromat[3][75] = 9'b111111111;
assign micromat[3][76] = 9'b111111111;
assign micromat[3][77] = 9'b111111111;
assign micromat[3][78] = 9'b111111111;
assign micromat[3][79] = 9'b111111111;
assign micromat[3][80] = 9'b111111111;
assign micromat[3][81] = 9'b111111111;
assign micromat[3][82] = 9'b111111111;
assign micromat[3][83] = 9'b111111111;
assign micromat[3][84] = 9'b111111111;
assign micromat[3][85] = 9'b111111111;
assign micromat[3][86] = 9'b111111111;
assign micromat[3][87] = 9'b111111111;
assign micromat[3][88] = 9'b111111111;
assign micromat[3][89] = 9'b111111111;
assign micromat[3][90] = 9'b111111111;
assign micromat[3][91] = 9'b111111111;
assign micromat[3][92] = 9'b111111111;
assign micromat[3][93] = 9'b111111111;
assign micromat[3][94] = 9'b111111111;
assign micromat[3][95] = 9'b111111111;
assign micromat[3][96] = 9'b111111111;
assign micromat[3][97] = 9'b111111111;
assign micromat[3][98] = 9'b111111111;
assign micromat[3][99] = 9'b111111111;
assign micromat[4][0] = 9'b111111111;
assign micromat[4][1] = 9'b111111111;
assign micromat[4][2] = 9'b111111111;
assign micromat[4][3] = 9'b111111111;
assign micromat[4][4] = 9'b111111111;
assign micromat[4][5] = 9'b111111111;
assign micromat[4][6] = 9'b111111111;
assign micromat[4][7] = 9'b111111111;
assign micromat[4][8] = 9'b111111111;
assign micromat[4][9] = 9'b111111111;
assign micromat[4][10] = 9'b111111111;
assign micromat[4][11] = 9'b111111111;
assign micromat[4][12] = 9'b111111111;
assign micromat[4][13] = 9'b111111111;
assign micromat[4][14] = 9'b111111111;
assign micromat[4][15] = 9'b111111111;
assign micromat[4][16] = 9'b111111111;
assign micromat[4][17] = 9'b111111111;
assign micromat[4][18] = 9'b111111111;
assign micromat[4][19] = 9'b111111111;
assign micromat[4][20] = 9'b111111111;
assign micromat[4][21] = 9'b111111111;
assign micromat[4][22] = 9'b111111111;
assign micromat[4][23] = 9'b111111111;
assign micromat[4][24] = 9'b111111111;
assign micromat[4][25] = 9'b111111111;
assign micromat[4][26] = 9'b111111111;
assign micromat[4][27] = 9'b111111111;
assign micromat[4][28] = 9'b111111111;
assign micromat[4][29] = 9'b111111111;
assign micromat[4][30] = 9'b111111111;
assign micromat[4][31] = 9'b111111111;
assign micromat[4][32] = 9'b111111111;
assign micromat[4][33] = 9'b111111111;
assign micromat[4][34] = 9'b111111111;
assign micromat[4][35] = 9'b111111111;
assign micromat[4][36] = 9'b111111111;
assign micromat[4][37] = 9'b111111111;
assign micromat[4][38] = 9'b111111111;
assign micromat[4][39] = 9'b111111111;
assign micromat[4][40] = 9'b111111111;
assign micromat[4][41] = 9'b111111111;
assign micromat[4][42] = 9'b111111111;
assign micromat[4][43] = 9'b111111111;
assign micromat[4][44] = 9'b111111111;
assign micromat[4][45] = 9'b111111111;
assign micromat[4][46] = 9'b111111111;
assign micromat[4][47] = 9'b111111111;
assign micromat[4][48] = 9'b111111111;
assign micromat[4][49] = 9'b111111111;
assign micromat[4][50] = 9'b111111111;
assign micromat[4][51] = 9'b111111111;
assign micromat[4][52] = 9'b111111111;
assign micromat[4][53] = 9'b111111111;
assign micromat[4][54] = 9'b111111111;
assign micromat[4][55] = 9'b111111111;
assign micromat[4][56] = 9'b111111111;
assign micromat[4][57] = 9'b111111111;
assign micromat[4][58] = 9'b111111111;
assign micromat[4][59] = 9'b111111111;
assign micromat[4][60] = 9'b111111111;
assign micromat[4][61] = 9'b111111111;
assign micromat[4][62] = 9'b111111111;
assign micromat[4][63] = 9'b111111111;
assign micromat[4][64] = 9'b111111111;
assign micromat[4][65] = 9'b111111111;
assign micromat[4][66] = 9'b111111111;
assign micromat[4][67] = 9'b111111111;
assign micromat[4][68] = 9'b111111111;
assign micromat[4][69] = 9'b111111111;
assign micromat[4][70] = 9'b111111111;
assign micromat[4][71] = 9'b111111111;
assign micromat[4][72] = 9'b111111111;
assign micromat[4][73] = 9'b111111111;
assign micromat[4][74] = 9'b111111111;
assign micromat[4][75] = 9'b111111111;
assign micromat[4][76] = 9'b111111111;
assign micromat[4][77] = 9'b111111111;
assign micromat[4][78] = 9'b111111111;
assign micromat[4][79] = 9'b111111111;
assign micromat[4][80] = 9'b111111111;
assign micromat[4][81] = 9'b111111111;
assign micromat[4][82] = 9'b111111111;
assign micromat[4][83] = 9'b111111111;
assign micromat[4][84] = 9'b111111111;
assign micromat[4][85] = 9'b111111111;
assign micromat[4][86] = 9'b111111111;
assign micromat[4][87] = 9'b111111111;
assign micromat[4][88] = 9'b111111111;
assign micromat[4][89] = 9'b111111111;
assign micromat[4][90] = 9'b111111111;
assign micromat[4][91] = 9'b111111111;
assign micromat[4][92] = 9'b111111111;
assign micromat[4][93] = 9'b111111111;
assign micromat[4][94] = 9'b111111111;
assign micromat[4][95] = 9'b111111111;
assign micromat[4][96] = 9'b111111111;
assign micromat[4][97] = 9'b111111111;
assign micromat[4][98] = 9'b111111111;
assign micromat[4][99] = 9'b111111111;
assign micromat[5][0] = 9'b111111111;
assign micromat[5][1] = 9'b111111111;
assign micromat[5][2] = 9'b111111111;
assign micromat[5][3] = 9'b111111111;
assign micromat[5][4] = 9'b111111111;
assign micromat[5][5] = 9'b111111111;
assign micromat[5][6] = 9'b111111111;
assign micromat[5][7] = 9'b111111111;
assign micromat[5][8] = 9'b111111111;
assign micromat[5][9] = 9'b111111111;
assign micromat[5][10] = 9'b111111111;
assign micromat[5][11] = 9'b111111111;
assign micromat[5][12] = 9'b111111111;
assign micromat[5][13] = 9'b111111111;
assign micromat[5][14] = 9'b111111111;
assign micromat[5][15] = 9'b111111111;
assign micromat[5][16] = 9'b111111111;
assign micromat[5][17] = 9'b111111111;
assign micromat[5][18] = 9'b111111111;
assign micromat[5][19] = 9'b111111111;
assign micromat[5][20] = 9'b111111111;
assign micromat[5][21] = 9'b111111111;
assign micromat[5][22] = 9'b111111111;
assign micromat[5][23] = 9'b111111111;
assign micromat[5][24] = 9'b111111111;
assign micromat[5][25] = 9'b111111111;
assign micromat[5][26] = 9'b111111111;
assign micromat[5][27] = 9'b111111111;
assign micromat[5][28] = 9'b111111111;
assign micromat[5][29] = 9'b111111111;
assign micromat[5][30] = 9'b111111111;
assign micromat[5][31] = 9'b111111111;
assign micromat[5][32] = 9'b111111111;
assign micromat[5][33] = 9'b111111111;
assign micromat[5][34] = 9'b111111111;
assign micromat[5][35] = 9'b111111111;
assign micromat[5][36] = 9'b111111111;
assign micromat[5][37] = 9'b111111111;
assign micromat[5][38] = 9'b111111111;
assign micromat[5][39] = 9'b111111111;
assign micromat[5][40] = 9'b111111111;
assign micromat[5][41] = 9'b111111111;
assign micromat[5][42] = 9'b111111111;
assign micromat[5][43] = 9'b111111111;
assign micromat[5][44] = 9'b111111111;
assign micromat[5][45] = 9'b111111111;
assign micromat[5][46] = 9'b111111111;
assign micromat[5][47] = 9'b111111111;
assign micromat[5][48] = 9'b111111111;
assign micromat[5][49] = 9'b111111111;
assign micromat[5][50] = 9'b111111111;
assign micromat[5][51] = 9'b111111111;
assign micromat[5][52] = 9'b111111111;
assign micromat[5][53] = 9'b111111111;
assign micromat[5][54] = 9'b111111111;
assign micromat[5][55] = 9'b111111111;
assign micromat[5][56] = 9'b111111111;
assign micromat[5][57] = 9'b111111111;
assign micromat[5][58] = 9'b111111111;
assign micromat[5][59] = 9'b111111111;
assign micromat[5][60] = 9'b111111111;
assign micromat[5][61] = 9'b111111111;
assign micromat[5][62] = 9'b111111111;
assign micromat[5][63] = 9'b111111111;
assign micromat[5][64] = 9'b111111111;
assign micromat[5][65] = 9'b111111111;
assign micromat[5][66] = 9'b111111111;
assign micromat[5][67] = 9'b111111111;
assign micromat[5][68] = 9'b111111111;
assign micromat[5][69] = 9'b111111111;
assign micromat[5][70] = 9'b111111111;
assign micromat[5][71] = 9'b111111111;
assign micromat[5][72] = 9'b111111111;
assign micromat[5][73] = 9'b111111111;
assign micromat[5][74] = 9'b111111111;
assign micromat[5][75] = 9'b111111111;
assign micromat[5][76] = 9'b111111111;
assign micromat[5][77] = 9'b111111111;
assign micromat[5][78] = 9'b111111111;
assign micromat[5][79] = 9'b111111111;
assign micromat[5][80] = 9'b111111111;
assign micromat[5][81] = 9'b111111111;
assign micromat[5][82] = 9'b111111111;
assign micromat[5][83] = 9'b111111111;
assign micromat[5][84] = 9'b111111111;
assign micromat[5][85] = 9'b111111111;
assign micromat[5][86] = 9'b111111111;
assign micromat[5][87] = 9'b111111111;
assign micromat[5][88] = 9'b111111111;
assign micromat[5][89] = 9'b111111111;
assign micromat[5][90] = 9'b111111111;
assign micromat[5][91] = 9'b111111111;
assign micromat[5][92] = 9'b111111111;
assign micromat[5][93] = 9'b111111111;
assign micromat[5][94] = 9'b111111111;
assign micromat[5][95] = 9'b111111111;
assign micromat[5][96] = 9'b111111111;
assign micromat[5][97] = 9'b111111111;
assign micromat[5][98] = 9'b111111111;
assign micromat[5][99] = 9'b111111111;
assign micromat[6][0] = 9'b111111111;
assign micromat[6][1] = 9'b111111111;
assign micromat[6][2] = 9'b111111111;
assign micromat[6][3] = 9'b111111111;
assign micromat[6][4] = 9'b111111111;
assign micromat[6][5] = 9'b111111111;
assign micromat[6][6] = 9'b111111111;
assign micromat[6][7] = 9'b111111111;
assign micromat[6][8] = 9'b111111111;
assign micromat[6][9] = 9'b111111111;
assign micromat[6][10] = 9'b111111111;
assign micromat[6][11] = 9'b111111111;
assign micromat[6][12] = 9'b111111111;
assign micromat[6][13] = 9'b111111111;
assign micromat[6][14] = 9'b111111111;
assign micromat[6][15] = 9'b111111111;
assign micromat[6][16] = 9'b111111111;
assign micromat[6][17] = 9'b111111111;
assign micromat[6][18] = 9'b111111111;
assign micromat[6][19] = 9'b111111111;
assign micromat[6][20] = 9'b111111111;
assign micromat[6][21] = 9'b111111111;
assign micromat[6][22] = 9'b111111111;
assign micromat[6][23] = 9'b111111111;
assign micromat[6][24] = 9'b111111111;
assign micromat[6][25] = 9'b111111111;
assign micromat[6][26] = 9'b111111111;
assign micromat[6][27] = 9'b111111111;
assign micromat[6][28] = 9'b111111111;
assign micromat[6][29] = 9'b111111111;
assign micromat[6][30] = 9'b111111111;
assign micromat[6][31] = 9'b111111111;
assign micromat[6][32] = 9'b111111111;
assign micromat[6][33] = 9'b111111111;
assign micromat[6][34] = 9'b111111111;
assign micromat[6][35] = 9'b111111111;
assign micromat[6][36] = 9'b111111111;
assign micromat[6][37] = 9'b111111111;
assign micromat[6][38] = 9'b111111111;
assign micromat[6][39] = 9'b111111111;
assign micromat[6][40] = 9'b111111111;
assign micromat[6][41] = 9'b111111111;
assign micromat[6][42] = 9'b111111111;
assign micromat[6][43] = 9'b111111111;
assign micromat[6][44] = 9'b111111111;
assign micromat[6][45] = 9'b111111111;
assign micromat[6][46] = 9'b111111111;
assign micromat[6][47] = 9'b111111111;
assign micromat[6][48] = 9'b111111111;
assign micromat[6][49] = 9'b111111111;
assign micromat[6][50] = 9'b111111111;
assign micromat[6][51] = 9'b111111111;
assign micromat[6][52] = 9'b111111111;
assign micromat[6][53] = 9'b111111111;
assign micromat[6][54] = 9'b111111111;
assign micromat[6][55] = 9'b111111111;
assign micromat[6][56] = 9'b111111111;
assign micromat[6][57] = 9'b111111111;
assign micromat[6][58] = 9'b111111111;
assign micromat[6][59] = 9'b111111111;
assign micromat[6][60] = 9'b111111111;
assign micromat[6][61] = 9'b111111111;
assign micromat[6][62] = 9'b111111111;
assign micromat[6][63] = 9'b111111111;
assign micromat[6][64] = 9'b111111111;
assign micromat[6][65] = 9'b111111111;
assign micromat[6][66] = 9'b111111111;
assign micromat[6][67] = 9'b111111111;
assign micromat[6][68] = 9'b111111111;
assign micromat[6][69] = 9'b111111111;
assign micromat[6][70] = 9'b111111111;
assign micromat[6][71] = 9'b111111111;
assign micromat[6][72] = 9'b111111111;
assign micromat[6][73] = 9'b111111111;
assign micromat[6][74] = 9'b111111111;
assign micromat[6][75] = 9'b111111111;
assign micromat[6][76] = 9'b111111111;
assign micromat[6][77] = 9'b111111111;
assign micromat[6][78] = 9'b111111111;
assign micromat[6][79] = 9'b111111111;
assign micromat[6][80] = 9'b111111111;
assign micromat[6][81] = 9'b111111111;
assign micromat[6][82] = 9'b111111111;
assign micromat[6][83] = 9'b111111111;
assign micromat[6][84] = 9'b111111111;
assign micromat[6][85] = 9'b111111111;
assign micromat[6][86] = 9'b111111111;
assign micromat[6][87] = 9'b111111111;
assign micromat[6][88] = 9'b111111111;
assign micromat[6][89] = 9'b111111111;
assign micromat[6][90] = 9'b111111111;
assign micromat[6][91] = 9'b111111111;
assign micromat[6][92] = 9'b111111111;
assign micromat[6][93] = 9'b111111111;
assign micromat[6][94] = 9'b111111111;
assign micromat[6][95] = 9'b111111111;
assign micromat[6][96] = 9'b111111111;
assign micromat[6][97] = 9'b111111111;
assign micromat[6][98] = 9'b111111111;
assign micromat[6][99] = 9'b111111111;
assign micromat[7][0] = 9'b111111111;
assign micromat[7][1] = 9'b111111111;
assign micromat[7][2] = 9'b111111111;
assign micromat[7][3] = 9'b111111111;
assign micromat[7][4] = 9'b111111111;
assign micromat[7][5] = 9'b111111111;
assign micromat[7][6] = 9'b111111111;
assign micromat[7][7] = 9'b111111111;
assign micromat[7][8] = 9'b111111111;
assign micromat[7][9] = 9'b111111111;
assign micromat[7][10] = 9'b111111111;
assign micromat[7][11] = 9'b111111111;
assign micromat[7][12] = 9'b111111111;
assign micromat[7][13] = 9'b111111111;
assign micromat[7][14] = 9'b111111111;
assign micromat[7][15] = 9'b111111111;
assign micromat[7][16] = 9'b111111111;
assign micromat[7][17] = 9'b111111111;
assign micromat[7][18] = 9'b111111111;
assign micromat[7][19] = 9'b111111111;
assign micromat[7][20] = 9'b111111111;
assign micromat[7][21] = 9'b111111111;
assign micromat[7][22] = 9'b111111111;
assign micromat[7][23] = 9'b111111111;
assign micromat[7][24] = 9'b111111111;
assign micromat[7][25] = 9'b111111111;
assign micromat[7][26] = 9'b111111111;
assign micromat[7][27] = 9'b111111111;
assign micromat[7][28] = 9'b111111111;
assign micromat[7][29] = 9'b111111111;
assign micromat[7][30] = 9'b111111111;
assign micromat[7][31] = 9'b111111111;
assign micromat[7][32] = 9'b111111111;
assign micromat[7][33] = 9'b111111111;
assign micromat[7][34] = 9'b111111111;
assign micromat[7][35] = 9'b111111111;
assign micromat[7][36] = 9'b111111111;
assign micromat[7][37] = 9'b111111111;
assign micromat[7][38] = 9'b111111111;
assign micromat[7][39] = 9'b111111111;
assign micromat[7][40] = 9'b111111111;
assign micromat[7][41] = 9'b111111111;
assign micromat[7][42] = 9'b111111111;
assign micromat[7][43] = 9'b111111111;
assign micromat[7][44] = 9'b111111111;
assign micromat[7][45] = 9'b111111111;
assign micromat[7][46] = 9'b111111111;
assign micromat[7][47] = 9'b111111111;
assign micromat[7][48] = 9'b111111111;
assign micromat[7][49] = 9'b111111111;
assign micromat[7][50] = 9'b111111111;
assign micromat[7][51] = 9'b111111111;
assign micromat[7][52] = 9'b111111111;
assign micromat[7][53] = 9'b111111111;
assign micromat[7][54] = 9'b111111111;
assign micromat[7][55] = 9'b111111111;
assign micromat[7][56] = 9'b111111111;
assign micromat[7][57] = 9'b111111111;
assign micromat[7][58] = 9'b111111111;
assign micromat[7][59] = 9'b111111111;
assign micromat[7][60] = 9'b111111111;
assign micromat[7][61] = 9'b111111111;
assign micromat[7][62] = 9'b111111111;
assign micromat[7][63] = 9'b111111111;
assign micromat[7][64] = 9'b111111111;
assign micromat[7][65] = 9'b111111111;
assign micromat[7][66] = 9'b111111111;
assign micromat[7][67] = 9'b111111111;
assign micromat[7][68] = 9'b111111111;
assign micromat[7][69] = 9'b111111111;
assign micromat[7][70] = 9'b111111111;
assign micromat[7][71] = 9'b111111111;
assign micromat[7][72] = 9'b111111111;
assign micromat[7][73] = 9'b111111111;
assign micromat[7][74] = 9'b111111111;
assign micromat[7][75] = 9'b111111111;
assign micromat[7][76] = 9'b111111111;
assign micromat[7][77] = 9'b111111111;
assign micromat[7][78] = 9'b111111111;
assign micromat[7][79] = 9'b111111111;
assign micromat[7][80] = 9'b111111111;
assign micromat[7][81] = 9'b111111111;
assign micromat[7][82] = 9'b111111111;
assign micromat[7][83] = 9'b111111111;
assign micromat[7][84] = 9'b111111111;
assign micromat[7][85] = 9'b111111111;
assign micromat[7][86] = 9'b111111111;
assign micromat[7][87] = 9'b111111111;
assign micromat[7][88] = 9'b111111111;
assign micromat[7][89] = 9'b111111111;
assign micromat[7][90] = 9'b111111111;
assign micromat[7][91] = 9'b111111111;
assign micromat[7][92] = 9'b111111111;
assign micromat[7][93] = 9'b111111111;
assign micromat[7][94] = 9'b111111111;
assign micromat[7][95] = 9'b111111111;
assign micromat[7][96] = 9'b111111111;
assign micromat[7][97] = 9'b111111111;
assign micromat[7][98] = 9'b111111111;
assign micromat[7][99] = 9'b111111111;
assign micromat[8][0] = 9'b111111111;
assign micromat[8][1] = 9'b111111111;
assign micromat[8][2] = 9'b111111111;
assign micromat[8][3] = 9'b111111111;
assign micromat[8][4] = 9'b111111111;
assign micromat[8][5] = 9'b111111111;
assign micromat[8][6] = 9'b111111111;
assign micromat[8][7] = 9'b111111111;
assign micromat[8][8] = 9'b111111111;
assign micromat[8][9] = 9'b111111111;
assign micromat[8][10] = 9'b111111111;
assign micromat[8][11] = 9'b111111111;
assign micromat[8][12] = 9'b111111111;
assign micromat[8][13] = 9'b111111111;
assign micromat[8][14] = 9'b111111111;
assign micromat[8][15] = 9'b111111111;
assign micromat[8][16] = 9'b111111111;
assign micromat[8][17] = 9'b111111111;
assign micromat[8][18] = 9'b111111111;
assign micromat[8][19] = 9'b111111111;
assign micromat[8][20] = 9'b111111111;
assign micromat[8][21] = 9'b111111111;
assign micromat[8][22] = 9'b111111111;
assign micromat[8][23] = 9'b111111111;
assign micromat[8][24] = 9'b111111111;
assign micromat[8][25] = 9'b111111111;
assign micromat[8][26] = 9'b111111111;
assign micromat[8][27] = 9'b111111111;
assign micromat[8][28] = 9'b111111111;
assign micromat[8][29] = 9'b111111111;
assign micromat[8][30] = 9'b111111111;
assign micromat[8][31] = 9'b111111111;
assign micromat[8][32] = 9'b111111111;
assign micromat[8][33] = 9'b111111111;
assign micromat[8][34] = 9'b111111111;
assign micromat[8][35] = 9'b111111111;
assign micromat[8][36] = 9'b111111111;
assign micromat[8][37] = 9'b111111111;
assign micromat[8][38] = 9'b111111111;
assign micromat[8][39] = 9'b111111111;
assign micromat[8][40] = 9'b111111111;
assign micromat[8][41] = 9'b111111111;
assign micromat[8][42] = 9'b111111111;
assign micromat[8][43] = 9'b111111111;
assign micromat[8][44] = 9'b111111111;
assign micromat[8][45] = 9'b111111111;
assign micromat[8][46] = 9'b111111111;
assign micromat[8][47] = 9'b111111111;
assign micromat[8][48] = 9'b111111111;
assign micromat[8][49] = 9'b111111111;
assign micromat[8][50] = 9'b111111111;
assign micromat[8][51] = 9'b111111111;
assign micromat[8][52] = 9'b111111111;
assign micromat[8][53] = 9'b111111111;
assign micromat[8][54] = 9'b111111111;
assign micromat[8][55] = 9'b111111111;
assign micromat[8][56] = 9'b111111111;
assign micromat[8][57] = 9'b111111111;
assign micromat[8][58] = 9'b111111111;
assign micromat[8][59] = 9'b111111111;
assign micromat[8][60] = 9'b111111111;
assign micromat[8][61] = 9'b111111111;
assign micromat[8][62] = 9'b111111111;
assign micromat[8][63] = 9'b111111111;
assign micromat[8][64] = 9'b111111111;
assign micromat[8][65] = 9'b111111111;
assign micromat[8][66] = 9'b111111111;
assign micromat[8][67] = 9'b111111111;
assign micromat[8][68] = 9'b111111111;
assign micromat[8][69] = 9'b111111111;
assign micromat[8][70] = 9'b111111111;
assign micromat[8][71] = 9'b111111111;
assign micromat[8][72] = 9'b111111111;
assign micromat[8][73] = 9'b111111111;
assign micromat[8][74] = 9'b111111111;
assign micromat[8][75] = 9'b111111111;
assign micromat[8][76] = 9'b111111111;
assign micromat[8][77] = 9'b111111111;
assign micromat[8][78] = 9'b111111111;
assign micromat[8][79] = 9'b111111111;
assign micromat[8][80] = 9'b111111111;
assign micromat[8][81] = 9'b111111111;
assign micromat[8][82] = 9'b111111111;
assign micromat[8][83] = 9'b111111111;
assign micromat[8][84] = 9'b111111111;
assign micromat[8][85] = 9'b111111111;
assign micromat[8][86] = 9'b111111111;
assign micromat[8][87] = 9'b111111111;
assign micromat[8][88] = 9'b111111111;
assign micromat[8][89] = 9'b111111111;
assign micromat[8][90] = 9'b111111111;
assign micromat[8][91] = 9'b111111111;
assign micromat[8][92] = 9'b111111111;
assign micromat[8][93] = 9'b111111111;
assign micromat[8][94] = 9'b111111111;
assign micromat[8][95] = 9'b111111111;
assign micromat[8][96] = 9'b111111111;
assign micromat[8][97] = 9'b111111111;
assign micromat[8][98] = 9'b111111111;
assign micromat[8][99] = 9'b111111111;
assign micromat[9][0] = 9'b111111111;
assign micromat[9][1] = 9'b111111111;
assign micromat[9][2] = 9'b111111111;
assign micromat[9][3] = 9'b111111111;
assign micromat[9][4] = 9'b111111111;
assign micromat[9][5] = 9'b111111111;
assign micromat[9][6] = 9'b111111111;
assign micromat[9][7] = 9'b111111111;
assign micromat[9][8] = 9'b111111111;
assign micromat[9][9] = 9'b111111111;
assign micromat[9][10] = 9'b111111111;
assign micromat[9][11] = 9'b111111111;
assign micromat[9][12] = 9'b111111111;
assign micromat[9][13] = 9'b111111111;
assign micromat[9][14] = 9'b111111111;
assign micromat[9][15] = 9'b111111111;
assign micromat[9][16] = 9'b111111111;
assign micromat[9][17] = 9'b111111111;
assign micromat[9][18] = 9'b111111111;
assign micromat[9][19] = 9'b111111111;
assign micromat[9][20] = 9'b111111111;
assign micromat[9][21] = 9'b111111111;
assign micromat[9][22] = 9'b111111111;
assign micromat[9][23] = 9'b111111111;
assign micromat[9][24] = 9'b111111111;
assign micromat[9][25] = 9'b111111111;
assign micromat[9][26] = 9'b111111111;
assign micromat[9][27] = 9'b111111111;
assign micromat[9][28] = 9'b111111111;
assign micromat[9][29] = 9'b111111111;
assign micromat[9][30] = 9'b111111111;
assign micromat[9][31] = 9'b111111111;
assign micromat[9][32] = 9'b111111111;
assign micromat[9][33] = 9'b111111111;
assign micromat[9][34] = 9'b111111111;
assign micromat[9][35] = 9'b111111111;
assign micromat[9][36] = 9'b111111111;
assign micromat[9][37] = 9'b111111111;
assign micromat[9][38] = 9'b111111111;
assign micromat[9][39] = 9'b111111111;
assign micromat[9][40] = 9'b111111111;
assign micromat[9][41] = 9'b111111111;
assign micromat[9][42] = 9'b111111111;
assign micromat[9][43] = 9'b111111111;
assign micromat[9][44] = 9'b111111111;
assign micromat[9][45] = 9'b111111111;
assign micromat[9][46] = 9'b111111111;
assign micromat[9][47] = 9'b111111111;
assign micromat[9][48] = 9'b111111111;
assign micromat[9][49] = 9'b111111111;
assign micromat[9][50] = 9'b111111111;
assign micromat[9][51] = 9'b111111111;
assign micromat[9][52] = 9'b111111111;
assign micromat[9][53] = 9'b111111111;
assign micromat[9][54] = 9'b111111111;
assign micromat[9][55] = 9'b111111111;
assign micromat[9][56] = 9'b111111111;
assign micromat[9][57] = 9'b111111111;
assign micromat[9][58] = 9'b111111111;
assign micromat[9][59] = 9'b111111111;
assign micromat[9][60] = 9'b111111111;
assign micromat[9][61] = 9'b111111111;
assign micromat[9][62] = 9'b111111111;
assign micromat[9][63] = 9'b111111111;
assign micromat[9][64] = 9'b111111111;
assign micromat[9][65] = 9'b111111111;
assign micromat[9][66] = 9'b111111111;
assign micromat[9][67] = 9'b111111111;
assign micromat[9][68] = 9'b111111111;
assign micromat[9][69] = 9'b111111111;
assign micromat[9][70] = 9'b111111111;
assign micromat[9][71] = 9'b111111111;
assign micromat[9][72] = 9'b111111111;
assign micromat[9][73] = 9'b111111111;
assign micromat[9][74] = 9'b111111111;
assign micromat[9][75] = 9'b111111111;
assign micromat[9][76] = 9'b111111111;
assign micromat[9][77] = 9'b111111111;
assign micromat[9][78] = 9'b111111111;
assign micromat[9][79] = 9'b111111111;
assign micromat[9][80] = 9'b111111111;
assign micromat[9][81] = 9'b111111111;
assign micromat[9][82] = 9'b111111111;
assign micromat[9][83] = 9'b111111111;
assign micromat[9][84] = 9'b111111111;
assign micromat[9][85] = 9'b111111111;
assign micromat[9][86] = 9'b111111111;
assign micromat[9][87] = 9'b111111111;
assign micromat[9][88] = 9'b111111111;
assign micromat[9][89] = 9'b111111111;
assign micromat[9][90] = 9'b111111111;
assign micromat[9][91] = 9'b111111111;
assign micromat[9][92] = 9'b111111111;
assign micromat[9][93] = 9'b111111111;
assign micromat[9][94] = 9'b111111111;
assign micromat[9][95] = 9'b111111111;
assign micromat[9][96] = 9'b111111111;
assign micromat[9][97] = 9'b111111111;
assign micromat[9][98] = 9'b111111111;
assign micromat[9][99] = 9'b111111111;
assign micromat[10][0] = 9'b111111111;
assign micromat[10][1] = 9'b111111111;
assign micromat[10][2] = 9'b111111111;
assign micromat[10][3] = 9'b111111111;
assign micromat[10][4] = 9'b111111111;
assign micromat[10][5] = 9'b111111111;
assign micromat[10][6] = 9'b111111111;
assign micromat[10][7] = 9'b111111111;
assign micromat[10][8] = 9'b111111111;
assign micromat[10][9] = 9'b111111111;
assign micromat[10][10] = 9'b111111111;
assign micromat[10][11] = 9'b111111111;
assign micromat[10][12] = 9'b111111111;
assign micromat[10][13] = 9'b111111111;
assign micromat[10][14] = 9'b111111111;
assign micromat[10][15] = 9'b111111111;
assign micromat[10][16] = 9'b111111111;
assign micromat[10][17] = 9'b111111111;
assign micromat[10][18] = 9'b111111111;
assign micromat[10][19] = 9'b111111111;
assign micromat[10][20] = 9'b111111111;
assign micromat[10][21] = 9'b111111111;
assign micromat[10][22] = 9'b111111111;
assign micromat[10][23] = 9'b111111111;
assign micromat[10][24] = 9'b111111111;
assign micromat[10][25] = 9'b111111111;
assign micromat[10][26] = 9'b111111111;
assign micromat[10][27] = 9'b111111111;
assign micromat[10][28] = 9'b111111111;
assign micromat[10][29] = 9'b111111111;
assign micromat[10][30] = 9'b111111111;
assign micromat[10][31] = 9'b111111111;
assign micromat[10][32] = 9'b111111111;
assign micromat[10][33] = 9'b111111111;
assign micromat[10][34] = 9'b111111111;
assign micromat[10][35] = 9'b111111111;
assign micromat[10][36] = 9'b111111111;
assign micromat[10][37] = 9'b111111111;
assign micromat[10][38] = 9'b111111111;
assign micromat[10][39] = 9'b111111111;
assign micromat[10][40] = 9'b111111111;
assign micromat[10][41] = 9'b111111111;
assign micromat[10][42] = 9'b111111111;
assign micromat[10][43] = 9'b111111111;
assign micromat[10][44] = 9'b111111111;
assign micromat[10][45] = 9'b111111111;
assign micromat[10][46] = 9'b111111111;
assign micromat[10][47] = 9'b111111111;
assign micromat[10][48] = 9'b111111111;
assign micromat[10][49] = 9'b111111111;
assign micromat[10][50] = 9'b111111111;
assign micromat[10][51] = 9'b111111111;
assign micromat[10][52] = 9'b111111111;
assign micromat[10][53] = 9'b111111111;
assign micromat[10][54] = 9'b111111111;
assign micromat[10][55] = 9'b111111111;
assign micromat[10][56] = 9'b111111111;
assign micromat[10][57] = 9'b111111111;
assign micromat[10][58] = 9'b111111111;
assign micromat[10][59] = 9'b111111111;
assign micromat[10][60] = 9'b111111111;
assign micromat[10][61] = 9'b111111111;
assign micromat[10][62] = 9'b111111111;
assign micromat[10][63] = 9'b111111111;
assign micromat[10][64] = 9'b111111111;
assign micromat[10][65] = 9'b111111111;
assign micromat[10][66] = 9'b111111111;
assign micromat[10][67] = 9'b111111111;
assign micromat[10][68] = 9'b111111111;
assign micromat[10][69] = 9'b111111111;
assign micromat[10][70] = 9'b111111111;
assign micromat[10][71] = 9'b111111111;
assign micromat[10][72] = 9'b111111111;
assign micromat[10][73] = 9'b111111111;
assign micromat[10][74] = 9'b111111111;
assign micromat[10][75] = 9'b111111111;
assign micromat[10][76] = 9'b111111111;
assign micromat[10][77] = 9'b111111111;
assign micromat[10][78] = 9'b111111111;
assign micromat[10][79] = 9'b111111111;
assign micromat[10][80] = 9'b111111111;
assign micromat[10][81] = 9'b111111111;
assign micromat[10][82] = 9'b111111111;
assign micromat[10][83] = 9'b111111111;
assign micromat[10][84] = 9'b111111111;
assign micromat[10][85] = 9'b111111111;
assign micromat[10][86] = 9'b111111111;
assign micromat[10][87] = 9'b111111111;
assign micromat[10][88] = 9'b111111111;
assign micromat[10][89] = 9'b111111111;
assign micromat[10][90] = 9'b111111111;
assign micromat[10][91] = 9'b111111111;
assign micromat[10][92] = 9'b111111111;
assign micromat[10][93] = 9'b111111111;
assign micromat[10][94] = 9'b111111111;
assign micromat[10][95] = 9'b111111111;
assign micromat[10][96] = 9'b111111111;
assign micromat[10][97] = 9'b111111111;
assign micromat[10][98] = 9'b111111111;
assign micromat[10][99] = 9'b111111111;
assign micromat[11][0] = 9'b111111111;
assign micromat[11][1] = 9'b111111111;
assign micromat[11][2] = 9'b111111111;
assign micromat[11][3] = 9'b111111111;
assign micromat[11][4] = 9'b111111111;
assign micromat[11][5] = 9'b111111111;
assign micromat[11][6] = 9'b111111111;
assign micromat[11][7] = 9'b111111111;
assign micromat[11][8] = 9'b111111111;
assign micromat[11][9] = 9'b111111111;
assign micromat[11][10] = 9'b111111111;
assign micromat[11][11] = 9'b111111111;
assign micromat[11][12] = 9'b111111111;
assign micromat[11][13] = 9'b111111111;
assign micromat[11][14] = 9'b111111111;
assign micromat[11][15] = 9'b111111111;
assign micromat[11][16] = 9'b111111111;
assign micromat[11][17] = 9'b111111111;
assign micromat[11][18] = 9'b111111111;
assign micromat[11][19] = 9'b111111111;
assign micromat[11][20] = 9'b111111111;
assign micromat[11][21] = 9'b111111111;
assign micromat[11][22] = 9'b111111111;
assign micromat[11][23] = 9'b111111111;
assign micromat[11][24] = 9'b111111111;
assign micromat[11][25] = 9'b111111111;
assign micromat[11][26] = 9'b111111111;
assign micromat[11][27] = 9'b111111111;
assign micromat[11][28] = 9'b111111111;
assign micromat[11][29] = 9'b111111111;
assign micromat[11][30] = 9'b111111111;
assign micromat[11][31] = 9'b111111111;
assign micromat[11][32] = 9'b111111111;
assign micromat[11][33] = 9'b111111111;
assign micromat[11][34] = 9'b111111111;
assign micromat[11][35] = 9'b111111111;
assign micromat[11][36] = 9'b111111111;
assign micromat[11][37] = 9'b111111111;
assign micromat[11][38] = 9'b111111111;
assign micromat[11][39] = 9'b111111111;
assign micromat[11][40] = 9'b111111111;
assign micromat[11][41] = 9'b111111111;
assign micromat[11][42] = 9'b111111111;
assign micromat[11][43] = 9'b111111111;
assign micromat[11][44] = 9'b111111111;
assign micromat[11][45] = 9'b111111111;
assign micromat[11][46] = 9'b111111111;
assign micromat[11][47] = 9'b111111111;
assign micromat[11][48] = 9'b111111111;
assign micromat[11][49] = 9'b111111111;
assign micromat[11][50] = 9'b111111111;
assign micromat[11][51] = 9'b111111111;
assign micromat[11][52] = 9'b111111111;
assign micromat[11][53] = 9'b111111111;
assign micromat[11][54] = 9'b111111111;
assign micromat[11][55] = 9'b111111111;
assign micromat[11][56] = 9'b111111111;
assign micromat[11][57] = 9'b111111111;
assign micromat[11][58] = 9'b111111111;
assign micromat[11][59] = 9'b111111111;
assign micromat[11][60] = 9'b111111111;
assign micromat[11][61] = 9'b111111111;
assign micromat[11][62] = 9'b111111111;
assign micromat[11][63] = 9'b111111111;
assign micromat[11][64] = 9'b111111111;
assign micromat[11][65] = 9'b111111111;
assign micromat[11][66] = 9'b111111111;
assign micromat[11][67] = 9'b111111111;
assign micromat[11][68] = 9'b111111111;
assign micromat[11][69] = 9'b111111111;
assign micromat[11][70] = 9'b111111111;
assign micromat[11][71] = 9'b111111111;
assign micromat[11][72] = 9'b111111111;
assign micromat[11][73] = 9'b111111111;
assign micromat[11][74] = 9'b111111111;
assign micromat[11][75] = 9'b111111111;
assign micromat[11][76] = 9'b111111111;
assign micromat[11][77] = 9'b111111111;
assign micromat[11][78] = 9'b111111111;
assign micromat[11][79] = 9'b111111111;
assign micromat[11][80] = 9'b111111111;
assign micromat[11][81] = 9'b111111111;
assign micromat[11][82] = 9'b111111111;
assign micromat[11][83] = 9'b111111111;
assign micromat[11][84] = 9'b111111111;
assign micromat[11][85] = 9'b111111111;
assign micromat[11][86] = 9'b111111111;
assign micromat[11][87] = 9'b111111111;
assign micromat[11][88] = 9'b111111111;
assign micromat[11][89] = 9'b111111111;
assign micromat[11][90] = 9'b111111111;
assign micromat[11][91] = 9'b111111111;
assign micromat[11][92] = 9'b111111111;
assign micromat[11][93] = 9'b111111111;
assign micromat[11][94] = 9'b111111111;
assign micromat[11][95] = 9'b111111111;
assign micromat[11][96] = 9'b111111111;
assign micromat[11][97] = 9'b111111111;
assign micromat[11][98] = 9'b111111111;
assign micromat[11][99] = 9'b111111111;
assign micromat[12][0] = 9'b111111111;
assign micromat[12][1] = 9'b111111111;
assign micromat[12][2] = 9'b111111111;
assign micromat[12][3] = 9'b111111111;
assign micromat[12][4] = 9'b111111111;
assign micromat[12][5] = 9'b111111111;
assign micromat[12][6] = 9'b111111111;
assign micromat[12][7] = 9'b111111111;
assign micromat[12][8] = 9'b111111111;
assign micromat[12][9] = 9'b111111111;
assign micromat[12][10] = 9'b111111111;
assign micromat[12][11] = 9'b111111111;
assign micromat[12][12] = 9'b111111111;
assign micromat[12][13] = 9'b111111111;
assign micromat[12][14] = 9'b111111111;
assign micromat[12][15] = 9'b111111111;
assign micromat[12][16] = 9'b111111111;
assign micromat[12][17] = 9'b111111111;
assign micromat[12][18] = 9'b111111111;
assign micromat[12][19] = 9'b111111111;
assign micromat[12][20] = 9'b111111111;
assign micromat[12][21] = 9'b111111111;
assign micromat[12][22] = 9'b111111111;
assign micromat[12][23] = 9'b111111111;
assign micromat[12][24] = 9'b111111111;
assign micromat[12][25] = 9'b111111111;
assign micromat[12][26] = 9'b111111111;
assign micromat[12][27] = 9'b111111111;
assign micromat[12][28] = 9'b111111111;
assign micromat[12][29] = 9'b111111111;
assign micromat[12][30] = 9'b111111111;
assign micromat[12][31] = 9'b111111111;
assign micromat[12][32] = 9'b111111111;
assign micromat[12][33] = 9'b111111111;
assign micromat[12][34] = 9'b111111111;
assign micromat[12][35] = 9'b111111111;
assign micromat[12][36] = 9'b111111111;
assign micromat[12][37] = 9'b111111111;
assign micromat[12][38] = 9'b111111111;
assign micromat[12][39] = 9'b111111111;
assign micromat[12][40] = 9'b111111111;
assign micromat[12][41] = 9'b111111111;
assign micromat[12][42] = 9'b111111111;
assign micromat[12][43] = 9'b111111111;
assign micromat[12][44] = 9'b111111111;
assign micromat[12][45] = 9'b111111111;
assign micromat[12][46] = 9'b111111111;
assign micromat[12][47] = 9'b111111111;
assign micromat[12][48] = 9'b111111111;
assign micromat[12][49] = 9'b111111111;
assign micromat[12][50] = 9'b111111111;
assign micromat[12][51] = 9'b111111111;
assign micromat[12][52] = 9'b111111111;
assign micromat[12][53] = 9'b111111111;
assign micromat[12][54] = 9'b111111111;
assign micromat[12][55] = 9'b111111111;
assign micromat[12][56] = 9'b111111111;
assign micromat[12][57] = 9'b111111111;
assign micromat[12][58] = 9'b111111111;
assign micromat[12][59] = 9'b111111111;
assign micromat[12][60] = 9'b111111111;
assign micromat[12][61] = 9'b111111111;
assign micromat[12][62] = 9'b111111111;
assign micromat[12][63] = 9'b111111111;
assign micromat[12][64] = 9'b111111111;
assign micromat[12][65] = 9'b111111111;
assign micromat[12][66] = 9'b111111111;
assign micromat[12][67] = 9'b111111111;
assign micromat[12][68] = 9'b111111111;
assign micromat[12][69] = 9'b111111111;
assign micromat[12][70] = 9'b111111111;
assign micromat[12][71] = 9'b111111111;
assign micromat[12][72] = 9'b111111111;
assign micromat[12][73] = 9'b111111111;
assign micromat[12][74] = 9'b111111111;
assign micromat[12][75] = 9'b111111111;
assign micromat[12][76] = 9'b111111111;
assign micromat[12][77] = 9'b111111111;
assign micromat[12][78] = 9'b111111111;
assign micromat[12][79] = 9'b111111111;
assign micromat[12][80] = 9'b111111111;
assign micromat[12][81] = 9'b111111111;
assign micromat[12][82] = 9'b111111111;
assign micromat[12][83] = 9'b111111111;
assign micromat[12][84] = 9'b111111111;
assign micromat[12][85] = 9'b111111111;
assign micromat[12][86] = 9'b111111111;
assign micromat[12][87] = 9'b111111111;
assign micromat[12][88] = 9'b111111111;
assign micromat[12][89] = 9'b111111111;
assign micromat[12][90] = 9'b111111111;
assign micromat[12][91] = 9'b111111111;
assign micromat[12][92] = 9'b111111111;
assign micromat[12][93] = 9'b111111111;
assign micromat[12][94] = 9'b111111111;
assign micromat[12][95] = 9'b111111111;
assign micromat[12][96] = 9'b111111111;
assign micromat[12][97] = 9'b111111111;
assign micromat[12][98] = 9'b111111111;
assign micromat[12][99] = 9'b111111111;
assign micromat[13][0] = 9'b111111111;
assign micromat[13][1] = 9'b111111111;
assign micromat[13][2] = 9'b111111111;
assign micromat[13][3] = 9'b111111111;
assign micromat[13][4] = 9'b111111111;
assign micromat[13][5] = 9'b111111111;
assign micromat[13][6] = 9'b111111111;
assign micromat[13][7] = 9'b111111111;
assign micromat[13][8] = 9'b111111111;
assign micromat[13][9] = 9'b111111111;
assign micromat[13][10] = 9'b111111111;
assign micromat[13][11] = 9'b111111111;
assign micromat[13][12] = 9'b111111111;
assign micromat[13][13] = 9'b111111111;
assign micromat[13][14] = 9'b111111111;
assign micromat[13][15] = 9'b111111111;
assign micromat[13][16] = 9'b111111111;
assign micromat[13][17] = 9'b111111111;
assign micromat[13][18] = 9'b111111111;
assign micromat[13][19] = 9'b111111111;
assign micromat[13][20] = 9'b111111111;
assign micromat[13][21] = 9'b111111111;
assign micromat[13][22] = 9'b111111111;
assign micromat[13][23] = 9'b111111111;
assign micromat[13][24] = 9'b111111111;
assign micromat[13][25] = 9'b111111111;
assign micromat[13][26] = 9'b111111111;
assign micromat[13][27] = 9'b111111111;
assign micromat[13][28] = 9'b111111111;
assign micromat[13][29] = 9'b111111111;
assign micromat[13][30] = 9'b111111111;
assign micromat[13][31] = 9'b111111111;
assign micromat[13][32] = 9'b111111111;
assign micromat[13][33] = 9'b111111111;
assign micromat[13][34] = 9'b111111111;
assign micromat[13][35] = 9'b111111111;
assign micromat[13][36] = 9'b111111111;
assign micromat[13][37] = 9'b111111111;
assign micromat[13][38] = 9'b111111111;
assign micromat[13][39] = 9'b111111111;
assign micromat[13][40] = 9'b111111111;
assign micromat[13][41] = 9'b111111111;
assign micromat[13][42] = 9'b111111111;
assign micromat[13][43] = 9'b111111111;
assign micromat[13][44] = 9'b111111111;
assign micromat[13][45] = 9'b111111111;
assign micromat[13][46] = 9'b111111111;
assign micromat[13][47] = 9'b111111111;
assign micromat[13][48] = 9'b111111111;
assign micromat[13][49] = 9'b111111111;
assign micromat[13][50] = 9'b111111111;
assign micromat[13][51] = 9'b111111111;
assign micromat[13][52] = 9'b111111111;
assign micromat[13][53] = 9'b111111111;
assign micromat[13][54] = 9'b111111111;
assign micromat[13][55] = 9'b111111111;
assign micromat[13][56] = 9'b111111111;
assign micromat[13][57] = 9'b111111111;
assign micromat[13][58] = 9'b111111111;
assign micromat[13][59] = 9'b111111111;
assign micromat[13][60] = 9'b111111111;
assign micromat[13][61] = 9'b111111111;
assign micromat[13][62] = 9'b111111111;
assign micromat[13][63] = 9'b111111111;
assign micromat[13][64] = 9'b111111111;
assign micromat[13][65] = 9'b111111111;
assign micromat[13][66] = 9'b111111111;
assign micromat[13][67] = 9'b111111111;
assign micromat[13][68] = 9'b111111111;
assign micromat[13][69] = 9'b111111111;
assign micromat[13][70] = 9'b111111111;
assign micromat[13][71] = 9'b111111111;
assign micromat[13][72] = 9'b111111111;
assign micromat[13][73] = 9'b111111111;
assign micromat[13][74] = 9'b111111111;
assign micromat[13][75] = 9'b111111111;
assign micromat[13][76] = 9'b111111111;
assign micromat[13][77] = 9'b111111111;
assign micromat[13][78] = 9'b111111111;
assign micromat[13][79] = 9'b111111111;
assign micromat[13][80] = 9'b111111111;
assign micromat[13][81] = 9'b111111111;
assign micromat[13][82] = 9'b111111111;
assign micromat[13][83] = 9'b111111111;
assign micromat[13][84] = 9'b111111111;
assign micromat[13][85] = 9'b111111111;
assign micromat[13][86] = 9'b111111111;
assign micromat[13][87] = 9'b111111111;
assign micromat[13][88] = 9'b111111111;
assign micromat[13][89] = 9'b111111111;
assign micromat[13][90] = 9'b111111111;
assign micromat[13][91] = 9'b111111111;
assign micromat[13][92] = 9'b111111111;
assign micromat[13][93] = 9'b111111111;
assign micromat[13][94] = 9'b111111111;
assign micromat[13][95] = 9'b111111111;
assign micromat[13][96] = 9'b111111111;
assign micromat[13][97] = 9'b111111111;
assign micromat[13][98] = 9'b111111111;
assign micromat[13][99] = 9'b111111111;
assign micromat[14][0] = 9'b111111111;
assign micromat[14][1] = 9'b111111111;
assign micromat[14][2] = 9'b111111111;
assign micromat[14][3] = 9'b111111111;
assign micromat[14][4] = 9'b111111111;
assign micromat[14][5] = 9'b111111111;
assign micromat[14][6] = 9'b111111111;
assign micromat[14][7] = 9'b111111111;
assign micromat[14][8] = 9'b111111111;
assign micromat[14][9] = 9'b111111111;
assign micromat[14][10] = 9'b111111111;
assign micromat[14][11] = 9'b111111111;
assign micromat[14][12] = 9'b111111111;
assign micromat[14][13] = 9'b111111111;
assign micromat[14][14] = 9'b111111111;
assign micromat[14][15] = 9'b111111111;
assign micromat[14][16] = 9'b111111111;
assign micromat[14][17] = 9'b111111111;
assign micromat[14][18] = 9'b111111111;
assign micromat[14][19] = 9'b111111111;
assign micromat[14][20] = 9'b111111111;
assign micromat[14][21] = 9'b111111111;
assign micromat[14][22] = 9'b111111111;
assign micromat[14][23] = 9'b111111111;
assign micromat[14][24] = 9'b111111111;
assign micromat[14][25] = 9'b111111111;
assign micromat[14][26] = 9'b111111111;
assign micromat[14][27] = 9'b111111111;
assign micromat[14][28] = 9'b111111111;
assign micromat[14][29] = 9'b111111111;
assign micromat[14][30] = 9'b111111111;
assign micromat[14][31] = 9'b111111111;
assign micromat[14][32] = 9'b111111111;
assign micromat[14][33] = 9'b111111111;
assign micromat[14][34] = 9'b111111111;
assign micromat[14][35] = 9'b111111111;
assign micromat[14][36] = 9'b111111111;
assign micromat[14][37] = 9'b111111111;
assign micromat[14][38] = 9'b111111111;
assign micromat[14][39] = 9'b111111111;
assign micromat[14][40] = 9'b111111111;
assign micromat[14][41] = 9'b111111111;
assign micromat[14][42] = 9'b111111111;
assign micromat[14][43] = 9'b111111111;
assign micromat[14][44] = 9'b111111111;
assign micromat[14][45] = 9'b111111111;
assign micromat[14][46] = 9'b111111111;
assign micromat[14][47] = 9'b111111111;
assign micromat[14][48] = 9'b111111111;
assign micromat[14][49] = 9'b111111111;
assign micromat[14][50] = 9'b111111111;
assign micromat[14][51] = 9'b111111111;
assign micromat[14][52] = 9'b111111111;
assign micromat[14][53] = 9'b111111111;
assign micromat[14][54] = 9'b111111111;
assign micromat[14][55] = 9'b111111111;
assign micromat[14][56] = 9'b111111111;
assign micromat[14][57] = 9'b111111111;
assign micromat[14][58] = 9'b111111111;
assign micromat[14][59] = 9'b111111111;
assign micromat[14][60] = 9'b111111111;
assign micromat[14][61] = 9'b111111111;
assign micromat[14][62] = 9'b111111111;
assign micromat[14][63] = 9'b111111111;
assign micromat[14][64] = 9'b111111111;
assign micromat[14][65] = 9'b111111111;
assign micromat[14][66] = 9'b111111111;
assign micromat[14][67] = 9'b111111111;
assign micromat[14][68] = 9'b111111111;
assign micromat[14][69] = 9'b111111111;
assign micromat[14][70] = 9'b111111111;
assign micromat[14][71] = 9'b111111111;
assign micromat[14][72] = 9'b111111111;
assign micromat[14][73] = 9'b111111111;
assign micromat[14][74] = 9'b111111111;
assign micromat[14][75] = 9'b111111111;
assign micromat[14][76] = 9'b111111111;
assign micromat[14][77] = 9'b111111111;
assign micromat[14][78] = 9'b111111111;
assign micromat[14][79] = 9'b111111111;
assign micromat[14][80] = 9'b111111111;
assign micromat[14][81] = 9'b111111111;
assign micromat[14][82] = 9'b111111111;
assign micromat[14][83] = 9'b111111111;
assign micromat[14][84] = 9'b111111111;
assign micromat[14][85] = 9'b111111111;
assign micromat[14][86] = 9'b111111111;
assign micromat[14][87] = 9'b111111111;
assign micromat[14][88] = 9'b111111111;
assign micromat[14][89] = 9'b111111111;
assign micromat[14][90] = 9'b111111111;
assign micromat[14][91] = 9'b111111111;
assign micromat[14][92] = 9'b111111111;
assign micromat[14][93] = 9'b111111111;
assign micromat[14][94] = 9'b111111111;
assign micromat[14][95] = 9'b111111111;
assign micromat[14][96] = 9'b111111111;
assign micromat[14][97] = 9'b111111111;
assign micromat[14][98] = 9'b111111111;
assign micromat[14][99] = 9'b111111111;
assign micromat[15][0] = 9'b111111111;
assign micromat[15][1] = 9'b111111111;
assign micromat[15][2] = 9'b111111111;
assign micromat[15][3] = 9'b111111111;
assign micromat[15][4] = 9'b111111111;
assign micromat[15][5] = 9'b111111111;
assign micromat[15][6] = 9'b111111111;
assign micromat[15][7] = 9'b111111111;
assign micromat[15][8] = 9'b111111111;
assign micromat[15][9] = 9'b111111111;
assign micromat[15][10] = 9'b111111111;
assign micromat[15][11] = 9'b111111111;
assign micromat[15][12] = 9'b111111111;
assign micromat[15][13] = 9'b111111111;
assign micromat[15][14] = 9'b111111111;
assign micromat[15][15] = 9'b111111111;
assign micromat[15][16] = 9'b111111111;
assign micromat[15][17] = 9'b111111111;
assign micromat[15][18] = 9'b111111111;
assign micromat[15][19] = 9'b111111111;
assign micromat[15][20] = 9'b111111111;
assign micromat[15][21] = 9'b111111111;
assign micromat[15][22] = 9'b111111111;
assign micromat[15][23] = 9'b111111111;
assign micromat[15][24] = 9'b111111111;
assign micromat[15][25] = 9'b111111111;
assign micromat[15][26] = 9'b111111111;
assign micromat[15][27] = 9'b111111111;
assign micromat[15][28] = 9'b111111111;
assign micromat[15][29] = 9'b111111111;
assign micromat[15][30] = 9'b111111111;
assign micromat[15][31] = 9'b111111111;
assign micromat[15][32] = 9'b111111111;
assign micromat[15][33] = 9'b111111111;
assign micromat[15][34] = 9'b111111111;
assign micromat[15][35] = 9'b111111111;
assign micromat[15][36] = 9'b111111111;
assign micromat[15][37] = 9'b111111111;
assign micromat[15][38] = 9'b111111111;
assign micromat[15][39] = 9'b111111111;
assign micromat[15][40] = 9'b111111111;
assign micromat[15][41] = 9'b111111111;
assign micromat[15][42] = 9'b111111111;
assign micromat[15][43] = 9'b111111111;
assign micromat[15][44] = 9'b111111111;
assign micromat[15][45] = 9'b111111111;
assign micromat[15][46] = 9'b111111111;
assign micromat[15][47] = 9'b111111111;
assign micromat[15][48] = 9'b111111111;
assign micromat[15][49] = 9'b111111111;
assign micromat[15][50] = 9'b111111111;
assign micromat[15][51] = 9'b111111111;
assign micromat[15][52] = 9'b111111111;
assign micromat[15][53] = 9'b111111111;
assign micromat[15][54] = 9'b111111111;
assign micromat[15][55] = 9'b111111111;
assign micromat[15][56] = 9'b111111111;
assign micromat[15][57] = 9'b111111111;
assign micromat[15][58] = 9'b111111111;
assign micromat[15][59] = 9'b111111111;
assign micromat[15][60] = 9'b111111111;
assign micromat[15][61] = 9'b111111111;
assign micromat[15][62] = 9'b111111111;
assign micromat[15][63] = 9'b111111111;
assign micromat[15][64] = 9'b111111111;
assign micromat[15][65] = 9'b111111111;
assign micromat[15][66] = 9'b111111111;
assign micromat[15][67] = 9'b111111111;
assign micromat[15][68] = 9'b111111111;
assign micromat[15][69] = 9'b111111111;
assign micromat[15][70] = 9'b111111111;
assign micromat[15][71] = 9'b111111111;
assign micromat[15][72] = 9'b111111111;
assign micromat[15][73] = 9'b111111111;
assign micromat[15][74] = 9'b111111111;
assign micromat[15][75] = 9'b111111111;
assign micromat[15][76] = 9'b111111111;
assign micromat[15][77] = 9'b111111111;
assign micromat[15][78] = 9'b111111111;
assign micromat[15][79] = 9'b111111111;
assign micromat[15][80] = 9'b111111111;
assign micromat[15][81] = 9'b111111111;
assign micromat[15][82] = 9'b111111111;
assign micromat[15][83] = 9'b111111111;
assign micromat[15][84] = 9'b111111111;
assign micromat[15][85] = 9'b111111111;
assign micromat[15][86] = 9'b111111111;
assign micromat[15][87] = 9'b111111111;
assign micromat[15][88] = 9'b111111111;
assign micromat[15][89] = 9'b111111111;
assign micromat[15][90] = 9'b111111111;
assign micromat[15][91] = 9'b111111111;
assign micromat[15][92] = 9'b111111111;
assign micromat[15][93] = 9'b111111111;
assign micromat[15][94] = 9'b111111111;
assign micromat[15][95] = 9'b111111111;
assign micromat[15][96] = 9'b111111111;
assign micromat[15][97] = 9'b111111111;
assign micromat[15][98] = 9'b111111111;
assign micromat[15][99] = 9'b111111111;
assign micromat[16][0] = 9'b111111111;
assign micromat[16][1] = 9'b111111111;
assign micromat[16][2] = 9'b111111111;
assign micromat[16][3] = 9'b111111111;
assign micromat[16][4] = 9'b111111111;
assign micromat[16][5] = 9'b111111111;
assign micromat[16][6] = 9'b111111111;
assign micromat[16][7] = 9'b111111111;
assign micromat[16][8] = 9'b111111111;
assign micromat[16][9] = 9'b111111111;
assign micromat[16][10] = 9'b111111111;
assign micromat[16][11] = 9'b111111111;
assign micromat[16][12] = 9'b111111111;
assign micromat[16][13] = 9'b111111111;
assign micromat[16][14] = 9'b111111111;
assign micromat[16][15] = 9'b111111111;
assign micromat[16][16] = 9'b111111111;
assign micromat[16][17] = 9'b111111111;
assign micromat[16][18] = 9'b111111111;
assign micromat[16][19] = 9'b111111111;
assign micromat[16][20] = 9'b111111111;
assign micromat[16][21] = 9'b111111111;
assign micromat[16][22] = 9'b111111111;
assign micromat[16][23] = 9'b111111111;
assign micromat[16][24] = 9'b111111111;
assign micromat[16][25] = 9'b111111111;
assign micromat[16][26] = 9'b111111111;
assign micromat[16][27] = 9'b111111111;
assign micromat[16][28] = 9'b111111111;
assign micromat[16][29] = 9'b111111111;
assign micromat[16][30] = 9'b111111111;
assign micromat[16][31] = 9'b111111111;
assign micromat[16][32] = 9'b111111111;
assign micromat[16][33] = 9'b111111111;
assign micromat[16][34] = 9'b111111111;
assign micromat[16][35] = 9'b111111111;
assign micromat[16][36] = 9'b111111111;
assign micromat[16][37] = 9'b111111111;
assign micromat[16][38] = 9'b111111111;
assign micromat[16][39] = 9'b111111111;
assign micromat[16][40] = 9'b111111111;
assign micromat[16][41] = 9'b111111111;
assign micromat[16][42] = 9'b111111111;
assign micromat[16][43] = 9'b111111111;
assign micromat[16][44] = 9'b111111111;
assign micromat[16][45] = 9'b111111111;
assign micromat[16][46] = 9'b111111111;
assign micromat[16][47] = 9'b111111111;
assign micromat[16][48] = 9'b111111111;
assign micromat[16][49] = 9'b111111111;
assign micromat[16][50] = 9'b111111111;
assign micromat[16][51] = 9'b111111111;
assign micromat[16][52] = 9'b111111111;
assign micromat[16][53] = 9'b111111111;
assign micromat[16][54] = 9'b111111111;
assign micromat[16][55] = 9'b111111111;
assign micromat[16][56] = 9'b111111111;
assign micromat[16][57] = 9'b111111111;
assign micromat[16][58] = 9'b111111111;
assign micromat[16][59] = 9'b111111111;
assign micromat[16][60] = 9'b111111111;
assign micromat[16][61] = 9'b111111111;
assign micromat[16][62] = 9'b111111111;
assign micromat[16][63] = 9'b111111111;
assign micromat[16][64] = 9'b111111111;
assign micromat[16][65] = 9'b111111111;
assign micromat[16][66] = 9'b111111111;
assign micromat[16][67] = 9'b111111111;
assign micromat[16][68] = 9'b111111111;
assign micromat[16][69] = 9'b111111111;
assign micromat[16][70] = 9'b111111111;
assign micromat[16][71] = 9'b111111111;
assign micromat[16][72] = 9'b111111111;
assign micromat[16][73] = 9'b111111111;
assign micromat[16][74] = 9'b111111111;
assign micromat[16][75] = 9'b111111111;
assign micromat[16][76] = 9'b111111111;
assign micromat[16][77] = 9'b111111111;
assign micromat[16][78] = 9'b111111111;
assign micromat[16][79] = 9'b111111111;
assign micromat[16][80] = 9'b111111111;
assign micromat[16][81] = 9'b111111111;
assign micromat[16][82] = 9'b111111111;
assign micromat[16][83] = 9'b111111111;
assign micromat[16][84] = 9'b111111111;
assign micromat[16][85] = 9'b111111111;
assign micromat[16][86] = 9'b111111111;
assign micromat[16][87] = 9'b111111111;
assign micromat[16][88] = 9'b111111111;
assign micromat[16][89] = 9'b111111111;
assign micromat[16][90] = 9'b111111111;
assign micromat[16][91] = 9'b111111111;
assign micromat[16][92] = 9'b111111111;
assign micromat[16][93] = 9'b111111111;
assign micromat[16][94] = 9'b111111111;
assign micromat[16][95] = 9'b111111111;
assign micromat[16][96] = 9'b111111111;
assign micromat[16][97] = 9'b111111111;
assign micromat[16][98] = 9'b111111111;
assign micromat[16][99] = 9'b111111111;
assign micromat[17][0] = 9'b111111111;
assign micromat[17][1] = 9'b111111111;
assign micromat[17][2] = 9'b111111111;
assign micromat[17][3] = 9'b111111111;
assign micromat[17][4] = 9'b111111111;
assign micromat[17][5] = 9'b111111111;
assign micromat[17][6] = 9'b111111111;
assign micromat[17][7] = 9'b111111111;
assign micromat[17][8] = 9'b111111111;
assign micromat[17][9] = 9'b111111111;
assign micromat[17][10] = 9'b111111111;
assign micromat[17][11] = 9'b111111111;
assign micromat[17][12] = 9'b111111111;
assign micromat[17][13] = 9'b111111111;
assign micromat[17][14] = 9'b111111111;
assign micromat[17][15] = 9'b111111111;
assign micromat[17][16] = 9'b111111111;
assign micromat[17][17] = 9'b111111111;
assign micromat[17][18] = 9'b111111111;
assign micromat[17][19] = 9'b111111111;
assign micromat[17][20] = 9'b111111111;
assign micromat[17][21] = 9'b111111111;
assign micromat[17][22] = 9'b111111111;
assign micromat[17][23] = 9'b111111111;
assign micromat[17][24] = 9'b111111111;
assign micromat[17][25] = 9'b111111111;
assign micromat[17][26] = 9'b111111111;
assign micromat[17][27] = 9'b111111111;
assign micromat[17][28] = 9'b111111111;
assign micromat[17][29] = 9'b111111111;
assign micromat[17][30] = 9'b111111111;
assign micromat[17][31] = 9'b111111111;
assign micromat[17][32] = 9'b111111111;
assign micromat[17][33] = 9'b111111111;
assign micromat[17][34] = 9'b111111111;
assign micromat[17][35] = 9'b111111111;
assign micromat[17][36] = 9'b111111111;
assign micromat[17][37] = 9'b111111111;
assign micromat[17][38] = 9'b111111111;
assign micromat[17][39] = 9'b111111111;
assign micromat[17][40] = 9'b111111111;
assign micromat[17][41] = 9'b111111111;
assign micromat[17][42] = 9'b111111111;
assign micromat[17][43] = 9'b111111111;
assign micromat[17][44] = 9'b111111111;
assign micromat[17][45] = 9'b111111111;
assign micromat[17][46] = 9'b111111111;
assign micromat[17][47] = 9'b111111111;
assign micromat[17][48] = 9'b111111111;
assign micromat[17][49] = 9'b111111111;
assign micromat[17][50] = 9'b111111111;
assign micromat[17][51] = 9'b111111111;
assign micromat[17][52] = 9'b111111111;
assign micromat[17][53] = 9'b111111111;
assign micromat[17][54] = 9'b111111111;
assign micromat[17][55] = 9'b111111111;
assign micromat[17][56] = 9'b111111111;
assign micromat[17][57] = 9'b111111111;
assign micromat[17][58] = 9'b111111111;
assign micromat[17][59] = 9'b111111111;
assign micromat[17][60] = 9'b111111111;
assign micromat[17][61] = 9'b111111111;
assign micromat[17][62] = 9'b111111111;
assign micromat[17][63] = 9'b111111111;
assign micromat[17][64] = 9'b111111111;
assign micromat[17][65] = 9'b111111111;
assign micromat[17][66] = 9'b111111111;
assign micromat[17][67] = 9'b111111111;
assign micromat[17][68] = 9'b111111111;
assign micromat[17][69] = 9'b111111111;
assign micromat[17][70] = 9'b111111111;
assign micromat[17][71] = 9'b111111111;
assign micromat[17][72] = 9'b111111111;
assign micromat[17][73] = 9'b111111111;
assign micromat[17][74] = 9'b111111111;
assign micromat[17][75] = 9'b111111111;
assign micromat[17][76] = 9'b111111111;
assign micromat[17][77] = 9'b111111111;
assign micromat[17][78] = 9'b111111111;
assign micromat[17][79] = 9'b111111111;
assign micromat[17][80] = 9'b111111111;
assign micromat[17][81] = 9'b111111111;
assign micromat[17][82] = 9'b111111111;
assign micromat[17][83] = 9'b111111111;
assign micromat[17][84] = 9'b111111111;
assign micromat[17][85] = 9'b111111111;
assign micromat[17][86] = 9'b111111111;
assign micromat[17][87] = 9'b111111111;
assign micromat[17][88] = 9'b111111111;
assign micromat[17][89] = 9'b111111111;
assign micromat[17][90] = 9'b111111111;
assign micromat[17][91] = 9'b111111111;
assign micromat[17][92] = 9'b111111111;
assign micromat[17][93] = 9'b111111111;
assign micromat[17][94] = 9'b111111111;
assign micromat[17][95] = 9'b111111111;
assign micromat[17][96] = 9'b111111111;
assign micromat[17][97] = 9'b111111111;
assign micromat[17][98] = 9'b111111111;
assign micromat[17][99] = 9'b111111111;
assign micromat[18][0] = 9'b111111111;
assign micromat[18][1] = 9'b111111111;
assign micromat[18][2] = 9'b111111111;
assign micromat[18][3] = 9'b111111111;
assign micromat[18][4] = 9'b111111111;
assign micromat[18][5] = 9'b111111111;
assign micromat[18][6] = 9'b111111111;
assign micromat[18][7] = 9'b111111111;
assign micromat[18][8] = 9'b111111111;
assign micromat[18][9] = 9'b111111111;
assign micromat[18][10] = 9'b111111111;
assign micromat[18][11] = 9'b111111111;
assign micromat[18][12] = 9'b111111111;
assign micromat[18][13] = 9'b111111111;
assign micromat[18][14] = 9'b111111111;
assign micromat[18][15] = 9'b111111111;
assign micromat[18][16] = 9'b111111111;
assign micromat[18][17] = 9'b111111111;
assign micromat[18][18] = 9'b111111111;
assign micromat[18][19] = 9'b111111111;
assign micromat[18][20] = 9'b111111111;
assign micromat[18][21] = 9'b111111111;
assign micromat[18][22] = 9'b111111111;
assign micromat[18][23] = 9'b111111111;
assign micromat[18][24] = 9'b111111111;
assign micromat[18][25] = 9'b111111111;
assign micromat[18][26] = 9'b111111111;
assign micromat[18][27] = 9'b111111111;
assign micromat[18][28] = 9'b111111111;
assign micromat[18][29] = 9'b111111111;
assign micromat[18][30] = 9'b111111111;
assign micromat[18][31] = 9'b111111111;
assign micromat[18][32] = 9'b111111111;
assign micromat[18][33] = 9'b111111111;
assign micromat[18][34] = 9'b111111111;
assign micromat[18][35] = 9'b111111111;
assign micromat[18][36] = 9'b111111111;
assign micromat[18][37] = 9'b111111111;
assign micromat[18][38] = 9'b111111111;
assign micromat[18][39] = 9'b111111111;
assign micromat[18][40] = 9'b111111111;
assign micromat[18][41] = 9'b111111111;
assign micromat[18][42] = 9'b111111111;
assign micromat[18][43] = 9'b111111111;
assign micromat[18][44] = 9'b111111111;
assign micromat[18][45] = 9'b111111111;
assign micromat[18][46] = 9'b111111111;
assign micromat[18][47] = 9'b111111111;
assign micromat[18][48] = 9'b111111111;
assign micromat[18][49] = 9'b111111111;
assign micromat[18][50] = 9'b111111111;
assign micromat[18][51] = 9'b111111111;
assign micromat[18][52] = 9'b111111111;
assign micromat[18][53] = 9'b111111111;
assign micromat[18][54] = 9'b111111111;
assign micromat[18][55] = 9'b111111111;
assign micromat[18][56] = 9'b111111111;
assign micromat[18][57] = 9'b111111111;
assign micromat[18][58] = 9'b111111111;
assign micromat[18][59] = 9'b111111111;
assign micromat[18][60] = 9'b111111111;
assign micromat[18][61] = 9'b111111111;
assign micromat[18][62] = 9'b111111111;
assign micromat[18][63] = 9'b111111111;
assign micromat[18][64] = 9'b111111111;
assign micromat[18][65] = 9'b111111111;
assign micromat[18][66] = 9'b111111111;
assign micromat[18][67] = 9'b111111111;
assign micromat[18][68] = 9'b111111111;
assign micromat[18][69] = 9'b111111111;
assign micromat[18][70] = 9'b111111111;
assign micromat[18][71] = 9'b111111111;
assign micromat[18][72] = 9'b111111111;
assign micromat[18][73] = 9'b111111111;
assign micromat[18][74] = 9'b111111111;
assign micromat[18][75] = 9'b111111111;
assign micromat[18][76] = 9'b111111111;
assign micromat[18][77] = 9'b111111111;
assign micromat[18][78] = 9'b111111111;
assign micromat[18][79] = 9'b111111111;
assign micromat[18][80] = 9'b111111111;
assign micromat[18][81] = 9'b111111111;
assign micromat[18][82] = 9'b111111111;
assign micromat[18][83] = 9'b111111111;
assign micromat[18][84] = 9'b111111111;
assign micromat[18][85] = 9'b111111111;
assign micromat[18][86] = 9'b111111111;
assign micromat[18][87] = 9'b111111111;
assign micromat[18][88] = 9'b111111111;
assign micromat[18][89] = 9'b111111111;
assign micromat[18][90] = 9'b111111111;
assign micromat[18][91] = 9'b111111111;
assign micromat[18][92] = 9'b111111111;
assign micromat[18][93] = 9'b111111111;
assign micromat[18][94] = 9'b111111111;
assign micromat[18][95] = 9'b111111111;
assign micromat[18][96] = 9'b111111111;
assign micromat[18][97] = 9'b111111111;
assign micromat[18][98] = 9'b111111111;
assign micromat[18][99] = 9'b111111111;
assign micromat[19][0] = 9'b111111111;
assign micromat[19][1] = 9'b111111111;
assign micromat[19][2] = 9'b111111111;
assign micromat[19][3] = 9'b111111111;
assign micromat[19][4] = 9'b111111111;
assign micromat[19][5] = 9'b111111111;
assign micromat[19][6] = 9'b111111111;
assign micromat[19][7] = 9'b111111111;
assign micromat[19][8] = 9'b111111111;
assign micromat[19][9] = 9'b111111111;
assign micromat[19][10] = 9'b111111111;
assign micromat[19][11] = 9'b111111111;
assign micromat[19][12] = 9'b111111111;
assign micromat[19][13] = 9'b111111111;
assign micromat[19][14] = 9'b111111111;
assign micromat[19][15] = 9'b111111111;
assign micromat[19][16] = 9'b111111111;
assign micromat[19][17] = 9'b111111111;
assign micromat[19][18] = 9'b111111111;
assign micromat[19][19] = 9'b111111111;
assign micromat[19][20] = 9'b111111111;
assign micromat[19][21] = 9'b111111111;
assign micromat[19][22] = 9'b111111111;
assign micromat[19][23] = 9'b111111111;
assign micromat[19][24] = 9'b111111111;
assign micromat[19][25] = 9'b111111111;
assign micromat[19][26] = 9'b111111111;
assign micromat[19][27] = 9'b111111111;
assign micromat[19][28] = 9'b111111111;
assign micromat[19][29] = 9'b111111111;
assign micromat[19][30] = 9'b111111111;
assign micromat[19][31] = 9'b111111111;
assign micromat[19][32] = 9'b111111111;
assign micromat[19][33] = 9'b111111111;
assign micromat[19][34] = 9'b111111111;
assign micromat[19][35] = 9'b111111111;
assign micromat[19][36] = 9'b111111111;
assign micromat[19][37] = 9'b111111111;
assign micromat[19][38] = 9'b111111111;
assign micromat[19][39] = 9'b111111111;
assign micromat[19][40] = 9'b111111111;
assign micromat[19][41] = 9'b111111111;
assign micromat[19][42] = 9'b111111111;
assign micromat[19][43] = 9'b111111111;
assign micromat[19][44] = 9'b111111111;
assign micromat[19][45] = 9'b111111111;
assign micromat[19][46] = 9'b111111111;
assign micromat[19][47] = 9'b111111111;
assign micromat[19][48] = 9'b111111111;
assign micromat[19][49] = 9'b111111111;
assign micromat[19][50] = 9'b111111111;
assign micromat[19][51] = 9'b111111111;
assign micromat[19][52] = 9'b111111111;
assign micromat[19][53] = 9'b111111111;
assign micromat[19][54] = 9'b111111111;
assign micromat[19][55] = 9'b111111111;
assign micromat[19][56] = 9'b111111111;
assign micromat[19][57] = 9'b111111111;
assign micromat[19][58] = 9'b111111111;
assign micromat[19][59] = 9'b111111111;
assign micromat[19][60] = 9'b111111111;
assign micromat[19][61] = 9'b111111111;
assign micromat[19][62] = 9'b111111111;
assign micromat[19][63] = 9'b111111111;
assign micromat[19][64] = 9'b111111111;
assign micromat[19][65] = 9'b111111111;
assign micromat[19][66] = 9'b111111111;
assign micromat[19][67] = 9'b111111111;
assign micromat[19][68] = 9'b111111111;
assign micromat[19][69] = 9'b111111111;
assign micromat[19][70] = 9'b111111111;
assign micromat[19][71] = 9'b111111111;
assign micromat[19][72] = 9'b111111111;
assign micromat[19][73] = 9'b111111111;
assign micromat[19][74] = 9'b111111111;
assign micromat[19][75] = 9'b111111111;
assign micromat[19][76] = 9'b111111111;
assign micromat[19][77] = 9'b111111111;
assign micromat[19][78] = 9'b111111111;
assign micromat[19][79] = 9'b111111111;
assign micromat[19][80] = 9'b111111111;
assign micromat[19][81] = 9'b111111111;
assign micromat[19][82] = 9'b111111111;
assign micromat[19][83] = 9'b111111111;
assign micromat[19][84] = 9'b111111111;
assign micromat[19][85] = 9'b111111111;
assign micromat[19][86] = 9'b111111111;
assign micromat[19][87] = 9'b111111111;
assign micromat[19][88] = 9'b111111111;
assign micromat[19][89] = 9'b111111111;
assign micromat[19][90] = 9'b111111111;
assign micromat[19][91] = 9'b111111111;
assign micromat[19][92] = 9'b111111111;
assign micromat[19][93] = 9'b111111111;
assign micromat[19][94] = 9'b111111111;
assign micromat[19][95] = 9'b111111111;
assign micromat[19][96] = 9'b111111111;
assign micromat[19][97] = 9'b111111111;
assign micromat[19][98] = 9'b111111111;
assign micromat[19][99] = 9'b111111111;
assign micromat[20][0] = 9'b111111111;
assign micromat[20][1] = 9'b111111111;
assign micromat[20][2] = 9'b111111111;
assign micromat[20][3] = 9'b111111111;
assign micromat[20][4] = 9'b111111111;
assign micromat[20][5] = 9'b111111111;
assign micromat[20][6] = 9'b111111111;
assign micromat[20][7] = 9'b111111111;
assign micromat[20][8] = 9'b111111111;
assign micromat[20][9] = 9'b111111111;
assign micromat[20][10] = 9'b111111111;
assign micromat[20][11] = 9'b111111111;
assign micromat[20][12] = 9'b111111111;
assign micromat[20][13] = 9'b111111111;
assign micromat[20][14] = 9'b111111111;
assign micromat[20][15] = 9'b111111111;
assign micromat[20][16] = 9'b111111111;
assign micromat[20][17] = 9'b111111111;
assign micromat[20][18] = 9'b111111111;
assign micromat[20][19] = 9'b111111111;
assign micromat[20][20] = 9'b111111111;
assign micromat[20][21] = 9'b111111111;
assign micromat[20][22] = 9'b111111111;
assign micromat[20][23] = 9'b111111111;
assign micromat[20][24] = 9'b111111111;
assign micromat[20][25] = 9'b111111111;
assign micromat[20][26] = 9'b111111111;
assign micromat[20][27] = 9'b111111111;
assign micromat[20][28] = 9'b111111111;
assign micromat[20][29] = 9'b111111111;
assign micromat[20][30] = 9'b111111111;
assign micromat[20][31] = 9'b111111111;
assign micromat[20][32] = 9'b111111111;
assign micromat[20][33] = 9'b111111111;
assign micromat[20][34] = 9'b111111111;
assign micromat[20][35] = 9'b111111111;
assign micromat[20][36] = 9'b111111111;
assign micromat[20][37] = 9'b111111111;
assign micromat[20][38] = 9'b111111111;
assign micromat[20][39] = 9'b111111111;
assign micromat[20][40] = 9'b111111111;
assign micromat[20][41] = 9'b111111111;
assign micromat[20][42] = 9'b111111111;
assign micromat[20][43] = 9'b111111111;
assign micromat[20][44] = 9'b111111111;
assign micromat[20][45] = 9'b111111111;
assign micromat[20][46] = 9'b111111111;
assign micromat[20][47] = 9'b111111111;
assign micromat[20][48] = 9'b111111111;
assign micromat[20][49] = 9'b111111111;
assign micromat[20][50] = 9'b111111111;
assign micromat[20][51] = 9'b111111111;
assign micromat[20][52] = 9'b111111111;
assign micromat[20][53] = 9'b111111111;
assign micromat[20][54] = 9'b111111111;
assign micromat[20][55] = 9'b111111111;
assign micromat[20][56] = 9'b111111111;
assign micromat[20][57] = 9'b111111111;
assign micromat[20][58] = 9'b111111111;
assign micromat[20][59] = 9'b111111111;
assign micromat[20][60] = 9'b111111111;
assign micromat[20][61] = 9'b111111111;
assign micromat[20][62] = 9'b111111111;
assign micromat[20][63] = 9'b111111111;
assign micromat[20][64] = 9'b111111111;
assign micromat[20][65] = 9'b111111111;
assign micromat[20][66] = 9'b111111111;
assign micromat[20][67] = 9'b111111111;
assign micromat[20][68] = 9'b111111111;
assign micromat[20][69] = 9'b111111111;
assign micromat[20][70] = 9'b111111111;
assign micromat[20][71] = 9'b111111111;
assign micromat[20][72] = 9'b111111111;
assign micromat[20][73] = 9'b111111111;
assign micromat[20][74] = 9'b111111111;
assign micromat[20][75] = 9'b111111111;
assign micromat[20][76] = 9'b111111111;
assign micromat[20][77] = 9'b111111111;
assign micromat[20][78] = 9'b111111111;
assign micromat[20][79] = 9'b111111111;
assign micromat[20][80] = 9'b111111111;
assign micromat[20][81] = 9'b111111111;
assign micromat[20][82] = 9'b111111111;
assign micromat[20][83] = 9'b111111111;
assign micromat[20][84] = 9'b111111111;
assign micromat[20][85] = 9'b111111111;
assign micromat[20][86] = 9'b111111111;
assign micromat[20][87] = 9'b111111111;
assign micromat[20][88] = 9'b111111111;
assign micromat[20][89] = 9'b111111111;
assign micromat[20][90] = 9'b111111111;
assign micromat[20][91] = 9'b111111111;
assign micromat[20][92] = 9'b111111111;
assign micromat[20][93] = 9'b111111111;
assign micromat[20][94] = 9'b111111111;
assign micromat[20][95] = 9'b111111111;
assign micromat[20][96] = 9'b111111111;
assign micromat[20][97] = 9'b111111111;
assign micromat[20][98] = 9'b111111111;
assign micromat[20][99] = 9'b111111111;
assign micromat[21][0] = 9'b111111111;
assign micromat[21][1] = 9'b111111111;
assign micromat[21][2] = 9'b111111111;
assign micromat[21][3] = 9'b111111111;
assign micromat[21][4] = 9'b111111111;
assign micromat[21][5] = 9'b111111111;
assign micromat[21][6] = 9'b111111111;
assign micromat[21][7] = 9'b111111111;
assign micromat[21][8] = 9'b111111111;
assign micromat[21][9] = 9'b111111111;
assign micromat[21][10] = 9'b111111111;
assign micromat[21][11] = 9'b111111111;
assign micromat[21][12] = 9'b111111111;
assign micromat[21][13] = 9'b111111111;
assign micromat[21][14] = 9'b111111111;
assign micromat[21][15] = 9'b111111111;
assign micromat[21][16] = 9'b111111111;
assign micromat[21][17] = 9'b111111111;
assign micromat[21][18] = 9'b111111111;
assign micromat[21][19] = 9'b111111111;
assign micromat[21][20] = 9'b111111111;
assign micromat[21][21] = 9'b111111111;
assign micromat[21][22] = 9'b111111111;
assign micromat[21][23] = 9'b111111111;
assign micromat[21][24] = 9'b111111111;
assign micromat[21][25] = 9'b111111111;
assign micromat[21][26] = 9'b111111111;
assign micromat[21][27] = 9'b111111111;
assign micromat[21][28] = 9'b111111111;
assign micromat[21][29] = 9'b111111111;
assign micromat[21][30] = 9'b111111111;
assign micromat[21][31] = 9'b111111111;
assign micromat[21][32] = 9'b111111111;
assign micromat[21][33] = 9'b111111111;
assign micromat[21][34] = 9'b111111111;
assign micromat[21][35] = 9'b111111111;
assign micromat[21][36] = 9'b111111111;
assign micromat[21][37] = 9'b111111111;
assign micromat[21][38] = 9'b111111111;
assign micromat[21][39] = 9'b111111111;
assign micromat[21][40] = 9'b111111111;
assign micromat[21][41] = 9'b111111111;
assign micromat[21][42] = 9'b111111111;
assign micromat[21][43] = 9'b111111111;
assign micromat[21][44] = 9'b111111111;
assign micromat[21][45] = 9'b111111111;
assign micromat[21][46] = 9'b111111111;
assign micromat[21][47] = 9'b111111111;
assign micromat[21][48] = 9'b111111111;
assign micromat[21][49] = 9'b111111111;
assign micromat[21][50] = 9'b111111111;
assign micromat[21][51] = 9'b111111111;
assign micromat[21][52] = 9'b111111111;
assign micromat[21][53] = 9'b111111111;
assign micromat[21][54] = 9'b111111111;
assign micromat[21][55] = 9'b111111111;
assign micromat[21][56] = 9'b111111111;
assign micromat[21][57] = 9'b111111111;
assign micromat[21][58] = 9'b111111111;
assign micromat[21][59] = 9'b111111111;
assign micromat[21][60] = 9'b111111111;
assign micromat[21][61] = 9'b111111111;
assign micromat[21][62] = 9'b111111111;
assign micromat[21][63] = 9'b111111111;
assign micromat[21][64] = 9'b111111111;
assign micromat[21][65] = 9'b111111111;
assign micromat[21][66] = 9'b111111111;
assign micromat[21][67] = 9'b111111111;
assign micromat[21][68] = 9'b111111111;
assign micromat[21][69] = 9'b111111111;
assign micromat[21][70] = 9'b111111111;
assign micromat[21][71] = 9'b111111111;
assign micromat[21][72] = 9'b111111111;
assign micromat[21][73] = 9'b111111111;
assign micromat[21][74] = 9'b111111111;
assign micromat[21][75] = 9'b111111111;
assign micromat[21][76] = 9'b111111111;
assign micromat[21][77] = 9'b111111111;
assign micromat[21][78] = 9'b111111111;
assign micromat[21][79] = 9'b111111111;
assign micromat[21][80] = 9'b111111111;
assign micromat[21][81] = 9'b111111111;
assign micromat[21][82] = 9'b111111111;
assign micromat[21][83] = 9'b111111111;
assign micromat[21][84] = 9'b111111111;
assign micromat[21][85] = 9'b111111111;
assign micromat[21][86] = 9'b111111111;
assign micromat[21][87] = 9'b111111111;
assign micromat[21][88] = 9'b111111111;
assign micromat[21][89] = 9'b111111111;
assign micromat[21][90] = 9'b111111111;
assign micromat[21][91] = 9'b111111111;
assign micromat[21][92] = 9'b111111111;
assign micromat[21][93] = 9'b111111111;
assign micromat[21][94] = 9'b111111111;
assign micromat[21][95] = 9'b111111111;
assign micromat[21][96] = 9'b111111111;
assign micromat[21][97] = 9'b111111111;
assign micromat[21][98] = 9'b111111111;
assign micromat[21][99] = 9'b111111111;
assign micromat[22][0] = 9'b111111111;
assign micromat[22][1] = 9'b111111111;
assign micromat[22][2] = 9'b111111111;
assign micromat[22][3] = 9'b111111111;
assign micromat[22][4] = 9'b111111111;
assign micromat[22][5] = 9'b111111111;
assign micromat[22][6] = 9'b111111111;
assign micromat[22][7] = 9'b111111111;
assign micromat[22][8] = 9'b111111111;
assign micromat[22][9] = 9'b111111111;
assign micromat[22][10] = 9'b111111111;
assign micromat[22][11] = 9'b111111111;
assign micromat[22][12] = 9'b111111111;
assign micromat[22][13] = 9'b111111111;
assign micromat[22][14] = 9'b111111111;
assign micromat[22][15] = 9'b111111111;
assign micromat[22][16] = 9'b111111111;
assign micromat[22][17] = 9'b111111111;
assign micromat[22][18] = 9'b111111111;
assign micromat[22][19] = 9'b111111111;
assign micromat[22][20] = 9'b111111111;
assign micromat[22][21] = 9'b111111111;
assign micromat[22][22] = 9'b111111111;
assign micromat[22][23] = 9'b111111111;
assign micromat[22][24] = 9'b111111111;
assign micromat[22][25] = 9'b111111111;
assign micromat[22][26] = 9'b111111111;
assign micromat[22][27] = 9'b111111111;
assign micromat[22][28] = 9'b111111111;
assign micromat[22][29] = 9'b111111111;
assign micromat[22][30] = 9'b111111111;
assign micromat[22][31] = 9'b111111111;
assign micromat[22][32] = 9'b111111111;
assign micromat[22][33] = 9'b111111111;
assign micromat[22][34] = 9'b111111111;
assign micromat[22][35] = 9'b111111111;
assign micromat[22][36] = 9'b111111111;
assign micromat[22][37] = 9'b111111111;
assign micromat[22][38] = 9'b111111111;
assign micromat[22][39] = 9'b111111111;
assign micromat[22][40] = 9'b111111111;
assign micromat[22][41] = 9'b111111111;
assign micromat[22][42] = 9'b111111111;
assign micromat[22][43] = 9'b111111111;
assign micromat[22][44] = 9'b111111111;
assign micromat[22][45] = 9'b111111111;
assign micromat[22][46] = 9'b111111111;
assign micromat[22][47] = 9'b111111111;
assign micromat[22][48] = 9'b111111111;
assign micromat[22][49] = 9'b111111111;
assign micromat[22][50] = 9'b111111111;
assign micromat[22][51] = 9'b111111111;
assign micromat[22][52] = 9'b111111111;
assign micromat[22][53] = 9'b111111111;
assign micromat[22][54] = 9'b111111111;
assign micromat[22][55] = 9'b111111111;
assign micromat[22][56] = 9'b111111111;
assign micromat[22][57] = 9'b111111111;
assign micromat[22][58] = 9'b111111111;
assign micromat[22][59] = 9'b111111111;
assign micromat[22][60] = 9'b111111111;
assign micromat[22][61] = 9'b111111111;
assign micromat[22][62] = 9'b111111111;
assign micromat[22][63] = 9'b111111111;
assign micromat[22][64] = 9'b111111111;
assign micromat[22][65] = 9'b111111111;
assign micromat[22][66] = 9'b111111111;
assign micromat[22][67] = 9'b111111111;
assign micromat[22][68] = 9'b111111111;
assign micromat[22][69] = 9'b111111111;
assign micromat[22][70] = 9'b111111111;
assign micromat[22][71] = 9'b111111111;
assign micromat[22][72] = 9'b111111111;
assign micromat[22][73] = 9'b111111111;
assign micromat[22][74] = 9'b111111111;
assign micromat[22][75] = 9'b111111111;
assign micromat[22][76] = 9'b111111111;
assign micromat[22][77] = 9'b111111111;
assign micromat[22][78] = 9'b111111111;
assign micromat[22][79] = 9'b111111111;
assign micromat[22][80] = 9'b111111111;
assign micromat[22][81] = 9'b111111111;
assign micromat[22][82] = 9'b111111111;
assign micromat[22][83] = 9'b111111111;
assign micromat[22][84] = 9'b111111111;
assign micromat[22][85] = 9'b111111111;
assign micromat[22][86] = 9'b111111111;
assign micromat[22][87] = 9'b111111111;
assign micromat[22][88] = 9'b111111111;
assign micromat[22][89] = 9'b111111111;
assign micromat[22][90] = 9'b111111111;
assign micromat[22][91] = 9'b111111111;
assign micromat[22][92] = 9'b111111111;
assign micromat[22][93] = 9'b111111111;
assign micromat[22][94] = 9'b111111111;
assign micromat[22][95] = 9'b111111111;
assign micromat[22][96] = 9'b111111111;
assign micromat[22][97] = 9'b111111111;
assign micromat[22][98] = 9'b111111111;
assign micromat[22][99] = 9'b111111111;
assign micromat[23][0] = 9'b111111111;
assign micromat[23][1] = 9'b111111111;
assign micromat[23][2] = 9'b111111111;
assign micromat[23][3] = 9'b111111111;
assign micromat[23][4] = 9'b111111111;
assign micromat[23][5] = 9'b111111111;
assign micromat[23][6] = 9'b111111111;
assign micromat[23][7] = 9'b111111111;
assign micromat[23][8] = 9'b111111111;
assign micromat[23][9] = 9'b111111111;
assign micromat[23][10] = 9'b111111111;
assign micromat[23][11] = 9'b111111111;
assign micromat[23][12] = 9'b111111111;
assign micromat[23][13] = 9'b111111111;
assign micromat[23][14] = 9'b111111111;
assign micromat[23][15] = 9'b111111111;
assign micromat[23][16] = 9'b111111111;
assign micromat[23][17] = 9'b111111111;
assign micromat[23][18] = 9'b111111111;
assign micromat[23][19] = 9'b111111111;
assign micromat[23][20] = 9'b111111111;
assign micromat[23][21] = 9'b111111111;
assign micromat[23][22] = 9'b111111111;
assign micromat[23][23] = 9'b111111111;
assign micromat[23][24] = 9'b111111111;
assign micromat[23][25] = 9'b111111111;
assign micromat[23][26] = 9'b111111111;
assign micromat[23][27] = 9'b111111111;
assign micromat[23][28] = 9'b111111111;
assign micromat[23][29] = 9'b111111111;
assign micromat[23][30] = 9'b111111111;
assign micromat[23][31] = 9'b111111111;
assign micromat[23][32] = 9'b111111111;
assign micromat[23][33] = 9'b111111111;
assign micromat[23][34] = 9'b111111111;
assign micromat[23][35] = 9'b111111111;
assign micromat[23][36] = 9'b111111111;
assign micromat[23][37] = 9'b111111111;
assign micromat[23][38] = 9'b111111111;
assign micromat[23][39] = 9'b111111111;
assign micromat[23][40] = 9'b111111111;
assign micromat[23][41] = 9'b111111111;
assign micromat[23][42] = 9'b111111111;
assign micromat[23][43] = 9'b111111111;
assign micromat[23][44] = 9'b111111111;
assign micromat[23][45] = 9'b111111111;
assign micromat[23][46] = 9'b111111111;
assign micromat[23][47] = 9'b111111111;
assign micromat[23][48] = 9'b111111111;
assign micromat[23][49] = 9'b111111111;
assign micromat[23][50] = 9'b111111111;
assign micromat[23][51] = 9'b111111111;
assign micromat[23][52] = 9'b111111111;
assign micromat[23][53] = 9'b111111111;
assign micromat[23][54] = 9'b111111111;
assign micromat[23][55] = 9'b111111111;
assign micromat[23][56] = 9'b111111111;
assign micromat[23][57] = 9'b111111111;
assign micromat[23][58] = 9'b111111111;
assign micromat[23][59] = 9'b111111111;
assign micromat[23][60] = 9'b111111111;
assign micromat[23][61] = 9'b111111111;
assign micromat[23][62] = 9'b111111111;
assign micromat[23][63] = 9'b111111111;
assign micromat[23][64] = 9'b111111111;
assign micromat[23][65] = 9'b111111111;
assign micromat[23][66] = 9'b111111111;
assign micromat[23][67] = 9'b111111111;
assign micromat[23][68] = 9'b111111111;
assign micromat[23][69] = 9'b111111111;
assign micromat[23][70] = 9'b111111111;
assign micromat[23][71] = 9'b111111111;
assign micromat[23][72] = 9'b111111111;
assign micromat[23][73] = 9'b111111111;
assign micromat[23][74] = 9'b111111111;
assign micromat[23][75] = 9'b111111111;
assign micromat[23][76] = 9'b111111111;
assign micromat[23][77] = 9'b111111111;
assign micromat[23][78] = 9'b111111111;
assign micromat[23][79] = 9'b111111111;
assign micromat[23][80] = 9'b111111111;
assign micromat[23][81] = 9'b111111111;
assign micromat[23][82] = 9'b111111111;
assign micromat[23][83] = 9'b111111111;
assign micromat[23][84] = 9'b111111111;
assign micromat[23][85] = 9'b111111111;
assign micromat[23][86] = 9'b111111111;
assign micromat[23][87] = 9'b111111111;
assign micromat[23][88] = 9'b111111111;
assign micromat[23][89] = 9'b111111111;
assign micromat[23][90] = 9'b111111111;
assign micromat[23][91] = 9'b111111111;
assign micromat[23][92] = 9'b111111111;
assign micromat[23][93] = 9'b111111111;
assign micromat[23][94] = 9'b111111111;
assign micromat[23][95] = 9'b111111111;
assign micromat[23][96] = 9'b111111111;
assign micromat[23][97] = 9'b111111111;
assign micromat[23][98] = 9'b111111111;
assign micromat[23][99] = 9'b111111111;
assign micromat[24][0] = 9'b111111111;
assign micromat[24][1] = 9'b111111111;
assign micromat[24][2] = 9'b111111111;
assign micromat[24][3] = 9'b111111111;
assign micromat[24][4] = 9'b111111111;
assign micromat[24][5] = 9'b111111111;
assign micromat[24][6] = 9'b111111111;
assign micromat[24][7] = 9'b111111111;
assign micromat[24][8] = 9'b111111111;
assign micromat[24][9] = 9'b111111111;
assign micromat[24][10] = 9'b111111111;
assign micromat[24][11] = 9'b111111111;
assign micromat[24][12] = 9'b111111111;
assign micromat[24][13] = 9'b111111111;
assign micromat[24][14] = 9'b111111111;
assign micromat[24][15] = 9'b111111111;
assign micromat[24][16] = 9'b111111111;
assign micromat[24][17] = 9'b111111111;
assign micromat[24][18] = 9'b111111111;
assign micromat[24][19] = 9'b111111111;
assign micromat[24][20] = 9'b111111111;
assign micromat[24][21] = 9'b111111111;
assign micromat[24][22] = 9'b111111111;
assign micromat[24][23] = 9'b111111111;
assign micromat[24][24] = 9'b111111111;
assign micromat[24][25] = 9'b111111111;
assign micromat[24][26] = 9'b111111111;
assign micromat[24][27] = 9'b111111111;
assign micromat[24][28] = 9'b111111111;
assign micromat[24][29] = 9'b111111111;
assign micromat[24][30] = 9'b111111111;
assign micromat[24][31] = 9'b111111111;
assign micromat[24][32] = 9'b111111111;
assign micromat[24][33] = 9'b111111111;
assign micromat[24][34] = 9'b111111111;
assign micromat[24][35] = 9'b111111111;
assign micromat[24][36] = 9'b111111111;
assign micromat[24][37] = 9'b111111111;
assign micromat[24][38] = 9'b111111111;
assign micromat[24][39] = 9'b111111111;
assign micromat[24][40] = 9'b111111111;
assign micromat[24][41] = 9'b111111111;
assign micromat[24][42] = 9'b111111111;
assign micromat[24][43] = 9'b111111111;
assign micromat[24][44] = 9'b111111111;
assign micromat[24][45] = 9'b111111111;
assign micromat[24][46] = 9'b111111111;
assign micromat[24][47] = 9'b111111111;
assign micromat[24][48] = 9'b111111111;
assign micromat[24][49] = 9'b111111111;
assign micromat[24][50] = 9'b111111111;
assign micromat[24][51] = 9'b111111111;
assign micromat[24][52] = 9'b111111111;
assign micromat[24][53] = 9'b111111111;
assign micromat[24][54] = 9'b111111111;
assign micromat[24][55] = 9'b111111111;
assign micromat[24][56] = 9'b111111111;
assign micromat[24][57] = 9'b111111111;
assign micromat[24][58] = 9'b111111111;
assign micromat[24][59] = 9'b111111111;
assign micromat[24][60] = 9'b111111111;
assign micromat[24][61] = 9'b111111111;
assign micromat[24][62] = 9'b111111111;
assign micromat[24][63] = 9'b111111111;
assign micromat[24][64] = 9'b111111111;
assign micromat[24][65] = 9'b111111111;
assign micromat[24][66] = 9'b111111111;
assign micromat[24][67] = 9'b111111111;
assign micromat[24][68] = 9'b111111111;
assign micromat[24][69] = 9'b111111111;
assign micromat[24][70] = 9'b111111111;
assign micromat[24][71] = 9'b111111111;
assign micromat[24][72] = 9'b111111111;
assign micromat[24][73] = 9'b111111111;
assign micromat[24][74] = 9'b111111111;
assign micromat[24][75] = 9'b111111111;
assign micromat[24][76] = 9'b111111111;
assign micromat[24][77] = 9'b111111111;
assign micromat[24][78] = 9'b111111111;
assign micromat[24][79] = 9'b111111111;
assign micromat[24][80] = 9'b111111111;
assign micromat[24][81] = 9'b111111111;
assign micromat[24][82] = 9'b111111111;
assign micromat[24][83] = 9'b111111111;
assign micromat[24][84] = 9'b111111111;
assign micromat[24][85] = 9'b111111111;
assign micromat[24][86] = 9'b111111111;
assign micromat[24][87] = 9'b111111111;
assign micromat[24][88] = 9'b111111111;
assign micromat[24][89] = 9'b111111111;
assign micromat[24][90] = 9'b111111111;
assign micromat[24][91] = 9'b111111111;
assign micromat[24][92] = 9'b111111111;
assign micromat[24][93] = 9'b111111111;
assign micromat[24][94] = 9'b111111111;
assign micromat[24][95] = 9'b111111111;
assign micromat[24][96] = 9'b111111111;
assign micromat[24][97] = 9'b111111111;
assign micromat[24][98] = 9'b111111111;
assign micromat[24][99] = 9'b111111111;
assign micromat[25][0] = 9'b111111111;
assign micromat[25][1] = 9'b111111111;
assign micromat[25][2] = 9'b111111111;
assign micromat[25][3] = 9'b111111111;
assign micromat[25][4] = 9'b111111111;
assign micromat[25][5] = 9'b111111111;
assign micromat[25][6] = 9'b111111111;
assign micromat[25][7] = 9'b111111111;
assign micromat[25][8] = 9'b111111111;
assign micromat[25][9] = 9'b111111111;
assign micromat[25][10] = 9'b111111111;
assign micromat[25][11] = 9'b111111111;
assign micromat[25][12] = 9'b111111111;
assign micromat[25][13] = 9'b111111111;
assign micromat[25][14] = 9'b111111111;
assign micromat[25][15] = 9'b111111111;
assign micromat[25][16] = 9'b111111111;
assign micromat[25][17] = 9'b111111111;
assign micromat[25][18] = 9'b111111111;
assign micromat[25][19] = 9'b111111111;
assign micromat[25][20] = 9'b111111111;
assign micromat[25][21] = 9'b111111111;
assign micromat[25][22] = 9'b111111111;
assign micromat[25][23] = 9'b111111111;
assign micromat[25][24] = 9'b111111111;
assign micromat[25][25] = 9'b111111111;
assign micromat[25][26] = 9'b111111111;
assign micromat[25][27] = 9'b111111111;
assign micromat[25][28] = 9'b111111111;
assign micromat[25][29] = 9'b111111111;
assign micromat[25][30] = 9'b111111111;
assign micromat[25][31] = 9'b111111111;
assign micromat[25][32] = 9'b111111111;
assign micromat[25][33] = 9'b111111111;
assign micromat[25][34] = 9'b111111111;
assign micromat[25][35] = 9'b111111111;
assign micromat[25][36] = 9'b111111111;
assign micromat[25][37] = 9'b111111111;
assign micromat[25][38] = 9'b111111111;
assign micromat[25][39] = 9'b111111111;
assign micromat[25][40] = 9'b111111111;
assign micromat[25][41] = 9'b111111111;
assign micromat[25][42] = 9'b111111111;
assign micromat[25][43] = 9'b111111111;
assign micromat[25][44] = 9'b111111111;
assign micromat[25][45] = 9'b111111111;
assign micromat[25][46] = 9'b111111111;
assign micromat[25][47] = 9'b111111111;
assign micromat[25][48] = 9'b111111111;
assign micromat[25][49] = 9'b111111111;
assign micromat[25][50] = 9'b111111111;
assign micromat[25][51] = 9'b111111111;
assign micromat[25][52] = 9'b111111111;
assign micromat[25][53] = 9'b111111111;
assign micromat[25][54] = 9'b111111111;
assign micromat[25][55] = 9'b111111111;
assign micromat[25][56] = 9'b111111111;
assign micromat[25][57] = 9'b111111111;
assign micromat[25][58] = 9'b111111111;
assign micromat[25][59] = 9'b111111111;
assign micromat[25][60] = 9'b111111111;
assign micromat[25][61] = 9'b111111111;
assign micromat[25][62] = 9'b111111111;
assign micromat[25][63] = 9'b111111111;
assign micromat[25][64] = 9'b111111111;
assign micromat[25][65] = 9'b111111111;
assign micromat[25][66] = 9'b111111111;
assign micromat[25][67] = 9'b111111111;
assign micromat[25][68] = 9'b111111111;
assign micromat[25][69] = 9'b111111111;
assign micromat[25][70] = 9'b111111111;
assign micromat[25][71] = 9'b111111111;
assign micromat[25][72] = 9'b111111111;
assign micromat[25][73] = 9'b111111111;
assign micromat[25][74] = 9'b111111111;
assign micromat[25][75] = 9'b111111111;
assign micromat[25][76] = 9'b111111111;
assign micromat[25][77] = 9'b111111111;
assign micromat[25][78] = 9'b111111111;
assign micromat[25][79] = 9'b111111111;
assign micromat[25][80] = 9'b111111111;
assign micromat[25][81] = 9'b111111111;
assign micromat[25][82] = 9'b111111111;
assign micromat[25][83] = 9'b111111111;
assign micromat[25][84] = 9'b111111111;
assign micromat[25][85] = 9'b111111111;
assign micromat[25][86] = 9'b111111111;
assign micromat[25][87] = 9'b111111111;
assign micromat[25][88] = 9'b111111111;
assign micromat[25][89] = 9'b111111111;
assign micromat[25][90] = 9'b111111111;
assign micromat[25][91] = 9'b111111111;
assign micromat[25][92] = 9'b111111111;
assign micromat[25][93] = 9'b111111111;
assign micromat[25][94] = 9'b111111111;
assign micromat[25][95] = 9'b111111111;
assign micromat[25][96] = 9'b111111111;
assign micromat[25][97] = 9'b111111111;
assign micromat[25][98] = 9'b111111111;
assign micromat[25][99] = 9'b111111111;
assign micromat[26][0] = 9'b111111111;
assign micromat[26][1] = 9'b111111111;
assign micromat[26][2] = 9'b111111111;
assign micromat[26][3] = 9'b111111111;
assign micromat[26][4] = 9'b111111111;
assign micromat[26][5] = 9'b111111111;
assign micromat[26][6] = 9'b111111111;
assign micromat[26][7] = 9'b111111111;
assign micromat[26][8] = 9'b111111111;
assign micromat[26][9] = 9'b111111111;
assign micromat[26][10] = 9'b111111111;
assign micromat[26][11] = 9'b111111111;
assign micromat[26][12] = 9'b111111111;
assign micromat[26][13] = 9'b111111111;
assign micromat[26][14] = 9'b111111111;
assign micromat[26][15] = 9'b111111111;
assign micromat[26][16] = 9'b111111111;
assign micromat[26][17] = 9'b111111111;
assign micromat[26][18] = 9'b111111111;
assign micromat[26][19] = 9'b111111111;
assign micromat[26][20] = 9'b111111111;
assign micromat[26][21] = 9'b111111111;
assign micromat[26][22] = 9'b111111111;
assign micromat[26][23] = 9'b111111111;
assign micromat[26][24] = 9'b111111111;
assign micromat[26][25] = 9'b111111111;
assign micromat[26][26] = 9'b111111111;
assign micromat[26][27] = 9'b111111111;
assign micromat[26][28] = 9'b111111111;
assign micromat[26][29] = 9'b111111111;
assign micromat[26][30] = 9'b111111111;
assign micromat[26][31] = 9'b111111111;
assign micromat[26][32] = 9'b111111111;
assign micromat[26][33] = 9'b111111111;
assign micromat[26][34] = 9'b111111111;
assign micromat[26][35] = 9'b111111111;
assign micromat[26][36] = 9'b111111111;
assign micromat[26][37] = 9'b111111111;
assign micromat[26][38] = 9'b111111111;
assign micromat[26][39] = 9'b111111111;
assign micromat[26][40] = 9'b111111111;
assign micromat[26][41] = 9'b111111111;
assign micromat[26][42] = 9'b111111111;
assign micromat[26][43] = 9'b111111111;
assign micromat[26][44] = 9'b111111111;
assign micromat[26][45] = 9'b111111111;
assign micromat[26][46] = 9'b111111111;
assign micromat[26][47] = 9'b111111111;
assign micromat[26][48] = 9'b111111111;
assign micromat[26][49] = 9'b111111111;
assign micromat[26][50] = 9'b111111111;
assign micromat[26][51] = 9'b111111111;
assign micromat[26][52] = 9'b111111111;
assign micromat[26][53] = 9'b111111111;
assign micromat[26][54] = 9'b111111111;
assign micromat[26][55] = 9'b111111111;
assign micromat[26][56] = 9'b111111111;
assign micromat[26][57] = 9'b111111111;
assign micromat[26][58] = 9'b111111111;
assign micromat[26][59] = 9'b111111111;
assign micromat[26][60] = 9'b111111111;
assign micromat[26][61] = 9'b111111111;
assign micromat[26][62] = 9'b111111111;
assign micromat[26][63] = 9'b111111111;
assign micromat[26][64] = 9'b111111111;
assign micromat[26][65] = 9'b111111111;
assign micromat[26][66] = 9'b111111111;
assign micromat[26][67] = 9'b111111111;
assign micromat[26][68] = 9'b111111111;
assign micromat[26][69] = 9'b111111111;
assign micromat[26][70] = 9'b111111111;
assign micromat[26][71] = 9'b111111111;
assign micromat[26][72] = 9'b111111111;
assign micromat[26][73] = 9'b111111111;
assign micromat[26][74] = 9'b111111111;
assign micromat[26][75] = 9'b111111111;
assign micromat[26][76] = 9'b111111111;
assign micromat[26][77] = 9'b111111111;
assign micromat[26][78] = 9'b111111111;
assign micromat[26][79] = 9'b111111111;
assign micromat[26][80] = 9'b111111111;
assign micromat[26][81] = 9'b111111111;
assign micromat[26][82] = 9'b111111111;
assign micromat[26][83] = 9'b111111111;
assign micromat[26][84] = 9'b111111111;
assign micromat[26][85] = 9'b111111111;
assign micromat[26][86] = 9'b111111111;
assign micromat[26][87] = 9'b111111111;
assign micromat[26][88] = 9'b111111111;
assign micromat[26][89] = 9'b111111111;
assign micromat[26][90] = 9'b111111111;
assign micromat[26][91] = 9'b111111111;
assign micromat[26][92] = 9'b111111111;
assign micromat[26][93] = 9'b111111111;
assign micromat[26][94] = 9'b111111111;
assign micromat[26][95] = 9'b111111111;
assign micromat[26][96] = 9'b111111111;
assign micromat[26][97] = 9'b111111111;
assign micromat[26][98] = 9'b111111111;
assign micromat[26][99] = 9'b111111111;
assign micromat[27][0] = 9'b111111111;
assign micromat[27][1] = 9'b111111111;
assign micromat[27][2] = 9'b111111111;
assign micromat[27][3] = 9'b111111111;
assign micromat[27][4] = 9'b111111111;
assign micromat[27][5] = 9'b111111111;
assign micromat[27][6] = 9'b111111111;
assign micromat[27][7] = 9'b111111111;
assign micromat[27][8] = 9'b111111111;
assign micromat[27][9] = 9'b111111111;
assign micromat[27][10] = 9'b111111111;
assign micromat[27][11] = 9'b111111111;
assign micromat[27][12] = 9'b111111111;
assign micromat[27][13] = 9'b111111111;
assign micromat[27][14] = 9'b111111111;
assign micromat[27][15] = 9'b111111111;
assign micromat[27][16] = 9'b111111111;
assign micromat[27][17] = 9'b111111111;
assign micromat[27][18] = 9'b111111111;
assign micromat[27][19] = 9'b111111111;
assign micromat[27][20] = 9'b111111111;
assign micromat[27][21] = 9'b111111111;
assign micromat[27][22] = 9'b111111111;
assign micromat[27][23] = 9'b111111111;
assign micromat[27][24] = 9'b111111111;
assign micromat[27][25] = 9'b111111111;
assign micromat[27][26] = 9'b111111111;
assign micromat[27][27] = 9'b111111111;
assign micromat[27][28] = 9'b111111111;
assign micromat[27][29] = 9'b111111111;
assign micromat[27][30] = 9'b111111111;
assign micromat[27][31] = 9'b111111111;
assign micromat[27][32] = 9'b111111111;
assign micromat[27][33] = 9'b111111111;
assign micromat[27][34] = 9'b111111111;
assign micromat[27][35] = 9'b111111111;
assign micromat[27][36] = 9'b111111111;
assign micromat[27][37] = 9'b111111111;
assign micromat[27][38] = 9'b111111111;
assign micromat[27][39] = 9'b111111111;
assign micromat[27][40] = 9'b111111111;
assign micromat[27][41] = 9'b111111111;
assign micromat[27][42] = 9'b111111111;
assign micromat[27][43] = 9'b111111111;
assign micromat[27][44] = 9'b111111111;
assign micromat[27][45] = 9'b111111111;
assign micromat[27][46] = 9'b111111111;
assign micromat[27][47] = 9'b111111111;
assign micromat[27][48] = 9'b111111111;
assign micromat[27][49] = 9'b111111111;
assign micromat[27][50] = 9'b111111111;
assign micromat[27][51] = 9'b111111111;
assign micromat[27][52] = 9'b111111111;
assign micromat[27][53] = 9'b111111111;
assign micromat[27][54] = 9'b111111111;
assign micromat[27][55] = 9'b111111111;
assign micromat[27][56] = 9'b111111111;
assign micromat[27][57] = 9'b111111111;
assign micromat[27][58] = 9'b111111111;
assign micromat[27][59] = 9'b111111111;
assign micromat[27][60] = 9'b111111111;
assign micromat[27][61] = 9'b111111111;
assign micromat[27][62] = 9'b111111111;
assign micromat[27][63] = 9'b111111111;
assign micromat[27][64] = 9'b111111111;
assign micromat[27][65] = 9'b111111111;
assign micromat[27][66] = 9'b111111111;
assign micromat[27][67] = 9'b111111111;
assign micromat[27][68] = 9'b111111111;
assign micromat[27][69] = 9'b111111111;
assign micromat[27][70] = 9'b111111111;
assign micromat[27][71] = 9'b111111111;
assign micromat[27][72] = 9'b111111111;
assign micromat[27][73] = 9'b111111111;
assign micromat[27][74] = 9'b111111111;
assign micromat[27][75] = 9'b111111111;
assign micromat[27][76] = 9'b111111111;
assign micromat[27][77] = 9'b111111111;
assign micromat[27][78] = 9'b111111111;
assign micromat[27][79] = 9'b111111111;
assign micromat[27][80] = 9'b111111111;
assign micromat[27][81] = 9'b111111111;
assign micromat[27][82] = 9'b111111111;
assign micromat[27][83] = 9'b111111111;
assign micromat[27][84] = 9'b111111111;
assign micromat[27][85] = 9'b111111111;
assign micromat[27][86] = 9'b111111111;
assign micromat[27][87] = 9'b111111111;
assign micromat[27][88] = 9'b111111111;
assign micromat[27][89] = 9'b111111111;
assign micromat[27][90] = 9'b111111111;
assign micromat[27][91] = 9'b111111111;
assign micromat[27][92] = 9'b111111111;
assign micromat[27][93] = 9'b111111111;
assign micromat[27][94] = 9'b111111111;
assign micromat[27][95] = 9'b111111111;
assign micromat[27][96] = 9'b111111111;
assign micromat[27][97] = 9'b111111111;
assign micromat[27][98] = 9'b111111111;
assign micromat[27][99] = 9'b111111111;
assign micromat[28][0] = 9'b111111111;
assign micromat[28][1] = 9'b111111111;
assign micromat[28][2] = 9'b111111111;
assign micromat[28][3] = 9'b111111111;
assign micromat[28][4] = 9'b111111111;
assign micromat[28][5] = 9'b111111111;
assign micromat[28][6] = 9'b111111111;
assign micromat[28][7] = 9'b111111111;
assign micromat[28][8] = 9'b111111111;
assign micromat[28][9] = 9'b111111111;
assign micromat[28][10] = 9'b111111111;
assign micromat[28][11] = 9'b111111111;
assign micromat[28][12] = 9'b111111111;
assign micromat[28][13] = 9'b111111111;
assign micromat[28][14] = 9'b111111111;
assign micromat[28][15] = 9'b111111111;
assign micromat[28][16] = 9'b110110110;
assign micromat[28][17] = 9'b101101101;
assign micromat[28][18] = 9'b101101101;
assign micromat[28][19] = 9'b101101101;
assign micromat[28][20] = 9'b101101101;
assign micromat[28][21] = 9'b101101101;
assign micromat[28][22] = 9'b101101101;
assign micromat[28][23] = 9'b101101101;
assign micromat[28][24] = 9'b101101101;
assign micromat[28][25] = 9'b101101101;
assign micromat[28][26] = 9'b101101101;
assign micromat[28][27] = 9'b101101101;
assign micromat[28][28] = 9'b101101101;
assign micromat[28][29] = 9'b101101101;
assign micromat[28][30] = 9'b101101101;
assign micromat[28][31] = 9'b101101101;
assign micromat[28][32] = 9'b101101101;
assign micromat[28][33] = 9'b101101101;
assign micromat[28][34] = 9'b101101101;
assign micromat[28][35] = 9'b101101101;
assign micromat[28][36] = 9'b101101101;
assign micromat[28][37] = 9'b101101101;
assign micromat[28][38] = 9'b101101101;
assign micromat[28][39] = 9'b101101101;
assign micromat[28][40] = 9'b101101101;
assign micromat[28][41] = 9'b101101101;
assign micromat[28][42] = 9'b101101101;
assign micromat[28][43] = 9'b101101101;
assign micromat[28][44] = 9'b101101101;
assign micromat[28][45] = 9'b101101101;
assign micromat[28][46] = 9'b101101101;
assign micromat[28][47] = 9'b101101101;
assign micromat[28][48] = 9'b101101101;
assign micromat[28][49] = 9'b101101101;
assign micromat[28][50] = 9'b101101101;
assign micromat[28][51] = 9'b101101101;
assign micromat[28][52] = 9'b101101101;
assign micromat[28][53] = 9'b101101101;
assign micromat[28][54] = 9'b101101101;
assign micromat[28][55] = 9'b101101101;
assign micromat[28][56] = 9'b101101101;
assign micromat[28][57] = 9'b101101101;
assign micromat[28][58] = 9'b101101101;
assign micromat[28][59] = 9'b101101101;
assign micromat[28][60] = 9'b101101101;
assign micromat[28][61] = 9'b101101101;
assign micromat[28][62] = 9'b101101101;
assign micromat[28][63] = 9'b101101101;
assign micromat[28][64] = 9'b101101101;
assign micromat[28][65] = 9'b101101101;
assign micromat[28][66] = 9'b101101101;
assign micromat[28][67] = 9'b101101101;
assign micromat[28][68] = 9'b101101101;
assign micromat[28][69] = 9'b101101101;
assign micromat[28][70] = 9'b101101101;
assign micromat[28][71] = 9'b101101101;
assign micromat[28][72] = 9'b101101101;
assign micromat[28][73] = 9'b101101101;
assign micromat[28][74] = 9'b101101101;
assign micromat[28][75] = 9'b101101101;
assign micromat[28][76] = 9'b101101101;
assign micromat[28][77] = 9'b101101101;
assign micromat[28][78] = 9'b101101101;
assign micromat[28][79] = 9'b101101101;
assign micromat[28][80] = 9'b101101101;
assign micromat[28][81] = 9'b101101101;
assign micromat[28][82] = 9'b101101101;
assign micromat[28][83] = 9'b110110110;
assign micromat[28][84] = 9'b111111111;
assign micromat[28][85] = 9'b111111111;
assign micromat[28][86] = 9'b111111111;
assign micromat[28][87] = 9'b111111111;
assign micromat[28][88] = 9'b111111111;
assign micromat[28][89] = 9'b111111111;
assign micromat[28][90] = 9'b111111111;
assign micromat[28][91] = 9'b111111111;
assign micromat[28][92] = 9'b111111111;
assign micromat[28][93] = 9'b111111111;
assign micromat[28][94] = 9'b111111111;
assign micromat[28][95] = 9'b111111111;
assign micromat[28][96] = 9'b111111111;
assign micromat[28][97] = 9'b111111111;
assign micromat[28][98] = 9'b111111111;
assign micromat[28][99] = 9'b111111111;
assign micromat[29][0] = 9'b111111111;
assign micromat[29][1] = 9'b111111111;
assign micromat[29][2] = 9'b111111111;
assign micromat[29][3] = 9'b111111111;
assign micromat[29][4] = 9'b111111111;
assign micromat[29][5] = 9'b111111111;
assign micromat[29][6] = 9'b111111111;
assign micromat[29][7] = 9'b111111111;
assign micromat[29][8] = 9'b111111111;
assign micromat[29][9] = 9'b111111111;
assign micromat[29][10] = 9'b111111111;
assign micromat[29][11] = 9'b111111111;
assign micromat[29][12] = 9'b111111111;
assign micromat[29][13] = 9'b111111111;
assign micromat[29][14] = 9'b111111111;
assign micromat[29][15] = 9'b111111111;
assign micromat[29][16] = 9'b101101101;
assign micromat[29][17] = 9'b100000000;
assign micromat[29][18] = 9'b100000000;
assign micromat[29][19] = 9'b100000000;
assign micromat[29][20] = 9'b100000000;
assign micromat[29][21] = 9'b100000000;
assign micromat[29][22] = 9'b100000000;
assign micromat[29][23] = 9'b100000000;
assign micromat[29][24] = 9'b100000000;
assign micromat[29][25] = 9'b100000000;
assign micromat[29][26] = 9'b100000000;
assign micromat[29][27] = 9'b100000000;
assign micromat[29][28] = 9'b100000000;
assign micromat[29][29] = 9'b100000000;
assign micromat[29][30] = 9'b100000000;
assign micromat[29][31] = 9'b100000000;
assign micromat[29][32] = 9'b100000000;
assign micromat[29][33] = 9'b100000000;
assign micromat[29][34] = 9'b100000000;
assign micromat[29][35] = 9'b100000000;
assign micromat[29][36] = 9'b100000000;
assign micromat[29][37] = 9'b100000000;
assign micromat[29][38] = 9'b100000000;
assign micromat[29][39] = 9'b100000000;
assign micromat[29][40] = 9'b100000000;
assign micromat[29][41] = 9'b100000000;
assign micromat[29][42] = 9'b100000000;
assign micromat[29][43] = 9'b100000000;
assign micromat[29][44] = 9'b100000000;
assign micromat[29][45] = 9'b100000000;
assign micromat[29][46] = 9'b100000000;
assign micromat[29][47] = 9'b100000000;
assign micromat[29][48] = 9'b100000000;
assign micromat[29][49] = 9'b100000000;
assign micromat[29][50] = 9'b100000000;
assign micromat[29][51] = 9'b100000000;
assign micromat[29][52] = 9'b100000000;
assign micromat[29][53] = 9'b100000000;
assign micromat[29][54] = 9'b100000000;
assign micromat[29][55] = 9'b100000000;
assign micromat[29][56] = 9'b100000000;
assign micromat[29][57] = 9'b100000000;
assign micromat[29][58] = 9'b100000000;
assign micromat[29][59] = 9'b100000000;
assign micromat[29][60] = 9'b100000000;
assign micromat[29][61] = 9'b100000000;
assign micromat[29][62] = 9'b100000000;
assign micromat[29][63] = 9'b100000000;
assign micromat[29][64] = 9'b100000000;
assign micromat[29][65] = 9'b100000000;
assign micromat[29][66] = 9'b100000000;
assign micromat[29][67] = 9'b100000000;
assign micromat[29][68] = 9'b100000000;
assign micromat[29][69] = 9'b100000000;
assign micromat[29][70] = 9'b100000000;
assign micromat[29][71] = 9'b100000000;
assign micromat[29][72] = 9'b100000000;
assign micromat[29][73] = 9'b100000000;
assign micromat[29][74] = 9'b100000000;
assign micromat[29][75] = 9'b100000000;
assign micromat[29][76] = 9'b100000000;
assign micromat[29][77] = 9'b100000000;
assign micromat[29][78] = 9'b100000000;
assign micromat[29][79] = 9'b100000000;
assign micromat[29][80] = 9'b100000000;
assign micromat[29][81] = 9'b100000000;
assign micromat[29][82] = 9'b100000000;
assign micromat[29][83] = 9'b101101101;
assign micromat[29][84] = 9'b111111111;
assign micromat[29][85] = 9'b111111111;
assign micromat[29][86] = 9'b111111111;
assign micromat[29][87] = 9'b111111111;
assign micromat[29][88] = 9'b111111111;
assign micromat[29][89] = 9'b111111111;
assign micromat[29][90] = 9'b111111111;
assign micromat[29][91] = 9'b111111111;
assign micromat[29][92] = 9'b111111111;
assign micromat[29][93] = 9'b111111111;
assign micromat[29][94] = 9'b111111111;
assign micromat[29][95] = 9'b111111111;
assign micromat[29][96] = 9'b111111111;
assign micromat[29][97] = 9'b111111111;
assign micromat[29][98] = 9'b111111111;
assign micromat[29][99] = 9'b111111111;
assign micromat[30][0] = 9'b111111111;
assign micromat[30][1] = 9'b111111111;
assign micromat[30][2] = 9'b111111111;
assign micromat[30][3] = 9'b111111111;
assign micromat[30][4] = 9'b111111111;
assign micromat[30][5] = 9'b111111111;
assign micromat[30][6] = 9'b111111111;
assign micromat[30][7] = 9'b111111111;
assign micromat[30][8] = 9'b111111111;
assign micromat[30][9] = 9'b111111111;
assign micromat[30][10] = 9'b111111111;
assign micromat[30][11] = 9'b111111111;
assign micromat[30][12] = 9'b111111111;
assign micromat[30][13] = 9'b111111111;
assign micromat[30][14] = 9'b111111111;
assign micromat[30][15] = 9'b111111111;
assign micromat[30][16] = 9'b101101101;
assign micromat[30][17] = 9'b100100100;
assign micromat[30][18] = 9'b100100100;
assign micromat[30][19] = 9'b100100100;
assign micromat[30][20] = 9'b100100100;
assign micromat[30][21] = 9'b100100100;
assign micromat[30][22] = 9'b100100100;
assign micromat[30][23] = 9'b100100100;
assign micromat[30][24] = 9'b100100100;
assign micromat[30][25] = 9'b100100100;
assign micromat[30][26] = 9'b100100100;
assign micromat[30][27] = 9'b100100100;
assign micromat[30][28] = 9'b100100100;
assign micromat[30][29] = 9'b100100100;
assign micromat[30][30] = 9'b100100100;
assign micromat[30][31] = 9'b100100100;
assign micromat[30][32] = 9'b100100100;
assign micromat[30][33] = 9'b100100100;
assign micromat[30][34] = 9'b100100100;
assign micromat[30][35] = 9'b100100100;
assign micromat[30][36] = 9'b100100100;
assign micromat[30][37] = 9'b100100100;
assign micromat[30][38] = 9'b100100100;
assign micromat[30][39] = 9'b100100100;
assign micromat[30][40] = 9'b100100100;
assign micromat[30][41] = 9'b100100100;
assign micromat[30][42] = 9'b100100100;
assign micromat[30][43] = 9'b100100100;
assign micromat[30][44] = 9'b100100100;
assign micromat[30][45] = 9'b100100100;
assign micromat[30][46] = 9'b100100100;
assign micromat[30][47] = 9'b100100100;
assign micromat[30][48] = 9'b100100100;
assign micromat[30][49] = 9'b100100100;
assign micromat[30][50] = 9'b100100100;
assign micromat[30][51] = 9'b100100100;
assign micromat[30][52] = 9'b100100100;
assign micromat[30][53] = 9'b100100100;
assign micromat[30][54] = 9'b100100100;
assign micromat[30][55] = 9'b100100100;
assign micromat[30][56] = 9'b100100100;
assign micromat[30][57] = 9'b100100100;
assign micromat[30][58] = 9'b100100100;
assign micromat[30][59] = 9'b100100100;
assign micromat[30][60] = 9'b100100100;
assign micromat[30][61] = 9'b100100100;
assign micromat[30][62] = 9'b100100100;
assign micromat[30][63] = 9'b100100100;
assign micromat[30][64] = 9'b100100100;
assign micromat[30][65] = 9'b100100100;
assign micromat[30][66] = 9'b100000000;
assign micromat[30][67] = 9'b100000000;
assign micromat[30][68] = 9'b100000000;
assign micromat[30][69] = 9'b100100100;
assign micromat[30][70] = 9'b100100100;
assign micromat[30][71] = 9'b100100100;
assign micromat[30][72] = 9'b100100100;
assign micromat[30][73] = 9'b100100100;
assign micromat[30][74] = 9'b100100100;
assign micromat[30][75] = 9'b100100100;
assign micromat[30][76] = 9'b100100100;
assign micromat[30][77] = 9'b100100100;
assign micromat[30][78] = 9'b100100100;
assign micromat[30][79] = 9'b100100100;
assign micromat[30][80] = 9'b100100100;
assign micromat[30][81] = 9'b100100100;
assign micromat[30][82] = 9'b100100100;
assign micromat[30][83] = 9'b101101101;
assign micromat[30][84] = 9'b111111111;
assign micromat[30][85] = 9'b111111111;
assign micromat[30][86] = 9'b111111111;
assign micromat[30][87] = 9'b111111111;
assign micromat[30][88] = 9'b111111111;
assign micromat[30][89] = 9'b111111111;
assign micromat[30][90] = 9'b111111111;
assign micromat[30][91] = 9'b111111111;
assign micromat[30][92] = 9'b111111111;
assign micromat[30][93] = 9'b111111111;
assign micromat[30][94] = 9'b111111111;
assign micromat[30][95] = 9'b111111111;
assign micromat[30][96] = 9'b111111111;
assign micromat[30][97] = 9'b111111111;
assign micromat[30][98] = 9'b111111111;
assign micromat[30][99] = 9'b111111111;
assign micromat[31][0] = 9'b111111111;
assign micromat[31][1] = 9'b111111111;
assign micromat[31][2] = 9'b111111111;
assign micromat[31][3] = 9'b111111111;
assign micromat[31][4] = 9'b111111111;
assign micromat[31][5] = 9'b111111111;
assign micromat[31][6] = 9'b111111111;
assign micromat[31][7] = 9'b111111111;
assign micromat[31][8] = 9'b111111111;
assign micromat[31][9] = 9'b111111111;
assign micromat[31][10] = 9'b111111111;
assign micromat[31][11] = 9'b111111111;
assign micromat[31][12] = 9'b111111111;
assign micromat[31][13] = 9'b111111111;
assign micromat[31][14] = 9'b100100100;
assign micromat[31][15] = 9'b100000000;
assign micromat[31][16] = 9'b101101101;
assign micromat[31][17] = 9'b111111111;
assign micromat[31][18] = 9'b111111111;
assign micromat[31][19] = 9'b111111111;
assign micromat[31][20] = 9'b111111111;
assign micromat[31][21] = 9'b111111111;
assign micromat[31][22] = 9'b111111111;
assign micromat[31][23] = 9'b111111111;
assign micromat[31][24] = 9'b111111111;
assign micromat[31][25] = 9'b111111111;
assign micromat[31][26] = 9'b111111111;
assign micromat[31][27] = 9'b111111111;
assign micromat[31][28] = 9'b111111111;
assign micromat[31][29] = 9'b111111111;
assign micromat[31][30] = 9'b111111111;
assign micromat[31][31] = 9'b111111111;
assign micromat[31][32] = 9'b111111111;
assign micromat[31][33] = 9'b111111111;
assign micromat[31][34] = 9'b111111111;
assign micromat[31][35] = 9'b111111111;
assign micromat[31][36] = 9'b111111111;
assign micromat[31][37] = 9'b111111111;
assign micromat[31][38] = 9'b111111111;
assign micromat[31][39] = 9'b111111111;
assign micromat[31][40] = 9'b111111111;
assign micromat[31][41] = 9'b111111111;
assign micromat[31][42] = 9'b111111111;
assign micromat[31][43] = 9'b111111111;
assign micromat[31][44] = 9'b111111111;
assign micromat[31][45] = 9'b111111111;
assign micromat[31][46] = 9'b111111111;
assign micromat[31][47] = 9'b111111111;
assign micromat[31][48] = 9'b111111111;
assign micromat[31][49] = 9'b111111111;
assign micromat[31][50] = 9'b111111111;
assign micromat[31][51] = 9'b111111111;
assign micromat[31][52] = 9'b111111111;
assign micromat[31][53] = 9'b111111111;
assign micromat[31][54] = 9'b111111111;
assign micromat[31][55] = 9'b111111111;
assign micromat[31][56] = 9'b111111111;
assign micromat[31][57] = 9'b111111111;
assign micromat[31][58] = 9'b111111111;
assign micromat[31][59] = 9'b111111111;
assign micromat[31][60] = 9'b111111111;
assign micromat[31][61] = 9'b111111111;
assign micromat[31][62] = 9'b111111111;
assign micromat[31][63] = 9'b111111111;
assign micromat[31][64] = 9'b111111111;
assign micromat[31][65] = 9'b111111111;
assign micromat[31][66] = 9'b110010010;
assign micromat[31][67] = 9'b100000000;
assign micromat[31][68] = 9'b100000000;
assign micromat[31][69] = 9'b111111111;
assign micromat[31][70] = 9'b111111111;
assign micromat[31][71] = 9'b111111111;
assign micromat[31][72] = 9'b111111111;
assign micromat[31][73] = 9'b111111111;
assign micromat[31][74] = 9'b111111111;
assign micromat[31][75] = 9'b111111111;
assign micromat[31][76] = 9'b111111111;
assign micromat[31][77] = 9'b111111111;
assign micromat[31][78] = 9'b111111111;
assign micromat[31][79] = 9'b111111111;
assign micromat[31][80] = 9'b111111111;
assign micromat[31][81] = 9'b111111111;
assign micromat[31][82] = 9'b111111111;
assign micromat[31][83] = 9'b101001101;
assign micromat[31][84] = 9'b100000000;
assign micromat[31][85] = 9'b100100100;
assign micromat[31][86] = 9'b111111111;
assign micromat[31][87] = 9'b111111111;
assign micromat[31][88] = 9'b111111111;
assign micromat[31][89] = 9'b111111111;
assign micromat[31][90] = 9'b111111111;
assign micromat[31][91] = 9'b111111111;
assign micromat[31][92] = 9'b111111111;
assign micromat[31][93] = 9'b111111111;
assign micromat[31][94] = 9'b111111111;
assign micromat[31][95] = 9'b111111111;
assign micromat[31][96] = 9'b111111111;
assign micromat[31][97] = 9'b111111111;
assign micromat[31][98] = 9'b111111111;
assign micromat[31][99] = 9'b111111111;
assign micromat[32][0] = 9'b111111111;
assign micromat[32][1] = 9'b111111111;
assign micromat[32][2] = 9'b111111111;
assign micromat[32][3] = 9'b111111111;
assign micromat[32][4] = 9'b111111111;
assign micromat[32][5] = 9'b111111111;
assign micromat[32][6] = 9'b111111111;
assign micromat[32][7] = 9'b111111111;
assign micromat[32][8] = 9'b111111111;
assign micromat[32][9] = 9'b111111111;
assign micromat[32][10] = 9'b111111111;
assign micromat[32][11] = 9'b111111111;
assign micromat[32][12] = 9'b111111111;
assign micromat[32][13] = 9'b111111111;
assign micromat[32][14] = 9'b100100100;
assign micromat[32][15] = 9'b100000000;
assign micromat[32][16] = 9'b101101101;
assign micromat[32][17] = 9'b111111111;
assign micromat[32][18] = 9'b111111111;
assign micromat[32][19] = 9'b111111111;
assign micromat[32][20] = 9'b111111111;
assign micromat[32][21] = 9'b111111111;
assign micromat[32][22] = 9'b111111111;
assign micromat[32][23] = 9'b111111111;
assign micromat[32][24] = 9'b111111111;
assign micromat[32][25] = 9'b111111111;
assign micromat[32][26] = 9'b111111111;
assign micromat[32][27] = 9'b111111111;
assign micromat[32][28] = 9'b111111111;
assign micromat[32][29] = 9'b111111111;
assign micromat[32][30] = 9'b111111111;
assign micromat[32][31] = 9'b111111111;
assign micromat[32][32] = 9'b111111111;
assign micromat[32][33] = 9'b111111111;
assign micromat[32][34] = 9'b111111111;
assign micromat[32][35] = 9'b111111111;
assign micromat[32][36] = 9'b111111111;
assign micromat[32][37] = 9'b111111111;
assign micromat[32][38] = 9'b111111111;
assign micromat[32][39] = 9'b111111111;
assign micromat[32][40] = 9'b111111111;
assign micromat[32][41] = 9'b111111111;
assign micromat[32][42] = 9'b111111111;
assign micromat[32][43] = 9'b111111111;
assign micromat[32][44] = 9'b111111111;
assign micromat[32][45] = 9'b111111111;
assign micromat[32][46] = 9'b111111111;
assign micromat[32][47] = 9'b111111111;
assign micromat[32][48] = 9'b111111111;
assign micromat[32][49] = 9'b111111111;
assign micromat[32][50] = 9'b111111111;
assign micromat[32][51] = 9'b111111111;
assign micromat[32][52] = 9'b111111111;
assign micromat[32][53] = 9'b111111111;
assign micromat[32][54] = 9'b111111111;
assign micromat[32][55] = 9'b111111111;
assign micromat[32][56] = 9'b111111111;
assign micromat[32][57] = 9'b111111111;
assign micromat[32][58] = 9'b111111111;
assign micromat[32][59] = 9'b111111111;
assign micromat[32][60] = 9'b111111111;
assign micromat[32][61] = 9'b111111111;
assign micromat[32][62] = 9'b111111111;
assign micromat[32][63] = 9'b111111111;
assign micromat[32][64] = 9'b111111111;
assign micromat[32][65] = 9'b111111111;
assign micromat[32][66] = 9'b110010010;
assign micromat[32][67] = 9'b100000000;
assign micromat[32][68] = 9'b100000000;
assign micromat[32][69] = 9'b111111111;
assign micromat[32][70] = 9'b111111111;
assign micromat[32][71] = 9'b111111111;
assign micromat[32][72] = 9'b111111111;
assign micromat[32][73] = 9'b111111111;
assign micromat[32][74] = 9'b111111111;
assign micromat[32][75] = 9'b111111111;
assign micromat[32][76] = 9'b111111111;
assign micromat[32][77] = 9'b111111111;
assign micromat[32][78] = 9'b111111111;
assign micromat[32][79] = 9'b111111111;
assign micromat[32][80] = 9'b111111111;
assign micromat[32][81] = 9'b111111111;
assign micromat[32][82] = 9'b111111111;
assign micromat[32][83] = 9'b101001101;
assign micromat[32][84] = 9'b100000000;
assign micromat[32][85] = 9'b100100100;
assign micromat[32][86] = 9'b111111111;
assign micromat[32][87] = 9'b111111111;
assign micromat[32][88] = 9'b111111111;
assign micromat[32][89] = 9'b111111111;
assign micromat[32][90] = 9'b111111111;
assign micromat[32][91] = 9'b111111111;
assign micromat[32][92] = 9'b111111111;
assign micromat[32][93] = 9'b111111111;
assign micromat[32][94] = 9'b111111111;
assign micromat[32][95] = 9'b111111111;
assign micromat[32][96] = 9'b111111111;
assign micromat[32][97] = 9'b111111111;
assign micromat[32][98] = 9'b111111111;
assign micromat[32][99] = 9'b111111111;
assign micromat[33][0] = 9'b111111111;
assign micromat[33][1] = 9'b111111111;
assign micromat[33][2] = 9'b111111111;
assign micromat[33][3] = 9'b111111111;
assign micromat[33][4] = 9'b111111111;
assign micromat[33][5] = 9'b111111111;
assign micromat[33][6] = 9'b111111111;
assign micromat[33][7] = 9'b111111111;
assign micromat[33][8] = 9'b111111111;
assign micromat[33][9] = 9'b111111111;
assign micromat[33][10] = 9'b111111111;
assign micromat[33][11] = 9'b111111111;
assign micromat[33][12] = 9'b111111111;
assign micromat[33][13] = 9'b111111111;
assign micromat[33][14] = 9'b100100100;
assign micromat[33][15] = 9'b100000000;
assign micromat[33][16] = 9'b101101101;
assign micromat[33][17] = 9'b111111111;
assign micromat[33][18] = 9'b111111111;
assign micromat[33][19] = 9'b111111111;
assign micromat[33][20] = 9'b111111111;
assign micromat[33][21] = 9'b111111111;
assign micromat[33][22] = 9'b111111111;
assign micromat[33][23] = 9'b111111111;
assign micromat[33][24] = 9'b111111111;
assign micromat[33][25] = 9'b111111111;
assign micromat[33][26] = 9'b111111111;
assign micromat[33][27] = 9'b111111111;
assign micromat[33][28] = 9'b111111111;
assign micromat[33][29] = 9'b111111111;
assign micromat[33][30] = 9'b111111111;
assign micromat[33][31] = 9'b111111111;
assign micromat[33][32] = 9'b111111111;
assign micromat[33][33] = 9'b111111111;
assign micromat[33][34] = 9'b111111111;
assign micromat[33][35] = 9'b111111111;
assign micromat[33][36] = 9'b111111111;
assign micromat[33][37] = 9'b111111111;
assign micromat[33][38] = 9'b111111111;
assign micromat[33][39] = 9'b111111111;
assign micromat[33][40] = 9'b111111111;
assign micromat[33][41] = 9'b111111111;
assign micromat[33][42] = 9'b111111111;
assign micromat[33][43] = 9'b111111111;
assign micromat[33][44] = 9'b111111111;
assign micromat[33][45] = 9'b111111111;
assign micromat[33][46] = 9'b111111111;
assign micromat[33][47] = 9'b111111111;
assign micromat[33][48] = 9'b111111111;
assign micromat[33][49] = 9'b111111111;
assign micromat[33][50] = 9'b111111111;
assign micromat[33][51] = 9'b111111111;
assign micromat[33][52] = 9'b111111111;
assign micromat[33][53] = 9'b111111111;
assign micromat[33][54] = 9'b111111111;
assign micromat[33][55] = 9'b111111111;
assign micromat[33][56] = 9'b111111111;
assign micromat[33][57] = 9'b111111111;
assign micromat[33][58] = 9'b111111111;
assign micromat[33][59] = 9'b111111111;
assign micromat[33][60] = 9'b111111111;
assign micromat[33][61] = 9'b111111111;
assign micromat[33][62] = 9'b111111111;
assign micromat[33][63] = 9'b111111111;
assign micromat[33][64] = 9'b110111111;
assign micromat[33][65] = 9'b110111111;
assign micromat[33][66] = 9'b101110001;
assign micromat[33][67] = 9'b100000000;
assign micromat[33][68] = 9'b100000000;
assign micromat[33][69] = 9'b111111111;
assign micromat[33][70] = 9'b111111111;
assign micromat[33][71] = 9'b111111111;
assign micromat[33][72] = 9'b111111111;
assign micromat[33][73] = 9'b110111111;
assign micromat[33][74] = 9'b101001001;
assign micromat[33][75] = 9'b101001000;
assign micromat[33][76] = 9'b101001000;
assign micromat[33][77] = 9'b100101000;
assign micromat[33][78] = 9'b101101101;
assign micromat[33][79] = 9'b111111111;
assign micromat[33][80] = 9'b111111111;
assign micromat[33][81] = 9'b110110111;
assign micromat[33][82] = 9'b111111111;
assign micromat[33][83] = 9'b101001001;
assign micromat[33][84] = 9'b100000000;
assign micromat[33][85] = 9'b100100100;
assign micromat[33][86] = 9'b111111111;
assign micromat[33][87] = 9'b111111111;
assign micromat[33][88] = 9'b111111111;
assign micromat[33][89] = 9'b111111111;
assign micromat[33][90] = 9'b111111111;
assign micromat[33][91] = 9'b111111111;
assign micromat[33][92] = 9'b111111111;
assign micromat[33][93] = 9'b111111111;
assign micromat[33][94] = 9'b111111111;
assign micromat[33][95] = 9'b111111111;
assign micromat[33][96] = 9'b111111111;
assign micromat[33][97] = 9'b111111111;
assign micromat[33][98] = 9'b111111111;
assign micromat[33][99] = 9'b111111111;
assign micromat[34][0] = 9'b111111111;
assign micromat[34][1] = 9'b111111111;
assign micromat[34][2] = 9'b111111111;
assign micromat[34][3] = 9'b111111111;
assign micromat[34][4] = 9'b111111111;
assign micromat[34][5] = 9'b111111111;
assign micromat[34][6] = 9'b111111111;
assign micromat[34][7] = 9'b111111111;
assign micromat[34][8] = 9'b111111111;
assign micromat[34][9] = 9'b111111111;
assign micromat[34][10] = 9'b111111111;
assign micromat[34][11] = 9'b111111111;
assign micromat[34][12] = 9'b111111111;
assign micromat[34][13] = 9'b111111111;
assign micromat[34][14] = 9'b100100100;
assign micromat[34][15] = 9'b100000000;
assign micromat[34][16] = 9'b101101101;
assign micromat[34][17] = 9'b111111111;
assign micromat[34][18] = 9'b111111111;
assign micromat[34][19] = 9'b111111111;
assign micromat[34][20] = 9'b111111111;
assign micromat[34][21] = 9'b111111111;
assign micromat[34][22] = 9'b111111111;
assign micromat[34][23] = 9'b111111111;
assign micromat[34][24] = 9'b111111111;
assign micromat[34][25] = 9'b111111111;
assign micromat[34][26] = 9'b111111111;
assign micromat[34][27] = 9'b111111111;
assign micromat[34][28] = 9'b111111111;
assign micromat[34][29] = 9'b111111111;
assign micromat[34][30] = 9'b111111111;
assign micromat[34][31] = 9'b111111111;
assign micromat[34][32] = 9'b111111111;
assign micromat[34][33] = 9'b111111111;
assign micromat[34][34] = 9'b111111111;
assign micromat[34][35] = 9'b111111111;
assign micromat[34][36] = 9'b111111111;
assign micromat[34][37] = 9'b111111111;
assign micromat[34][38] = 9'b111111111;
assign micromat[34][39] = 9'b111111111;
assign micromat[34][40] = 9'b111111111;
assign micromat[34][41] = 9'b111111111;
assign micromat[34][42] = 9'b111111111;
assign micromat[34][43] = 9'b111111111;
assign micromat[34][44] = 9'b111111111;
assign micromat[34][45] = 9'b111111111;
assign micromat[34][46] = 9'b111111111;
assign micromat[34][47] = 9'b111111111;
assign micromat[34][48] = 9'b111111111;
assign micromat[34][49] = 9'b111111111;
assign micromat[34][50] = 9'b111111111;
assign micromat[34][51] = 9'b111111111;
assign micromat[34][52] = 9'b111111111;
assign micromat[34][53] = 9'b111111111;
assign micromat[34][54] = 9'b111111111;
assign micromat[34][55] = 9'b111111111;
assign micromat[34][56] = 9'b111111111;
assign micromat[34][57] = 9'b111111111;
assign micromat[34][58] = 9'b111111111;
assign micromat[34][59] = 9'b111111111;
assign micromat[34][60] = 9'b111111111;
assign micromat[34][61] = 9'b111111111;
assign micromat[34][62] = 9'b111111111;
assign micromat[34][63] = 9'b111111111;
assign micromat[34][64] = 9'b110110111;
assign micromat[34][65] = 9'b110110111;
assign micromat[34][66] = 9'b101101101;
assign micromat[34][67] = 9'b100000000;
assign micromat[34][68] = 9'b100000000;
assign micromat[34][69] = 9'b111111111;
assign micromat[34][70] = 9'b111111111;
assign micromat[34][71] = 9'b111111111;
assign micromat[34][72] = 9'b111111111;
assign micromat[34][73] = 9'b110111111;
assign micromat[34][74] = 9'b100000000;
assign micromat[34][75] = 9'b100000000;
assign micromat[34][76] = 9'b100000000;
assign micromat[34][77] = 9'b100000000;
assign micromat[34][78] = 9'b100100100;
assign micromat[34][79] = 9'b111111111;
assign micromat[34][80] = 9'b111111111;
assign micromat[34][81] = 9'b110110111;
assign micromat[34][82] = 9'b110111111;
assign micromat[34][83] = 9'b101001001;
assign micromat[34][84] = 9'b100000000;
assign micromat[34][85] = 9'b100100100;
assign micromat[34][86] = 9'b111111111;
assign micromat[34][87] = 9'b111111111;
assign micromat[34][88] = 9'b111111111;
assign micromat[34][89] = 9'b111111111;
assign micromat[34][90] = 9'b111111111;
assign micromat[34][91] = 9'b111111111;
assign micromat[34][92] = 9'b111111111;
assign micromat[34][93] = 9'b111111111;
assign micromat[34][94] = 9'b111111111;
assign micromat[34][95] = 9'b111111111;
assign micromat[34][96] = 9'b111111111;
assign micromat[34][97] = 9'b111111111;
assign micromat[34][98] = 9'b111111111;
assign micromat[34][99] = 9'b111111111;
assign micromat[35][0] = 9'b111111111;
assign micromat[35][1] = 9'b111111111;
assign micromat[35][2] = 9'b111111111;
assign micromat[35][3] = 9'b111111111;
assign micromat[35][4] = 9'b111111111;
assign micromat[35][5] = 9'b111111111;
assign micromat[35][6] = 9'b111111111;
assign micromat[35][7] = 9'b111111111;
assign micromat[35][8] = 9'b111111111;
assign micromat[35][9] = 9'b111111111;
assign micromat[35][10] = 9'b111111111;
assign micromat[35][11] = 9'b111111111;
assign micromat[35][12] = 9'b111111111;
assign micromat[35][13] = 9'b111111111;
assign micromat[35][14] = 9'b100100100;
assign micromat[35][15] = 9'b100000000;
assign micromat[35][16] = 9'b101101101;
assign micromat[35][17] = 9'b111111111;
assign micromat[35][18] = 9'b111111111;
assign micromat[35][19] = 9'b111111111;
assign micromat[35][20] = 9'b111111111;
assign micromat[35][21] = 9'b110010010;
assign micromat[35][22] = 9'b101101101;
assign micromat[35][23] = 9'b101110001;
assign micromat[35][24] = 9'b101110001;
assign micromat[35][25] = 9'b101110001;
assign micromat[35][26] = 9'b101110001;
assign micromat[35][27] = 9'b101110001;
assign micromat[35][28] = 9'b101110001;
assign micromat[35][29] = 9'b101110001;
assign micromat[35][30] = 9'b101110001;
assign micromat[35][31] = 9'b101110001;
assign micromat[35][32] = 9'b101110001;
assign micromat[35][33] = 9'b101110001;
assign micromat[35][34] = 9'b101110001;
assign micromat[35][35] = 9'b101110001;
assign micromat[35][36] = 9'b101110001;
assign micromat[35][37] = 9'b101110001;
assign micromat[35][38] = 9'b101110001;
assign micromat[35][39] = 9'b101110001;
assign micromat[35][40] = 9'b101110001;
assign micromat[35][41] = 9'b101110001;
assign micromat[35][42] = 9'b101110001;
assign micromat[35][43] = 9'b101110001;
assign micromat[35][44] = 9'b101110001;
assign micromat[35][45] = 9'b101110001;
assign micromat[35][46] = 9'b101110001;
assign micromat[35][47] = 9'b101110001;
assign micromat[35][48] = 9'b101110001;
assign micromat[35][49] = 9'b101110001;
assign micromat[35][50] = 9'b101110001;
assign micromat[35][51] = 9'b101110001;
assign micromat[35][52] = 9'b101110001;
assign micromat[35][53] = 9'b101110001;
assign micromat[35][54] = 9'b101110001;
assign micromat[35][55] = 9'b101110001;
assign micromat[35][56] = 9'b101110001;
assign micromat[35][57] = 9'b101110001;
assign micromat[35][58] = 9'b101110001;
assign micromat[35][59] = 9'b101110001;
assign micromat[35][60] = 9'b101110001;
assign micromat[35][61] = 9'b110010001;
assign micromat[35][62] = 9'b111111111;
assign micromat[35][63] = 9'b111111111;
assign micromat[35][64] = 9'b110110111;
assign micromat[35][65] = 9'b110110111;
assign micromat[35][66] = 9'b101101101;
assign micromat[35][67] = 9'b100000000;
assign micromat[35][68] = 9'b100000000;
assign micromat[35][69] = 9'b111111111;
assign micromat[35][70] = 9'b111111111;
assign micromat[35][71] = 9'b110110111;
assign micromat[35][72] = 9'b101101101;
assign micromat[35][73] = 9'b101101101;
assign micromat[35][74] = 9'b101001001;
assign micromat[35][75] = 9'b101001001;
assign micromat[35][76] = 9'b101001001;
assign micromat[35][77] = 9'b101001001;
assign micromat[35][78] = 9'b101001001;
assign micromat[35][79] = 9'b101110001;
assign micromat[35][80] = 9'b101110001;
assign micromat[35][81] = 9'b110010110;
assign micromat[35][82] = 9'b110111111;
assign micromat[35][83] = 9'b101001001;
assign micromat[35][84] = 9'b100000000;
assign micromat[35][85] = 9'b100100100;
assign micromat[35][86] = 9'b111111111;
assign micromat[35][87] = 9'b111111111;
assign micromat[35][88] = 9'b111111111;
assign micromat[35][89] = 9'b111111111;
assign micromat[35][90] = 9'b111111111;
assign micromat[35][91] = 9'b111111111;
assign micromat[35][92] = 9'b111111111;
assign micromat[35][93] = 9'b111111111;
assign micromat[35][94] = 9'b111111111;
assign micromat[35][95] = 9'b111111111;
assign micromat[35][96] = 9'b111111111;
assign micromat[35][97] = 9'b111111111;
assign micromat[35][98] = 9'b111111111;
assign micromat[35][99] = 9'b111111111;
assign micromat[36][0] = 9'b111111111;
assign micromat[36][1] = 9'b111111111;
assign micromat[36][2] = 9'b111111111;
assign micromat[36][3] = 9'b111111111;
assign micromat[36][4] = 9'b111111111;
assign micromat[36][5] = 9'b111111111;
assign micromat[36][6] = 9'b111111111;
assign micromat[36][7] = 9'b111111111;
assign micromat[36][8] = 9'b111111111;
assign micromat[36][9] = 9'b111111111;
assign micromat[36][10] = 9'b111111111;
assign micromat[36][11] = 9'b111111111;
assign micromat[36][12] = 9'b111111111;
assign micromat[36][13] = 9'b111111111;
assign micromat[36][14] = 9'b100100100;
assign micromat[36][15] = 9'b100000000;
assign micromat[36][16] = 9'b101101101;
assign micromat[36][17] = 9'b111111111;
assign micromat[36][18] = 9'b111111111;
assign micromat[36][19] = 9'b111111111;
assign micromat[36][20] = 9'b111111111;
assign micromat[36][21] = 9'b100100100;
assign micromat[36][22] = 9'b100000000;
assign micromat[36][23] = 9'b100000000;
assign micromat[36][24] = 9'b100000000;
assign micromat[36][25] = 9'b100000000;
assign micromat[36][26] = 9'b100000000;
assign micromat[36][27] = 9'b100000000;
assign micromat[36][28] = 9'b100000000;
assign micromat[36][29] = 9'b100000000;
assign micromat[36][30] = 9'b100000000;
assign micromat[36][31] = 9'b100000000;
assign micromat[36][32] = 9'b100000000;
assign micromat[36][33] = 9'b100000000;
assign micromat[36][34] = 9'b100000000;
assign micromat[36][35] = 9'b100000000;
assign micromat[36][36] = 9'b100000000;
assign micromat[36][37] = 9'b100000000;
assign micromat[36][38] = 9'b100000000;
assign micromat[36][39] = 9'b100000000;
assign micromat[36][40] = 9'b100000000;
assign micromat[36][41] = 9'b100000000;
assign micromat[36][42] = 9'b100000000;
assign micromat[36][43] = 9'b100000000;
assign micromat[36][44] = 9'b100000000;
assign micromat[36][45] = 9'b100000000;
assign micromat[36][46] = 9'b100000000;
assign micromat[36][47] = 9'b100000000;
assign micromat[36][48] = 9'b100000000;
assign micromat[36][49] = 9'b100000000;
assign micromat[36][50] = 9'b100000000;
assign micromat[36][51] = 9'b100000000;
assign micromat[36][52] = 9'b100000000;
assign micromat[36][53] = 9'b100000000;
assign micromat[36][54] = 9'b100000000;
assign micromat[36][55] = 9'b100000000;
assign micromat[36][56] = 9'b100000000;
assign micromat[36][57] = 9'b100000000;
assign micromat[36][58] = 9'b100000000;
assign micromat[36][59] = 9'b100000000;
assign micromat[36][60] = 9'b100000000;
assign micromat[36][61] = 9'b100000000;
assign micromat[36][62] = 9'b110111111;
assign micromat[36][63] = 9'b111111111;
assign micromat[36][64] = 9'b110110111;
assign micromat[36][65] = 9'b110110111;
assign micromat[36][66] = 9'b101101101;
assign micromat[36][67] = 9'b100000000;
assign micromat[36][68] = 9'b100000000;
assign micromat[36][69] = 9'b111111111;
assign micromat[36][70] = 9'b111111111;
assign micromat[36][71] = 9'b101101101;
assign micromat[36][72] = 9'b100000000;
assign micromat[36][73] = 9'b100000000;
assign micromat[36][74] = 9'b111111111;
assign micromat[36][75] = 9'b111111111;
assign micromat[36][76] = 9'b111111111;
assign micromat[36][77] = 9'b111111111;
assign micromat[36][78] = 9'b110010010;
assign micromat[36][79] = 9'b100000000;
assign micromat[36][80] = 9'b100000000;
assign micromat[36][81] = 9'b110010010;
assign micromat[36][82] = 9'b111111111;
assign micromat[36][83] = 9'b101001001;
assign micromat[36][84] = 9'b100000000;
assign micromat[36][85] = 9'b100100100;
assign micromat[36][86] = 9'b111111111;
assign micromat[36][87] = 9'b111111111;
assign micromat[36][88] = 9'b111111111;
assign micromat[36][89] = 9'b111111111;
assign micromat[36][90] = 9'b111111111;
assign micromat[36][91] = 9'b111111111;
assign micromat[36][92] = 9'b111111111;
assign micromat[36][93] = 9'b111111111;
assign micromat[36][94] = 9'b111111111;
assign micromat[36][95] = 9'b111111111;
assign micromat[36][96] = 9'b111111111;
assign micromat[36][97] = 9'b111111111;
assign micromat[36][98] = 9'b111111111;
assign micromat[36][99] = 9'b111111111;
assign micromat[37][0] = 9'b111111111;
assign micromat[37][1] = 9'b111111111;
assign micromat[37][2] = 9'b111111111;
assign micromat[37][3] = 9'b111111111;
assign micromat[37][4] = 9'b111111111;
assign micromat[37][5] = 9'b111111111;
assign micromat[37][6] = 9'b111111111;
assign micromat[37][7] = 9'b111111111;
assign micromat[37][8] = 9'b111111111;
assign micromat[37][9] = 9'b111111111;
assign micromat[37][10] = 9'b111111111;
assign micromat[37][11] = 9'b111111111;
assign micromat[37][12] = 9'b111111111;
assign micromat[37][13] = 9'b111111111;
assign micromat[37][14] = 9'b100100100;
assign micromat[37][15] = 9'b100000000;
assign micromat[37][16] = 9'b101101101;
assign micromat[37][17] = 9'b111111111;
assign micromat[37][18] = 9'b111111111;
assign micromat[37][19] = 9'b111111111;
assign micromat[37][20] = 9'b111111111;
assign micromat[37][21] = 9'b100101000;
assign micromat[37][22] = 9'b100000000;
assign micromat[37][23] = 9'b100000000;
assign micromat[37][24] = 9'b100000000;
assign micromat[37][25] = 9'b100000000;
assign micromat[37][26] = 9'b100000000;
assign micromat[37][27] = 9'b100000000;
assign micromat[37][28] = 9'b100000000;
assign micromat[37][29] = 9'b100000000;
assign micromat[37][30] = 9'b100000000;
assign micromat[37][31] = 9'b100000000;
assign micromat[37][32] = 9'b100000000;
assign micromat[37][33] = 9'b100000000;
assign micromat[37][34] = 9'b100000000;
assign micromat[37][35] = 9'b100000000;
assign micromat[37][36] = 9'b100000000;
assign micromat[37][37] = 9'b100000000;
assign micromat[37][38] = 9'b100000000;
assign micromat[37][39] = 9'b100000000;
assign micromat[37][40] = 9'b100000000;
assign micromat[37][41] = 9'b100000000;
assign micromat[37][42] = 9'b100000000;
assign micromat[37][43] = 9'b100000000;
assign micromat[37][44] = 9'b100000000;
assign micromat[37][45] = 9'b100000000;
assign micromat[37][46] = 9'b100000000;
assign micromat[37][47] = 9'b100000000;
assign micromat[37][48] = 9'b100000000;
assign micromat[37][49] = 9'b100000000;
assign micromat[37][50] = 9'b100000000;
assign micromat[37][51] = 9'b100000000;
assign micromat[37][52] = 9'b100000000;
assign micromat[37][53] = 9'b100000000;
assign micromat[37][54] = 9'b100000000;
assign micromat[37][55] = 9'b100000000;
assign micromat[37][56] = 9'b100000000;
assign micromat[37][57] = 9'b100000000;
assign micromat[37][58] = 9'b100000000;
assign micromat[37][59] = 9'b100000000;
assign micromat[37][60] = 9'b100000000;
assign micromat[37][61] = 9'b100000000;
assign micromat[37][62] = 9'b110111111;
assign micromat[37][63] = 9'b111111111;
assign micromat[37][64] = 9'b110110111;
assign micromat[37][65] = 9'b110110111;
assign micromat[37][66] = 9'b101101101;
assign micromat[37][67] = 9'b100000000;
assign micromat[37][68] = 9'b100000000;
assign micromat[37][69] = 9'b111111111;
assign micromat[37][70] = 9'b111111111;
assign micromat[37][71] = 9'b101101101;
assign micromat[37][72] = 9'b100000000;
assign micromat[37][73] = 9'b100100100;
assign micromat[37][74] = 9'b111111111;
assign micromat[37][75] = 9'b111111111;
assign micromat[37][76] = 9'b111111111;
assign micromat[37][77] = 9'b111111111;
assign micromat[37][78] = 9'b110010001;
assign micromat[37][79] = 9'b100000000;
assign micromat[37][80] = 9'b100000000;
assign micromat[37][81] = 9'b110010010;
assign micromat[37][82] = 9'b111111111;
assign micromat[37][83] = 9'b101001001;
assign micromat[37][84] = 9'b100000000;
assign micromat[37][85] = 9'b100100100;
assign micromat[37][86] = 9'b111111111;
assign micromat[37][87] = 9'b111111111;
assign micromat[37][88] = 9'b111111111;
assign micromat[37][89] = 9'b111111111;
assign micromat[37][90] = 9'b111111111;
assign micromat[37][91] = 9'b111111111;
assign micromat[37][92] = 9'b111111111;
assign micromat[37][93] = 9'b111111111;
assign micromat[37][94] = 9'b111111111;
assign micromat[37][95] = 9'b111111111;
assign micromat[37][96] = 9'b111111111;
assign micromat[37][97] = 9'b111111111;
assign micromat[37][98] = 9'b111111111;
assign micromat[37][99] = 9'b111111111;
assign micromat[38][0] = 9'b111111111;
assign micromat[38][1] = 9'b111111111;
assign micromat[38][2] = 9'b111111111;
assign micromat[38][3] = 9'b111111111;
assign micromat[38][4] = 9'b111111111;
assign micromat[38][5] = 9'b111111111;
assign micromat[38][6] = 9'b111111111;
assign micromat[38][7] = 9'b111111111;
assign micromat[38][8] = 9'b111111111;
assign micromat[38][9] = 9'b111111111;
assign micromat[38][10] = 9'b111111111;
assign micromat[38][11] = 9'b111111111;
assign micromat[38][12] = 9'b111111111;
assign micromat[38][13] = 9'b111111111;
assign micromat[38][14] = 9'b100100100;
assign micromat[38][15] = 9'b100000000;
assign micromat[38][16] = 9'b101101101;
assign micromat[38][17] = 9'b111111111;
assign micromat[38][18] = 9'b111111111;
assign micromat[38][19] = 9'b111111111;
assign micromat[38][20] = 9'b111111111;
assign micromat[38][21] = 9'b100101000;
assign micromat[38][22] = 9'b100000000;
assign micromat[38][23] = 9'b100100100;
assign micromat[38][24] = 9'b101101101;
assign micromat[38][25] = 9'b101001001;
assign micromat[38][26] = 9'b101001001;
assign micromat[38][27] = 9'b101001001;
assign micromat[38][28] = 9'b101001001;
assign micromat[38][29] = 9'b101001001;
assign micromat[38][30] = 9'b101001001;
assign micromat[38][31] = 9'b101001001;
assign micromat[38][32] = 9'b101001001;
assign micromat[38][33] = 9'b101001001;
assign micromat[38][34] = 9'b101001001;
assign micromat[38][35] = 9'b101001001;
assign micromat[38][36] = 9'b101001001;
assign micromat[38][37] = 9'b101001001;
assign micromat[38][38] = 9'b101001001;
assign micromat[38][39] = 9'b101001001;
assign micromat[38][40] = 9'b101001001;
assign micromat[38][41] = 9'b101001001;
assign micromat[38][42] = 9'b101001001;
assign micromat[38][43] = 9'b101001001;
assign micromat[38][44] = 9'b101001001;
assign micromat[38][45] = 9'b101001001;
assign micromat[38][46] = 9'b101001001;
assign micromat[38][47] = 9'b101001001;
assign micromat[38][48] = 9'b101001001;
assign micromat[38][49] = 9'b101001001;
assign micromat[38][50] = 9'b101001001;
assign micromat[38][51] = 9'b101001001;
assign micromat[38][52] = 9'b101001001;
assign micromat[38][53] = 9'b101001001;
assign micromat[38][54] = 9'b101001001;
assign micromat[38][55] = 9'b101001001;
assign micromat[38][56] = 9'b101001001;
assign micromat[38][57] = 9'b101101101;
assign micromat[38][58] = 9'b101101101;
assign micromat[38][59] = 9'b100100100;
assign micromat[38][60] = 9'b100000000;
assign micromat[38][61] = 9'b100000000;
assign micromat[38][62] = 9'b110111111;
assign micromat[38][63] = 9'b111111111;
assign micromat[38][64] = 9'b110110111;
assign micromat[38][65] = 9'b110110111;
assign micromat[38][66] = 9'b101101101;
assign micromat[38][67] = 9'b100000000;
assign micromat[38][68] = 9'b100000000;
assign micromat[38][69] = 9'b111111111;
assign micromat[38][70] = 9'b111111111;
assign micromat[38][71] = 9'b101101101;
assign micromat[38][72] = 9'b100000000;
assign micromat[38][73] = 9'b100000000;
assign micromat[38][74] = 9'b111111111;
assign micromat[38][75] = 9'b111111111;
assign micromat[38][76] = 9'b110110111;
assign micromat[38][77] = 9'b110111111;
assign micromat[38][78] = 9'b101101101;
assign micromat[38][79] = 9'b100000000;
assign micromat[38][80] = 9'b100000000;
assign micromat[38][81] = 9'b110010010;
assign micromat[38][82] = 9'b111111111;
assign micromat[38][83] = 9'b101001001;
assign micromat[38][84] = 9'b100000000;
assign micromat[38][85] = 9'b100100100;
assign micromat[38][86] = 9'b111111111;
assign micromat[38][87] = 9'b111111111;
assign micromat[38][88] = 9'b111111111;
assign micromat[38][89] = 9'b111111111;
assign micromat[38][90] = 9'b111111111;
assign micromat[38][91] = 9'b111111111;
assign micromat[38][92] = 9'b111111111;
assign micromat[38][93] = 9'b111111111;
assign micromat[38][94] = 9'b111111111;
assign micromat[38][95] = 9'b111111111;
assign micromat[38][96] = 9'b111111111;
assign micromat[38][97] = 9'b111111111;
assign micromat[38][98] = 9'b111111111;
assign micromat[38][99] = 9'b111111111;
assign micromat[39][0] = 9'b111111111;
assign micromat[39][1] = 9'b111111111;
assign micromat[39][2] = 9'b111111111;
assign micromat[39][3] = 9'b111111111;
assign micromat[39][4] = 9'b111111111;
assign micromat[39][5] = 9'b111111111;
assign micromat[39][6] = 9'b111111111;
assign micromat[39][7] = 9'b111111111;
assign micromat[39][8] = 9'b111111111;
assign micromat[39][9] = 9'b111111111;
assign micromat[39][10] = 9'b111111111;
assign micromat[39][11] = 9'b111111111;
assign micromat[39][12] = 9'b111111111;
assign micromat[39][13] = 9'b111111111;
assign micromat[39][14] = 9'b100100100;
assign micromat[39][15] = 9'b100000000;
assign micromat[39][16] = 9'b101101101;
assign micromat[39][17] = 9'b111111111;
assign micromat[39][18] = 9'b111111111;
assign micromat[39][19] = 9'b111111111;
assign micromat[39][20] = 9'b111111111;
assign micromat[39][21] = 9'b100101000;
assign micromat[39][22] = 9'b100000000;
assign micromat[39][23] = 9'b100100100;
assign micromat[39][24] = 9'b101101101;
assign micromat[39][25] = 9'b101101101;
assign micromat[39][26] = 9'b101101101;
assign micromat[39][27] = 9'b101101101;
assign micromat[39][28] = 9'b101101101;
assign micromat[39][29] = 9'b101101101;
assign micromat[39][30] = 9'b101101101;
assign micromat[39][31] = 9'b101101101;
assign micromat[39][32] = 9'b101101101;
assign micromat[39][33] = 9'b101101101;
assign micromat[39][34] = 9'b101101101;
assign micromat[39][35] = 9'b101101101;
assign micromat[39][36] = 9'b101101101;
assign micromat[39][37] = 9'b101101101;
assign micromat[39][38] = 9'b101101101;
assign micromat[39][39] = 9'b101101101;
assign micromat[39][40] = 9'b101101101;
assign micromat[39][41] = 9'b101101101;
assign micromat[39][42] = 9'b101101101;
assign micromat[39][43] = 9'b101101101;
assign micromat[39][44] = 9'b101101101;
assign micromat[39][45] = 9'b101101101;
assign micromat[39][46] = 9'b101101101;
assign micromat[39][47] = 9'b101101101;
assign micromat[39][48] = 9'b101101101;
assign micromat[39][49] = 9'b101101101;
assign micromat[39][50] = 9'b101101101;
assign micromat[39][51] = 9'b101101101;
assign micromat[39][52] = 9'b101101101;
assign micromat[39][53] = 9'b101101101;
assign micromat[39][54] = 9'b101101101;
assign micromat[39][55] = 9'b101101101;
assign micromat[39][56] = 9'b101101101;
assign micromat[39][57] = 9'b101101101;
assign micromat[39][58] = 9'b101101101;
assign micromat[39][59] = 9'b101001000;
assign micromat[39][60] = 9'b100000000;
assign micromat[39][61] = 9'b100000000;
assign micromat[39][62] = 9'b110111111;
assign micromat[39][63] = 9'b111111111;
assign micromat[39][64] = 9'b110110111;
assign micromat[39][65] = 9'b110110111;
assign micromat[39][66] = 9'b101101101;
assign micromat[39][67] = 9'b100000000;
assign micromat[39][68] = 9'b100000000;
assign micromat[39][69] = 9'b111111111;
assign micromat[39][70] = 9'b111111111;
assign micromat[39][71] = 9'b101101101;
assign micromat[39][72] = 9'b100000000;
assign micromat[39][73] = 9'b100000000;
assign micromat[39][74] = 9'b111111111;
assign micromat[39][75] = 9'b111111111;
assign micromat[39][76] = 9'b111111111;
assign micromat[39][77] = 9'b111111111;
assign micromat[39][78] = 9'b101101101;
assign micromat[39][79] = 9'b100000000;
assign micromat[39][80] = 9'b100000000;
assign micromat[39][81] = 9'b110010010;
assign micromat[39][82] = 9'b111111111;
assign micromat[39][83] = 9'b101001001;
assign micromat[39][84] = 9'b100000000;
assign micromat[39][85] = 9'b100100100;
assign micromat[39][86] = 9'b111111111;
assign micromat[39][87] = 9'b111111111;
assign micromat[39][88] = 9'b111111111;
assign micromat[39][89] = 9'b111111111;
assign micromat[39][90] = 9'b111111111;
assign micromat[39][91] = 9'b111111111;
assign micromat[39][92] = 9'b111111111;
assign micromat[39][93] = 9'b111111111;
assign micromat[39][94] = 9'b111111111;
assign micromat[39][95] = 9'b111111111;
assign micromat[39][96] = 9'b111111111;
assign micromat[39][97] = 9'b111111111;
assign micromat[39][98] = 9'b111111111;
assign micromat[39][99] = 9'b111111111;
assign micromat[40][0] = 9'b111111111;
assign micromat[40][1] = 9'b111111111;
assign micromat[40][2] = 9'b111111111;
assign micromat[40][3] = 9'b111111111;
assign micromat[40][4] = 9'b111111111;
assign micromat[40][5] = 9'b111111111;
assign micromat[40][6] = 9'b111111111;
assign micromat[40][7] = 9'b111111111;
assign micromat[40][8] = 9'b111111111;
assign micromat[40][9] = 9'b111111111;
assign micromat[40][10] = 9'b111111111;
assign micromat[40][11] = 9'b111111111;
assign micromat[40][12] = 9'b111111111;
assign micromat[40][13] = 9'b111111111;
assign micromat[40][14] = 9'b100100100;
assign micromat[40][15] = 9'b100000000;
assign micromat[40][16] = 9'b101101101;
assign micromat[40][17] = 9'b111111111;
assign micromat[40][18] = 9'b111111111;
assign micromat[40][19] = 9'b111111111;
assign micromat[40][20] = 9'b111111111;
assign micromat[40][21] = 9'b100101000;
assign micromat[40][22] = 9'b100000000;
assign micromat[40][23] = 9'b100100100;
assign micromat[40][24] = 9'b101101101;
assign micromat[40][25] = 9'b101101101;
assign micromat[40][26] = 9'b101101101;
assign micromat[40][27] = 9'b101101101;
assign micromat[40][28] = 9'b101101101;
assign micromat[40][29] = 9'b101101101;
assign micromat[40][30] = 9'b101101101;
assign micromat[40][31] = 9'b101101101;
assign micromat[40][32] = 9'b101101101;
assign micromat[40][33] = 9'b101101101;
assign micromat[40][34] = 9'b101101101;
assign micromat[40][35] = 9'b101101101;
assign micromat[40][36] = 9'b101101101;
assign micromat[40][37] = 9'b101101101;
assign micromat[40][38] = 9'b101101101;
assign micromat[40][39] = 9'b101101101;
assign micromat[40][40] = 9'b101101101;
assign micromat[40][41] = 9'b101101101;
assign micromat[40][42] = 9'b101101101;
assign micromat[40][43] = 9'b101101101;
assign micromat[40][44] = 9'b101101101;
assign micromat[40][45] = 9'b101101101;
assign micromat[40][46] = 9'b101101101;
assign micromat[40][47] = 9'b101101101;
assign micromat[40][48] = 9'b101101101;
assign micromat[40][49] = 9'b101101101;
assign micromat[40][50] = 9'b101101101;
assign micromat[40][51] = 9'b101101101;
assign micromat[40][52] = 9'b101101101;
assign micromat[40][53] = 9'b101101101;
assign micromat[40][54] = 9'b101101101;
assign micromat[40][55] = 9'b101101101;
assign micromat[40][56] = 9'b101101101;
assign micromat[40][57] = 9'b110010001;
assign micromat[40][58] = 9'b110010001;
assign micromat[40][59] = 9'b101001001;
assign micromat[40][60] = 9'b100000000;
assign micromat[40][61] = 9'b100000000;
assign micromat[40][62] = 9'b110111111;
assign micromat[40][63] = 9'b111111111;
assign micromat[40][64] = 9'b110110111;
assign micromat[40][65] = 9'b110110111;
assign micromat[40][66] = 9'b101101101;
assign micromat[40][67] = 9'b100000000;
assign micromat[40][68] = 9'b100000000;
assign micromat[40][69] = 9'b111111111;
assign micromat[40][70] = 9'b111111111;
assign micromat[40][71] = 9'b110110110;
assign micromat[40][72] = 9'b101101101;
assign micromat[40][73] = 9'b101101101;
assign micromat[40][74] = 9'b101001001;
assign micromat[40][75] = 9'b101001001;
assign micromat[40][76] = 9'b101001001;
assign micromat[40][77] = 9'b101001001;
assign micromat[40][78] = 9'b101001001;
assign micromat[40][79] = 9'b101101101;
assign micromat[40][80] = 9'b101101101;
assign micromat[40][81] = 9'b110010010;
assign micromat[40][82] = 9'b110111111;
assign micromat[40][83] = 9'b101001001;
assign micromat[40][84] = 9'b100000000;
assign micromat[40][85] = 9'b100100100;
assign micromat[40][86] = 9'b111111111;
assign micromat[40][87] = 9'b111111111;
assign micromat[40][88] = 9'b111111111;
assign micromat[40][89] = 9'b111111111;
assign micromat[40][90] = 9'b111111111;
assign micromat[40][91] = 9'b111111111;
assign micromat[40][92] = 9'b111111111;
assign micromat[40][93] = 9'b111111111;
assign micromat[40][94] = 9'b111111111;
assign micromat[40][95] = 9'b111111111;
assign micromat[40][96] = 9'b111111111;
assign micromat[40][97] = 9'b111111111;
assign micromat[40][98] = 9'b111111111;
assign micromat[40][99] = 9'b111111111;
assign micromat[41][0] = 9'b111111111;
assign micromat[41][1] = 9'b111111111;
assign micromat[41][2] = 9'b111111111;
assign micromat[41][3] = 9'b111111111;
assign micromat[41][4] = 9'b111111111;
assign micromat[41][5] = 9'b111111111;
assign micromat[41][6] = 9'b111111111;
assign micromat[41][7] = 9'b111111111;
assign micromat[41][8] = 9'b111111111;
assign micromat[41][9] = 9'b111111111;
assign micromat[41][10] = 9'b111111111;
assign micromat[41][11] = 9'b111111111;
assign micromat[41][12] = 9'b111111111;
assign micromat[41][13] = 9'b111111111;
assign micromat[41][14] = 9'b100100100;
assign micromat[41][15] = 9'b100000000;
assign micromat[41][16] = 9'b101101101;
assign micromat[41][17] = 9'b111111111;
assign micromat[41][18] = 9'b111111111;
assign micromat[41][19] = 9'b111111111;
assign micromat[41][20] = 9'b111111111;
assign micromat[41][21] = 9'b100101000;
assign micromat[41][22] = 9'b100000000;
assign micromat[41][23] = 9'b100100100;
assign micromat[41][24] = 9'b101101101;
assign micromat[41][25] = 9'b101101101;
assign micromat[41][26] = 9'b101101101;
assign micromat[41][27] = 9'b101101101;
assign micromat[41][28] = 9'b101101101;
assign micromat[41][29] = 9'b101101101;
assign micromat[41][30] = 9'b101101101;
assign micromat[41][31] = 9'b101101101;
assign micromat[41][32] = 9'b101101101;
assign micromat[41][33] = 9'b101101101;
assign micromat[41][34] = 9'b101101101;
assign micromat[41][35] = 9'b101101101;
assign micromat[41][36] = 9'b101101101;
assign micromat[41][37] = 9'b101101101;
assign micromat[41][38] = 9'b101101101;
assign micromat[41][39] = 9'b101101101;
assign micromat[41][40] = 9'b101101101;
assign micromat[41][41] = 9'b101101101;
assign micromat[41][42] = 9'b101101101;
assign micromat[41][43] = 9'b101101101;
assign micromat[41][44] = 9'b101101101;
assign micromat[41][45] = 9'b101101101;
assign micromat[41][46] = 9'b101101101;
assign micromat[41][47] = 9'b101101101;
assign micromat[41][48] = 9'b101101101;
assign micromat[41][49] = 9'b101101101;
assign micromat[41][50] = 9'b101101101;
assign micromat[41][51] = 9'b101101101;
assign micromat[41][52] = 9'b101101101;
assign micromat[41][53] = 9'b101101101;
assign micromat[41][54] = 9'b101101101;
assign micromat[41][55] = 9'b101101101;
assign micromat[41][56] = 9'b101101101;
assign micromat[41][57] = 9'b110010001;
assign micromat[41][58] = 9'b110110110;
assign micromat[41][59] = 9'b101001001;
assign micromat[41][60] = 9'b100000000;
assign micromat[41][61] = 9'b100000000;
assign micromat[41][62] = 9'b110111111;
assign micromat[41][63] = 9'b111111111;
assign micromat[41][64] = 9'b110110111;
assign micromat[41][65] = 9'b110110111;
assign micromat[41][66] = 9'b101101101;
assign micromat[41][67] = 9'b100000000;
assign micromat[41][68] = 9'b100000000;
assign micromat[41][69] = 9'b111111111;
assign micromat[41][70] = 9'b111111111;
assign micromat[41][71] = 9'b111111111;
assign micromat[41][72] = 9'b111111111;
assign micromat[41][73] = 9'b110111111;
assign micromat[41][74] = 9'b100000000;
assign micromat[41][75] = 9'b100000000;
assign micromat[41][76] = 9'b100000000;
assign micromat[41][77] = 9'b100000000;
assign micromat[41][78] = 9'b100100100;
assign micromat[41][79] = 9'b111111111;
assign micromat[41][80] = 9'b111111111;
assign micromat[41][81] = 9'b110110111;
assign micromat[41][82] = 9'b110111111;
assign micromat[41][83] = 9'b101001001;
assign micromat[41][84] = 9'b100000000;
assign micromat[41][85] = 9'b100100100;
assign micromat[41][86] = 9'b111111111;
assign micromat[41][87] = 9'b111111111;
assign micromat[41][88] = 9'b111111111;
assign micromat[41][89] = 9'b111111111;
assign micromat[41][90] = 9'b111111111;
assign micromat[41][91] = 9'b111111111;
assign micromat[41][92] = 9'b111111111;
assign micromat[41][93] = 9'b111111111;
assign micromat[41][94] = 9'b111111111;
assign micromat[41][95] = 9'b111111111;
assign micromat[41][96] = 9'b111111111;
assign micromat[41][97] = 9'b111111111;
assign micromat[41][98] = 9'b111111111;
assign micromat[41][99] = 9'b111111111;
assign micromat[42][0] = 9'b111111111;
assign micromat[42][1] = 9'b111111111;
assign micromat[42][2] = 9'b111111111;
assign micromat[42][3] = 9'b111111111;
assign micromat[42][4] = 9'b111111111;
assign micromat[42][5] = 9'b111111111;
assign micromat[42][6] = 9'b111111111;
assign micromat[42][7] = 9'b111111111;
assign micromat[42][8] = 9'b111111111;
assign micromat[42][9] = 9'b111111111;
assign micromat[42][10] = 9'b111111111;
assign micromat[42][11] = 9'b111111111;
assign micromat[42][12] = 9'b111111111;
assign micromat[42][13] = 9'b111111111;
assign micromat[42][14] = 9'b100100100;
assign micromat[42][15] = 9'b100000000;
assign micromat[42][16] = 9'b101101101;
assign micromat[42][17] = 9'b111111111;
assign micromat[42][18] = 9'b111111111;
assign micromat[42][19] = 9'b111111111;
assign micromat[42][20] = 9'b111111111;
assign micromat[42][21] = 9'b100101000;
assign micromat[42][22] = 9'b100000000;
assign micromat[42][23] = 9'b100100100;
assign micromat[42][24] = 9'b101101101;
assign micromat[42][25] = 9'b101101101;
assign micromat[42][26] = 9'b101101101;
assign micromat[42][27] = 9'b101101101;
assign micromat[42][28] = 9'b101101101;
assign micromat[42][29] = 9'b101101101;
assign micromat[42][30] = 9'b101101101;
assign micromat[42][31] = 9'b101101101;
assign micromat[42][32] = 9'b101101101;
assign micromat[42][33] = 9'b101101101;
assign micromat[42][34] = 9'b101101101;
assign micromat[42][35] = 9'b101101101;
assign micromat[42][36] = 9'b101101101;
assign micromat[42][37] = 9'b101101101;
assign micromat[42][38] = 9'b101101101;
assign micromat[42][39] = 9'b101101101;
assign micromat[42][40] = 9'b101101101;
assign micromat[42][41] = 9'b101101101;
assign micromat[42][42] = 9'b101101101;
assign micromat[42][43] = 9'b101101101;
assign micromat[42][44] = 9'b101101101;
assign micromat[42][45] = 9'b101101101;
assign micromat[42][46] = 9'b101101101;
assign micromat[42][47] = 9'b101101101;
assign micromat[42][48] = 9'b101101101;
assign micromat[42][49] = 9'b101101101;
assign micromat[42][50] = 9'b101101101;
assign micromat[42][51] = 9'b101101101;
assign micromat[42][52] = 9'b101101101;
assign micromat[42][53] = 9'b101101101;
assign micromat[42][54] = 9'b101101101;
assign micromat[42][55] = 9'b101101101;
assign micromat[42][56] = 9'b101101101;
assign micromat[42][57] = 9'b110010001;
assign micromat[42][58] = 9'b110110110;
assign micromat[42][59] = 9'b101001001;
assign micromat[42][60] = 9'b100000000;
assign micromat[42][61] = 9'b100000000;
assign micromat[42][62] = 9'b110111111;
assign micromat[42][63] = 9'b111111111;
assign micromat[42][64] = 9'b110110111;
assign micromat[42][65] = 9'b110110111;
assign micromat[42][66] = 9'b101101101;
assign micromat[42][67] = 9'b100000000;
assign micromat[42][68] = 9'b100000000;
assign micromat[42][69] = 9'b111111111;
assign micromat[42][70] = 9'b111111111;
assign micromat[42][71] = 9'b111111111;
assign micromat[42][72] = 9'b111111111;
assign micromat[42][73] = 9'b110110111;
assign micromat[42][74] = 9'b100100100;
assign micromat[42][75] = 9'b100100100;
assign micromat[42][76] = 9'b100100100;
assign micromat[42][77] = 9'b100100100;
assign micromat[42][78] = 9'b101001001;
assign micromat[42][79] = 9'b111111111;
assign micromat[42][80] = 9'b111111111;
assign micromat[42][81] = 9'b110110111;
assign micromat[42][82] = 9'b110111111;
assign micromat[42][83] = 9'b101001001;
assign micromat[42][84] = 9'b100000000;
assign micromat[42][85] = 9'b100100100;
assign micromat[42][86] = 9'b111111111;
assign micromat[42][87] = 9'b111111111;
assign micromat[42][88] = 9'b111111111;
assign micromat[42][89] = 9'b111111111;
assign micromat[42][90] = 9'b111111111;
assign micromat[42][91] = 9'b111111111;
assign micromat[42][92] = 9'b111111111;
assign micromat[42][93] = 9'b111111111;
assign micromat[42][94] = 9'b111111111;
assign micromat[42][95] = 9'b111111111;
assign micromat[42][96] = 9'b111111111;
assign micromat[42][97] = 9'b111111111;
assign micromat[42][98] = 9'b111111111;
assign micromat[42][99] = 9'b111111111;
assign micromat[43][0] = 9'b111111111;
assign micromat[43][1] = 9'b111111111;
assign micromat[43][2] = 9'b111111111;
assign micromat[43][3] = 9'b111111111;
assign micromat[43][4] = 9'b111111111;
assign micromat[43][5] = 9'b111111111;
assign micromat[43][6] = 9'b111111111;
assign micromat[43][7] = 9'b111111111;
assign micromat[43][8] = 9'b111111111;
assign micromat[43][9] = 9'b111111111;
assign micromat[43][10] = 9'b111111111;
assign micromat[43][11] = 9'b111111111;
assign micromat[43][12] = 9'b111111111;
assign micromat[43][13] = 9'b111111111;
assign micromat[43][14] = 9'b100100100;
assign micromat[43][15] = 9'b100000000;
assign micromat[43][16] = 9'b101101101;
assign micromat[43][17] = 9'b111111111;
assign micromat[43][18] = 9'b111111111;
assign micromat[43][19] = 9'b111111111;
assign micromat[43][20] = 9'b111111111;
assign micromat[43][21] = 9'b100101000;
assign micromat[43][22] = 9'b100000000;
assign micromat[43][23] = 9'b100100100;
assign micromat[43][24] = 9'b101101101;
assign micromat[43][25] = 9'b101101101;
assign micromat[43][26] = 9'b101101101;
assign micromat[43][27] = 9'b101101101;
assign micromat[43][28] = 9'b101101101;
assign micromat[43][29] = 9'b101101101;
assign micromat[43][30] = 9'b101101101;
assign micromat[43][31] = 9'b101101101;
assign micromat[43][32] = 9'b101101101;
assign micromat[43][33] = 9'b101101101;
assign micromat[43][34] = 9'b101101101;
assign micromat[43][35] = 9'b101101101;
assign micromat[43][36] = 9'b101101101;
assign micromat[43][37] = 9'b101101101;
assign micromat[43][38] = 9'b101101101;
assign micromat[43][39] = 9'b101101101;
assign micromat[43][40] = 9'b101101101;
assign micromat[43][41] = 9'b101101101;
assign micromat[43][42] = 9'b101101101;
assign micromat[43][43] = 9'b101101101;
assign micromat[43][44] = 9'b101101101;
assign micromat[43][45] = 9'b101101101;
assign micromat[43][46] = 9'b101101101;
assign micromat[43][47] = 9'b101101101;
assign micromat[43][48] = 9'b101101101;
assign micromat[43][49] = 9'b101101101;
assign micromat[43][50] = 9'b101101101;
assign micromat[43][51] = 9'b101101101;
assign micromat[43][52] = 9'b101101101;
assign micromat[43][53] = 9'b101101101;
assign micromat[43][54] = 9'b101101101;
assign micromat[43][55] = 9'b101101101;
assign micromat[43][56] = 9'b101101101;
assign micromat[43][57] = 9'b110010001;
assign micromat[43][58] = 9'b110110110;
assign micromat[43][59] = 9'b101001001;
assign micromat[43][60] = 9'b100000000;
assign micromat[43][61] = 9'b100000000;
assign micromat[43][62] = 9'b110111111;
assign micromat[43][63] = 9'b111111111;
assign micromat[43][64] = 9'b110110111;
assign micromat[43][65] = 9'b110110111;
assign micromat[43][66] = 9'b101101101;
assign micromat[43][67] = 9'b100000000;
assign micromat[43][68] = 9'b100000000;
assign micromat[43][69] = 9'b111111111;
assign micromat[43][70] = 9'b111111111;
assign micromat[43][71] = 9'b111111111;
assign micromat[43][72] = 9'b111111111;
assign micromat[43][73] = 9'b111111111;
assign micromat[43][74] = 9'b111111111;
assign micromat[43][75] = 9'b111111111;
assign micromat[43][76] = 9'b111111111;
assign micromat[43][77] = 9'b111111111;
assign micromat[43][78] = 9'b111111111;
assign micromat[43][79] = 9'b111111111;
assign micromat[43][80] = 9'b111111111;
assign micromat[43][81] = 9'b110110111;
assign micromat[43][82] = 9'b110111111;
assign micromat[43][83] = 9'b101001001;
assign micromat[43][84] = 9'b100000000;
assign micromat[43][85] = 9'b100100100;
assign micromat[43][86] = 9'b111111111;
assign micromat[43][87] = 9'b111111111;
assign micromat[43][88] = 9'b111111111;
assign micromat[43][89] = 9'b111111111;
assign micromat[43][90] = 9'b111111111;
assign micromat[43][91] = 9'b111111111;
assign micromat[43][92] = 9'b111111111;
assign micromat[43][93] = 9'b111111111;
assign micromat[43][94] = 9'b111111111;
assign micromat[43][95] = 9'b111111111;
assign micromat[43][96] = 9'b111111111;
assign micromat[43][97] = 9'b111111111;
assign micromat[43][98] = 9'b111111111;
assign micromat[43][99] = 9'b111111111;
assign micromat[44][0] = 9'b111111111;
assign micromat[44][1] = 9'b111111111;
assign micromat[44][2] = 9'b111111111;
assign micromat[44][3] = 9'b111111111;
assign micromat[44][4] = 9'b111111111;
assign micromat[44][5] = 9'b111111111;
assign micromat[44][6] = 9'b111111111;
assign micromat[44][7] = 9'b111111111;
assign micromat[44][8] = 9'b111111111;
assign micromat[44][9] = 9'b111111111;
assign micromat[44][10] = 9'b111111111;
assign micromat[44][11] = 9'b111111111;
assign micromat[44][12] = 9'b111111111;
assign micromat[44][13] = 9'b111111111;
assign micromat[44][14] = 9'b100100100;
assign micromat[44][15] = 9'b100000000;
assign micromat[44][16] = 9'b101101101;
assign micromat[44][17] = 9'b111111111;
assign micromat[44][18] = 9'b111111111;
assign micromat[44][19] = 9'b111111111;
assign micromat[44][20] = 9'b111111111;
assign micromat[44][21] = 9'b100101000;
assign micromat[44][22] = 9'b100000000;
assign micromat[44][23] = 9'b100100100;
assign micromat[44][24] = 9'b101101101;
assign micromat[44][25] = 9'b101101101;
assign micromat[44][26] = 9'b101101101;
assign micromat[44][27] = 9'b101101101;
assign micromat[44][28] = 9'b101101101;
assign micromat[44][29] = 9'b101101101;
assign micromat[44][30] = 9'b101101101;
assign micromat[44][31] = 9'b101101101;
assign micromat[44][32] = 9'b101101101;
assign micromat[44][33] = 9'b101101101;
assign micromat[44][34] = 9'b101101101;
assign micromat[44][35] = 9'b101101101;
assign micromat[44][36] = 9'b101101101;
assign micromat[44][37] = 9'b101101101;
assign micromat[44][38] = 9'b101101101;
assign micromat[44][39] = 9'b101101101;
assign micromat[44][40] = 9'b101101101;
assign micromat[44][41] = 9'b101101101;
assign micromat[44][42] = 9'b101101101;
assign micromat[44][43] = 9'b101101101;
assign micromat[44][44] = 9'b101101101;
assign micromat[44][45] = 9'b101101101;
assign micromat[44][46] = 9'b101101101;
assign micromat[44][47] = 9'b101101101;
assign micromat[44][48] = 9'b101101101;
assign micromat[44][49] = 9'b101101101;
assign micromat[44][50] = 9'b101101101;
assign micromat[44][51] = 9'b101101101;
assign micromat[44][52] = 9'b101101101;
assign micromat[44][53] = 9'b101101101;
assign micromat[44][54] = 9'b101101101;
assign micromat[44][55] = 9'b101101101;
assign micromat[44][56] = 9'b101101101;
assign micromat[44][57] = 9'b110010001;
assign micromat[44][58] = 9'b110110110;
assign micromat[44][59] = 9'b101001001;
assign micromat[44][60] = 9'b100000000;
assign micromat[44][61] = 9'b100000000;
assign micromat[44][62] = 9'b110111111;
assign micromat[44][63] = 9'b111111111;
assign micromat[44][64] = 9'b110110111;
assign micromat[44][65] = 9'b110110111;
assign micromat[44][66] = 9'b101101101;
assign micromat[44][67] = 9'b100000000;
assign micromat[44][68] = 9'b100000000;
assign micromat[44][69] = 9'b111111111;
assign micromat[44][70] = 9'b111111111;
assign micromat[44][71] = 9'b111111111;
assign micromat[44][72] = 9'b111111111;
assign micromat[44][73] = 9'b111111111;
assign micromat[44][74] = 9'b111111111;
assign micromat[44][75] = 9'b111111111;
assign micromat[44][76] = 9'b111111111;
assign micromat[44][77] = 9'b111111111;
assign micromat[44][78] = 9'b111111111;
assign micromat[44][79] = 9'b111111111;
assign micromat[44][80] = 9'b111111111;
assign micromat[44][81] = 9'b110110111;
assign micromat[44][82] = 9'b110111111;
assign micromat[44][83] = 9'b101001001;
assign micromat[44][84] = 9'b100000000;
assign micromat[44][85] = 9'b100100100;
assign micromat[44][86] = 9'b111111111;
assign micromat[44][87] = 9'b111111111;
assign micromat[44][88] = 9'b111111111;
assign micromat[44][89] = 9'b111111111;
assign micromat[44][90] = 9'b111111111;
assign micromat[44][91] = 9'b111111111;
assign micromat[44][92] = 9'b111111111;
assign micromat[44][93] = 9'b111111111;
assign micromat[44][94] = 9'b111111111;
assign micromat[44][95] = 9'b111111111;
assign micromat[44][96] = 9'b111111111;
assign micromat[44][97] = 9'b111111111;
assign micromat[44][98] = 9'b111111111;
assign micromat[44][99] = 9'b111111111;
assign micromat[45][0] = 9'b111111111;
assign micromat[45][1] = 9'b111111111;
assign micromat[45][2] = 9'b111111111;
assign micromat[45][3] = 9'b111111111;
assign micromat[45][4] = 9'b111111111;
assign micromat[45][5] = 9'b111111111;
assign micromat[45][6] = 9'b111111111;
assign micromat[45][7] = 9'b111111111;
assign micromat[45][8] = 9'b111111111;
assign micromat[45][9] = 9'b111111111;
assign micromat[45][10] = 9'b111111111;
assign micromat[45][11] = 9'b111111111;
assign micromat[45][12] = 9'b111111111;
assign micromat[45][13] = 9'b111111111;
assign micromat[45][14] = 9'b100100100;
assign micromat[45][15] = 9'b100000000;
assign micromat[45][16] = 9'b101101101;
assign micromat[45][17] = 9'b111111111;
assign micromat[45][18] = 9'b111111111;
assign micromat[45][19] = 9'b111111111;
assign micromat[45][20] = 9'b111111111;
assign micromat[45][21] = 9'b100101000;
assign micromat[45][22] = 9'b100000000;
assign micromat[45][23] = 9'b100100100;
assign micromat[45][24] = 9'b101101101;
assign micromat[45][25] = 9'b101101101;
assign micromat[45][26] = 9'b101101101;
assign micromat[45][27] = 9'b101101101;
assign micromat[45][28] = 9'b101101101;
assign micromat[45][29] = 9'b101101101;
assign micromat[45][30] = 9'b101101101;
assign micromat[45][31] = 9'b101101101;
assign micromat[45][32] = 9'b101101101;
assign micromat[45][33] = 9'b101101101;
assign micromat[45][34] = 9'b101101101;
assign micromat[45][35] = 9'b101101101;
assign micromat[45][36] = 9'b101101101;
assign micromat[45][37] = 9'b101101101;
assign micromat[45][38] = 9'b101101101;
assign micromat[45][39] = 9'b101101101;
assign micromat[45][40] = 9'b101101101;
assign micromat[45][41] = 9'b101101101;
assign micromat[45][42] = 9'b101101101;
assign micromat[45][43] = 9'b101101101;
assign micromat[45][44] = 9'b101101101;
assign micromat[45][45] = 9'b101101101;
assign micromat[45][46] = 9'b101101101;
assign micromat[45][47] = 9'b101101101;
assign micromat[45][48] = 9'b101101101;
assign micromat[45][49] = 9'b101101101;
assign micromat[45][50] = 9'b101101101;
assign micromat[45][51] = 9'b101101101;
assign micromat[45][52] = 9'b101101101;
assign micromat[45][53] = 9'b101101101;
assign micromat[45][54] = 9'b101101101;
assign micromat[45][55] = 9'b101101101;
assign micromat[45][56] = 9'b101101101;
assign micromat[45][57] = 9'b110010001;
assign micromat[45][58] = 9'b110110110;
assign micromat[45][59] = 9'b101001001;
assign micromat[45][60] = 9'b100000000;
assign micromat[45][61] = 9'b100000000;
assign micromat[45][62] = 9'b110111111;
assign micromat[45][63] = 9'b111111111;
assign micromat[45][64] = 9'b110110111;
assign micromat[45][65] = 9'b110110111;
assign micromat[45][66] = 9'b101101101;
assign micromat[45][67] = 9'b100000000;
assign micromat[45][68] = 9'b100000000;
assign micromat[45][69] = 9'b111111111;
assign micromat[45][70] = 9'b111111111;
assign micromat[45][71] = 9'b111111111;
assign micromat[45][72] = 9'b111111111;
assign micromat[45][73] = 9'b110110111;
assign micromat[45][74] = 9'b100100100;
assign micromat[45][75] = 9'b100100100;
assign micromat[45][76] = 9'b100100100;
assign micromat[45][77] = 9'b100100100;
assign micromat[45][78] = 9'b101001101;
assign micromat[45][79] = 9'b111111111;
assign micromat[45][80] = 9'b111111111;
assign micromat[45][81] = 9'b110110111;
assign micromat[45][82] = 9'b110111111;
assign micromat[45][83] = 9'b101001001;
assign micromat[45][84] = 9'b100000000;
assign micromat[45][85] = 9'b100100100;
assign micromat[45][86] = 9'b111111111;
assign micromat[45][87] = 9'b111111111;
assign micromat[45][88] = 9'b111111111;
assign micromat[45][89] = 9'b111111111;
assign micromat[45][90] = 9'b111111111;
assign micromat[45][91] = 9'b111111111;
assign micromat[45][92] = 9'b111111111;
assign micromat[45][93] = 9'b111111111;
assign micromat[45][94] = 9'b111111111;
assign micromat[45][95] = 9'b111111111;
assign micromat[45][96] = 9'b111111111;
assign micromat[45][97] = 9'b111111111;
assign micromat[45][98] = 9'b111111111;
assign micromat[45][99] = 9'b111111111;
assign micromat[46][0] = 9'b111111111;
assign micromat[46][1] = 9'b111111111;
assign micromat[46][2] = 9'b111111111;
assign micromat[46][3] = 9'b111111111;
assign micromat[46][4] = 9'b111111111;
assign micromat[46][5] = 9'b111111111;
assign micromat[46][6] = 9'b111111111;
assign micromat[46][7] = 9'b111111111;
assign micromat[46][8] = 9'b111111111;
assign micromat[46][9] = 9'b111111111;
assign micromat[46][10] = 9'b111111111;
assign micromat[46][11] = 9'b111111111;
assign micromat[46][12] = 9'b111111111;
assign micromat[46][13] = 9'b111111111;
assign micromat[46][14] = 9'b100100100;
assign micromat[46][15] = 9'b100000000;
assign micromat[46][16] = 9'b101101101;
assign micromat[46][17] = 9'b111111111;
assign micromat[46][18] = 9'b111111111;
assign micromat[46][19] = 9'b111111111;
assign micromat[46][20] = 9'b111111111;
assign micromat[46][21] = 9'b100101000;
assign micromat[46][22] = 9'b100000000;
assign micromat[46][23] = 9'b100100100;
assign micromat[46][24] = 9'b101101101;
assign micromat[46][25] = 9'b101101101;
assign micromat[46][26] = 9'b101101101;
assign micromat[46][27] = 9'b101101101;
assign micromat[46][28] = 9'b101101101;
assign micromat[46][29] = 9'b101101101;
assign micromat[46][30] = 9'b101101101;
assign micromat[46][31] = 9'b101101101;
assign micromat[46][32] = 9'b101101101;
assign micromat[46][33] = 9'b101101101;
assign micromat[46][34] = 9'b101101101;
assign micromat[46][35] = 9'b101101101;
assign micromat[46][36] = 9'b101101101;
assign micromat[46][37] = 9'b101101101;
assign micromat[46][38] = 9'b101101101;
assign micromat[46][39] = 9'b101101101;
assign micromat[46][40] = 9'b101101101;
assign micromat[46][41] = 9'b101101101;
assign micromat[46][42] = 9'b101101101;
assign micromat[46][43] = 9'b101101101;
assign micromat[46][44] = 9'b101101101;
assign micromat[46][45] = 9'b101101101;
assign micromat[46][46] = 9'b101101101;
assign micromat[46][47] = 9'b101101101;
assign micromat[46][48] = 9'b101101101;
assign micromat[46][49] = 9'b101101101;
assign micromat[46][50] = 9'b101101101;
assign micromat[46][51] = 9'b101101101;
assign micromat[46][52] = 9'b101101101;
assign micromat[46][53] = 9'b101101101;
assign micromat[46][54] = 9'b101101101;
assign micromat[46][55] = 9'b101101101;
assign micromat[46][56] = 9'b101101101;
assign micromat[46][57] = 9'b110010001;
assign micromat[46][58] = 9'b110110110;
assign micromat[46][59] = 9'b101001001;
assign micromat[46][60] = 9'b100000000;
assign micromat[46][61] = 9'b100000000;
assign micromat[46][62] = 9'b110111111;
assign micromat[46][63] = 9'b111111111;
assign micromat[46][64] = 9'b110110111;
assign micromat[46][65] = 9'b110110111;
assign micromat[46][66] = 9'b101101101;
assign micromat[46][67] = 9'b100000000;
assign micromat[46][68] = 9'b100000000;
assign micromat[46][69] = 9'b111111111;
assign micromat[46][70] = 9'b111111111;
assign micromat[46][71] = 9'b111111111;
assign micromat[46][72] = 9'b111111111;
assign micromat[46][73] = 9'b110111111;
assign micromat[46][74] = 9'b100000000;
assign micromat[46][75] = 9'b100000000;
assign micromat[46][76] = 9'b100000000;
assign micromat[46][77] = 9'b100000000;
assign micromat[46][78] = 9'b100100100;
assign micromat[46][79] = 9'b111111111;
assign micromat[46][80] = 9'b111111111;
assign micromat[46][81] = 9'b110110111;
assign micromat[46][82] = 9'b110111111;
assign micromat[46][83] = 9'b101001001;
assign micromat[46][84] = 9'b100000000;
assign micromat[46][85] = 9'b100100100;
assign micromat[46][86] = 9'b111111111;
assign micromat[46][87] = 9'b111111111;
assign micromat[46][88] = 9'b111111111;
assign micromat[46][89] = 9'b111111111;
assign micromat[46][90] = 9'b111111111;
assign micromat[46][91] = 9'b111111111;
assign micromat[46][92] = 9'b111111111;
assign micromat[46][93] = 9'b111111111;
assign micromat[46][94] = 9'b111111111;
assign micromat[46][95] = 9'b111111111;
assign micromat[46][96] = 9'b111111111;
assign micromat[46][97] = 9'b111111111;
assign micromat[46][98] = 9'b111111111;
assign micromat[46][99] = 9'b111111111;
assign micromat[47][0] = 9'b111111111;
assign micromat[47][1] = 9'b111111111;
assign micromat[47][2] = 9'b111111111;
assign micromat[47][3] = 9'b111111111;
assign micromat[47][4] = 9'b111111111;
assign micromat[47][5] = 9'b111111111;
assign micromat[47][6] = 9'b111111111;
assign micromat[47][7] = 9'b111111111;
assign micromat[47][8] = 9'b111111111;
assign micromat[47][9] = 9'b111111111;
assign micromat[47][10] = 9'b111111111;
assign micromat[47][11] = 9'b111111111;
assign micromat[47][12] = 9'b111111111;
assign micromat[47][13] = 9'b111111111;
assign micromat[47][14] = 9'b100100100;
assign micromat[47][15] = 9'b100000000;
assign micromat[47][16] = 9'b101101101;
assign micromat[47][17] = 9'b111111111;
assign micromat[47][18] = 9'b111111111;
assign micromat[47][19] = 9'b111111111;
assign micromat[47][20] = 9'b111111111;
assign micromat[47][21] = 9'b100101000;
assign micromat[47][22] = 9'b100000000;
assign micromat[47][23] = 9'b100100100;
assign micromat[47][24] = 9'b101101101;
assign micromat[47][25] = 9'b101101101;
assign micromat[47][26] = 9'b101101101;
assign micromat[47][27] = 9'b101101101;
assign micromat[47][28] = 9'b101101101;
assign micromat[47][29] = 9'b101101101;
assign micromat[47][30] = 9'b101101101;
assign micromat[47][31] = 9'b101101101;
assign micromat[47][32] = 9'b101101101;
assign micromat[47][33] = 9'b101101101;
assign micromat[47][34] = 9'b101101101;
assign micromat[47][35] = 9'b101101101;
assign micromat[47][36] = 9'b101101101;
assign micromat[47][37] = 9'b101101101;
assign micromat[47][38] = 9'b101101101;
assign micromat[47][39] = 9'b101101101;
assign micromat[47][40] = 9'b101101101;
assign micromat[47][41] = 9'b101101101;
assign micromat[47][42] = 9'b101101101;
assign micromat[47][43] = 9'b101101101;
assign micromat[47][44] = 9'b101101101;
assign micromat[47][45] = 9'b101101101;
assign micromat[47][46] = 9'b101101101;
assign micromat[47][47] = 9'b101101101;
assign micromat[47][48] = 9'b101101101;
assign micromat[47][49] = 9'b101101101;
assign micromat[47][50] = 9'b101101101;
assign micromat[47][51] = 9'b101101101;
assign micromat[47][52] = 9'b101101101;
assign micromat[47][53] = 9'b101101101;
assign micromat[47][54] = 9'b101101101;
assign micromat[47][55] = 9'b101101101;
assign micromat[47][56] = 9'b101101101;
assign micromat[47][57] = 9'b110010001;
assign micromat[47][58] = 9'b110110110;
assign micromat[47][59] = 9'b101001001;
assign micromat[47][60] = 9'b100000000;
assign micromat[47][61] = 9'b100000000;
assign micromat[47][62] = 9'b110111111;
assign micromat[47][63] = 9'b111111111;
assign micromat[47][64] = 9'b110110111;
assign micromat[47][65] = 9'b110110111;
assign micromat[47][66] = 9'b101101101;
assign micromat[47][67] = 9'b100000000;
assign micromat[47][68] = 9'b100000000;
assign micromat[47][69] = 9'b111111111;
assign micromat[47][70] = 9'b111111111;
assign micromat[47][71] = 9'b110110111;
assign micromat[47][72] = 9'b101101101;
assign micromat[47][73] = 9'b101101101;
assign micromat[47][74] = 9'b101001001;
assign micromat[47][75] = 9'b101001001;
assign micromat[47][76] = 9'b101001001;
assign micromat[47][77] = 9'b101001001;
assign micromat[47][78] = 9'b101001001;
assign micromat[47][79] = 9'b101101101;
assign micromat[47][80] = 9'b101101101;
assign micromat[47][81] = 9'b110010110;
assign micromat[47][82] = 9'b110111111;
assign micromat[47][83] = 9'b101001001;
assign micromat[47][84] = 9'b100000000;
assign micromat[47][85] = 9'b100100100;
assign micromat[47][86] = 9'b111111111;
assign micromat[47][87] = 9'b111111111;
assign micromat[47][88] = 9'b111111111;
assign micromat[47][89] = 9'b111111111;
assign micromat[47][90] = 9'b111111111;
assign micromat[47][91] = 9'b111111111;
assign micromat[47][92] = 9'b111111111;
assign micromat[47][93] = 9'b111111111;
assign micromat[47][94] = 9'b111111111;
assign micromat[47][95] = 9'b111111111;
assign micromat[47][96] = 9'b111111111;
assign micromat[47][97] = 9'b111111111;
assign micromat[47][98] = 9'b111111111;
assign micromat[47][99] = 9'b111111111;
assign micromat[48][0] = 9'b111111111;
assign micromat[48][1] = 9'b111111111;
assign micromat[48][2] = 9'b111111111;
assign micromat[48][3] = 9'b111111111;
assign micromat[48][4] = 9'b111111111;
assign micromat[48][5] = 9'b111111111;
assign micromat[48][6] = 9'b111111111;
assign micromat[48][7] = 9'b111111111;
assign micromat[48][8] = 9'b111111111;
assign micromat[48][9] = 9'b111111111;
assign micromat[48][10] = 9'b111111111;
assign micromat[48][11] = 9'b111111111;
assign micromat[48][12] = 9'b111111111;
assign micromat[48][13] = 9'b111111111;
assign micromat[48][14] = 9'b100100100;
assign micromat[48][15] = 9'b100000000;
assign micromat[48][16] = 9'b101101101;
assign micromat[48][17] = 9'b111111111;
assign micromat[48][18] = 9'b111111111;
assign micromat[48][19] = 9'b111111111;
assign micromat[48][20] = 9'b111111111;
assign micromat[48][21] = 9'b100101000;
assign micromat[48][22] = 9'b100000000;
assign micromat[48][23] = 9'b100100100;
assign micromat[48][24] = 9'b101101101;
assign micromat[48][25] = 9'b101101101;
assign micromat[48][26] = 9'b101101101;
assign micromat[48][27] = 9'b101101101;
assign micromat[48][28] = 9'b101101101;
assign micromat[48][29] = 9'b101101101;
assign micromat[48][30] = 9'b101101101;
assign micromat[48][31] = 9'b101101101;
assign micromat[48][32] = 9'b101101101;
assign micromat[48][33] = 9'b101101101;
assign micromat[48][34] = 9'b101101101;
assign micromat[48][35] = 9'b101101101;
assign micromat[48][36] = 9'b101101101;
assign micromat[48][37] = 9'b101101101;
assign micromat[48][38] = 9'b101101101;
assign micromat[48][39] = 9'b101101101;
assign micromat[48][40] = 9'b101101101;
assign micromat[48][41] = 9'b101101101;
assign micromat[48][42] = 9'b101101101;
assign micromat[48][43] = 9'b101101101;
assign micromat[48][44] = 9'b101101101;
assign micromat[48][45] = 9'b101101101;
assign micromat[48][46] = 9'b101101101;
assign micromat[48][47] = 9'b101101101;
assign micromat[48][48] = 9'b101101101;
assign micromat[48][49] = 9'b101101101;
assign micromat[48][50] = 9'b101101101;
assign micromat[48][51] = 9'b101101101;
assign micromat[48][52] = 9'b101101101;
assign micromat[48][53] = 9'b101101101;
assign micromat[48][54] = 9'b101101101;
assign micromat[48][55] = 9'b101101101;
assign micromat[48][56] = 9'b101101101;
assign micromat[48][57] = 9'b110010001;
assign micromat[48][58] = 9'b110110110;
assign micromat[48][59] = 9'b101001001;
assign micromat[48][60] = 9'b100000000;
assign micromat[48][61] = 9'b100000000;
assign micromat[48][62] = 9'b110111111;
assign micromat[48][63] = 9'b111111111;
assign micromat[48][64] = 9'b110110111;
assign micromat[48][65] = 9'b110110111;
assign micromat[48][66] = 9'b101101101;
assign micromat[48][67] = 9'b100000000;
assign micromat[48][68] = 9'b100000000;
assign micromat[48][69] = 9'b111111111;
assign micromat[48][70] = 9'b111111111;
assign micromat[48][71] = 9'b101101101;
assign micromat[48][72] = 9'b100000000;
assign micromat[48][73] = 9'b100000000;
assign micromat[48][74] = 9'b111111111;
assign micromat[48][75] = 9'b111111111;
assign micromat[48][76] = 9'b111111111;
assign micromat[48][77] = 9'b111111111;
assign micromat[48][78] = 9'b110010010;
assign micromat[48][79] = 9'b100000000;
assign micromat[48][80] = 9'b100000000;
assign micromat[48][81] = 9'b110010010;
assign micromat[48][82] = 9'b111111111;
assign micromat[48][83] = 9'b101001001;
assign micromat[48][84] = 9'b100000000;
assign micromat[48][85] = 9'b100100100;
assign micromat[48][86] = 9'b111111111;
assign micromat[48][87] = 9'b111111111;
assign micromat[48][88] = 9'b111111111;
assign micromat[48][89] = 9'b111111111;
assign micromat[48][90] = 9'b111111111;
assign micromat[48][91] = 9'b111111111;
assign micromat[48][92] = 9'b111111111;
assign micromat[48][93] = 9'b111111111;
assign micromat[48][94] = 9'b111111111;
assign micromat[48][95] = 9'b111111111;
assign micromat[48][96] = 9'b111111111;
assign micromat[48][97] = 9'b111111111;
assign micromat[48][98] = 9'b111111111;
assign micromat[48][99] = 9'b111111111;
assign micromat[49][0] = 9'b111111111;
assign micromat[49][1] = 9'b111111111;
assign micromat[49][2] = 9'b111111111;
assign micromat[49][3] = 9'b111111111;
assign micromat[49][4] = 9'b111111111;
assign micromat[49][5] = 9'b111111111;
assign micromat[49][6] = 9'b111111111;
assign micromat[49][7] = 9'b111111111;
assign micromat[49][8] = 9'b111111111;
assign micromat[49][9] = 9'b111111111;
assign micromat[49][10] = 9'b111111111;
assign micromat[49][11] = 9'b111111111;
assign micromat[49][12] = 9'b111111111;
assign micromat[49][13] = 9'b111111111;
assign micromat[49][14] = 9'b100100100;
assign micromat[49][15] = 9'b100000000;
assign micromat[49][16] = 9'b101101101;
assign micromat[49][17] = 9'b111111111;
assign micromat[49][18] = 9'b111111111;
assign micromat[49][19] = 9'b111111111;
assign micromat[49][20] = 9'b111111111;
assign micromat[49][21] = 9'b100101000;
assign micromat[49][22] = 9'b100000000;
assign micromat[49][23] = 9'b100100100;
assign micromat[49][24] = 9'b101101101;
assign micromat[49][25] = 9'b101101101;
assign micromat[49][26] = 9'b101101101;
assign micromat[49][27] = 9'b101101101;
assign micromat[49][28] = 9'b101101101;
assign micromat[49][29] = 9'b101101101;
assign micromat[49][30] = 9'b101101101;
assign micromat[49][31] = 9'b101101101;
assign micromat[49][32] = 9'b101101101;
assign micromat[49][33] = 9'b101101101;
assign micromat[49][34] = 9'b101101101;
assign micromat[49][35] = 9'b101101101;
assign micromat[49][36] = 9'b101101101;
assign micromat[49][37] = 9'b101101101;
assign micromat[49][38] = 9'b101101101;
assign micromat[49][39] = 9'b101101101;
assign micromat[49][40] = 9'b101101101;
assign micromat[49][41] = 9'b101101101;
assign micromat[49][42] = 9'b101101101;
assign micromat[49][43] = 9'b101101101;
assign micromat[49][44] = 9'b101101101;
assign micromat[49][45] = 9'b101101101;
assign micromat[49][46] = 9'b101101101;
assign micromat[49][47] = 9'b101101101;
assign micromat[49][48] = 9'b101101101;
assign micromat[49][49] = 9'b101101101;
assign micromat[49][50] = 9'b101101101;
assign micromat[49][51] = 9'b101101101;
assign micromat[49][52] = 9'b101101101;
assign micromat[49][53] = 9'b101101101;
assign micromat[49][54] = 9'b101101101;
assign micromat[49][55] = 9'b101101101;
assign micromat[49][56] = 9'b101101101;
assign micromat[49][57] = 9'b110010001;
assign micromat[49][58] = 9'b110110110;
assign micromat[49][59] = 9'b101001001;
assign micromat[49][60] = 9'b100000000;
assign micromat[49][61] = 9'b100000000;
assign micromat[49][62] = 9'b110111111;
assign micromat[49][63] = 9'b111111111;
assign micromat[49][64] = 9'b110110111;
assign micromat[49][65] = 9'b110110111;
assign micromat[49][66] = 9'b101101101;
assign micromat[49][67] = 9'b100000000;
assign micromat[49][68] = 9'b100000000;
assign micromat[49][69] = 9'b111111111;
assign micromat[49][70] = 9'b111111111;
assign micromat[49][71] = 9'b101101101;
assign micromat[49][72] = 9'b100000000;
assign micromat[49][73] = 9'b100000100;
assign micromat[49][74] = 9'b111111111;
assign micromat[49][75] = 9'b111111111;
assign micromat[49][76] = 9'b111111111;
assign micromat[49][77] = 9'b111111111;
assign micromat[49][78] = 9'b110010001;
assign micromat[49][79] = 9'b100000000;
assign micromat[49][80] = 9'b100000000;
assign micromat[49][81] = 9'b110010010;
assign micromat[49][82] = 9'b111111111;
assign micromat[49][83] = 9'b101001001;
assign micromat[49][84] = 9'b100000000;
assign micromat[49][85] = 9'b100100100;
assign micromat[49][86] = 9'b111111111;
assign micromat[49][87] = 9'b111111111;
assign micromat[49][88] = 9'b111111111;
assign micromat[49][89] = 9'b111111111;
assign micromat[49][90] = 9'b111111111;
assign micromat[49][91] = 9'b111111111;
assign micromat[49][92] = 9'b111111111;
assign micromat[49][93] = 9'b111111111;
assign micromat[49][94] = 9'b111111111;
assign micromat[49][95] = 9'b111111111;
assign micromat[49][96] = 9'b111111111;
assign micromat[49][97] = 9'b111111111;
assign micromat[49][98] = 9'b111111111;
assign micromat[49][99] = 9'b111111111;
assign micromat[50][0] = 9'b111111111;
assign micromat[50][1] = 9'b111111111;
assign micromat[50][2] = 9'b111111111;
assign micromat[50][3] = 9'b111111111;
assign micromat[50][4] = 9'b111111111;
assign micromat[50][5] = 9'b111111111;
assign micromat[50][6] = 9'b111111111;
assign micromat[50][7] = 9'b111111111;
assign micromat[50][8] = 9'b111111111;
assign micromat[50][9] = 9'b111111111;
assign micromat[50][10] = 9'b111111111;
assign micromat[50][11] = 9'b111111111;
assign micromat[50][12] = 9'b111111111;
assign micromat[50][13] = 9'b111111111;
assign micromat[50][14] = 9'b100100100;
assign micromat[50][15] = 9'b100000000;
assign micromat[50][16] = 9'b101101101;
assign micromat[50][17] = 9'b111111111;
assign micromat[50][18] = 9'b111111111;
assign micromat[50][19] = 9'b111111111;
assign micromat[50][20] = 9'b111111111;
assign micromat[50][21] = 9'b100101000;
assign micromat[50][22] = 9'b100000000;
assign micromat[50][23] = 9'b100100100;
assign micromat[50][24] = 9'b101101101;
assign micromat[50][25] = 9'b101101101;
assign micromat[50][26] = 9'b101101101;
assign micromat[50][27] = 9'b101101101;
assign micromat[50][28] = 9'b101101101;
assign micromat[50][29] = 9'b101101101;
assign micromat[50][30] = 9'b101101101;
assign micromat[50][31] = 9'b101101101;
assign micromat[50][32] = 9'b101101101;
assign micromat[50][33] = 9'b101101101;
assign micromat[50][34] = 9'b101101101;
assign micromat[50][35] = 9'b101101101;
assign micromat[50][36] = 9'b101101101;
assign micromat[50][37] = 9'b101101101;
assign micromat[50][38] = 9'b101101101;
assign micromat[50][39] = 9'b101101101;
assign micromat[50][40] = 9'b101101101;
assign micromat[50][41] = 9'b101101101;
assign micromat[50][42] = 9'b101101101;
assign micromat[50][43] = 9'b101101101;
assign micromat[50][44] = 9'b101101101;
assign micromat[50][45] = 9'b101101101;
assign micromat[50][46] = 9'b101101101;
assign micromat[50][47] = 9'b101101101;
assign micromat[50][48] = 9'b101101101;
assign micromat[50][49] = 9'b101101101;
assign micromat[50][50] = 9'b101101101;
assign micromat[50][51] = 9'b101101101;
assign micromat[50][52] = 9'b101101101;
assign micromat[50][53] = 9'b101101101;
assign micromat[50][54] = 9'b101101101;
assign micromat[50][55] = 9'b101101101;
assign micromat[50][56] = 9'b101101101;
assign micromat[50][57] = 9'b110010001;
assign micromat[50][58] = 9'b110110110;
assign micromat[50][59] = 9'b101001001;
assign micromat[50][60] = 9'b100000000;
assign micromat[50][61] = 9'b100000000;
assign micromat[50][62] = 9'b110111111;
assign micromat[50][63] = 9'b111111111;
assign micromat[50][64] = 9'b110110111;
assign micromat[50][65] = 9'b110110111;
assign micromat[50][66] = 9'b101101101;
assign micromat[50][67] = 9'b100000000;
assign micromat[50][68] = 9'b100000000;
assign micromat[50][69] = 9'b111111111;
assign micromat[50][70] = 9'b111111111;
assign micromat[50][71] = 9'b101101101;
assign micromat[50][72] = 9'b100000000;
assign micromat[50][73] = 9'b100000000;
assign micromat[50][74] = 9'b111111111;
assign micromat[50][75] = 9'b111111111;
assign micromat[50][76] = 9'b110110111;
assign micromat[50][77] = 9'b110110111;
assign micromat[50][78] = 9'b101101101;
assign micromat[50][79] = 9'b100000000;
assign micromat[50][80] = 9'b100000000;
assign micromat[50][81] = 9'b110010010;
assign micromat[50][82] = 9'b111111111;
assign micromat[50][83] = 9'b101001001;
assign micromat[50][84] = 9'b100000000;
assign micromat[50][85] = 9'b100100100;
assign micromat[50][86] = 9'b111111111;
assign micromat[50][87] = 9'b111111111;
assign micromat[50][88] = 9'b111111111;
assign micromat[50][89] = 9'b111111111;
assign micromat[50][90] = 9'b111111111;
assign micromat[50][91] = 9'b111111111;
assign micromat[50][92] = 9'b111111111;
assign micromat[50][93] = 9'b111111111;
assign micromat[50][94] = 9'b111111111;
assign micromat[50][95] = 9'b111111111;
assign micromat[50][96] = 9'b111111111;
assign micromat[50][97] = 9'b111111111;
assign micromat[50][98] = 9'b111111111;
assign micromat[50][99] = 9'b111111111;
assign micromat[51][0] = 9'b111111111;
assign micromat[51][1] = 9'b111111111;
assign micromat[51][2] = 9'b111111111;
assign micromat[51][3] = 9'b111111111;
assign micromat[51][4] = 9'b111111111;
assign micromat[51][5] = 9'b111111111;
assign micromat[51][6] = 9'b111111111;
assign micromat[51][7] = 9'b111111111;
assign micromat[51][8] = 9'b111111111;
assign micromat[51][9] = 9'b111111111;
assign micromat[51][10] = 9'b111111111;
assign micromat[51][11] = 9'b111111111;
assign micromat[51][12] = 9'b111111111;
assign micromat[51][13] = 9'b111111111;
assign micromat[51][14] = 9'b100100100;
assign micromat[51][15] = 9'b100000000;
assign micromat[51][16] = 9'b101101101;
assign micromat[51][17] = 9'b111111111;
assign micromat[51][18] = 9'b111111111;
assign micromat[51][19] = 9'b111111111;
assign micromat[51][20] = 9'b111111111;
assign micromat[51][21] = 9'b100101000;
assign micromat[51][22] = 9'b100000000;
assign micromat[51][23] = 9'b100100100;
assign micromat[51][24] = 9'b101101101;
assign micromat[51][25] = 9'b101101101;
assign micromat[51][26] = 9'b101101101;
assign micromat[51][27] = 9'b101101101;
assign micromat[51][28] = 9'b101101101;
assign micromat[51][29] = 9'b101101101;
assign micromat[51][30] = 9'b101101101;
assign micromat[51][31] = 9'b101101101;
assign micromat[51][32] = 9'b101101101;
assign micromat[51][33] = 9'b101101101;
assign micromat[51][34] = 9'b101101101;
assign micromat[51][35] = 9'b101101101;
assign micromat[51][36] = 9'b101101101;
assign micromat[51][37] = 9'b101101101;
assign micromat[51][38] = 9'b101101101;
assign micromat[51][39] = 9'b101101101;
assign micromat[51][40] = 9'b101101101;
assign micromat[51][41] = 9'b101101101;
assign micromat[51][42] = 9'b101101101;
assign micromat[51][43] = 9'b101101101;
assign micromat[51][44] = 9'b101101101;
assign micromat[51][45] = 9'b101101101;
assign micromat[51][46] = 9'b101101101;
assign micromat[51][47] = 9'b101101101;
assign micromat[51][48] = 9'b101101101;
assign micromat[51][49] = 9'b101101101;
assign micromat[51][50] = 9'b101101101;
assign micromat[51][51] = 9'b101101101;
assign micromat[51][52] = 9'b101101101;
assign micromat[51][53] = 9'b101101101;
assign micromat[51][54] = 9'b101101101;
assign micromat[51][55] = 9'b101101101;
assign micromat[51][56] = 9'b101101101;
assign micromat[51][57] = 9'b110010001;
assign micromat[51][58] = 9'b110110110;
assign micromat[51][59] = 9'b101001001;
assign micromat[51][60] = 9'b100000000;
assign micromat[51][61] = 9'b100000000;
assign micromat[51][62] = 9'b110111111;
assign micromat[51][63] = 9'b111111111;
assign micromat[51][64] = 9'b110110111;
assign micromat[51][65] = 9'b110110111;
assign micromat[51][66] = 9'b101101101;
assign micromat[51][67] = 9'b100000000;
assign micromat[51][68] = 9'b100000000;
assign micromat[51][69] = 9'b111111111;
assign micromat[51][70] = 9'b111111111;
assign micromat[51][71] = 9'b101101101;
assign micromat[51][72] = 9'b100000000;
assign micromat[51][73] = 9'b100000000;
assign micromat[51][74] = 9'b111111111;
assign micromat[51][75] = 9'b111111111;
assign micromat[51][76] = 9'b111111111;
assign micromat[51][77] = 9'b111111111;
assign micromat[51][78] = 9'b101101101;
assign micromat[51][79] = 9'b100000000;
assign micromat[51][80] = 9'b100000000;
assign micromat[51][81] = 9'b110010010;
assign micromat[51][82] = 9'b111111111;
assign micromat[51][83] = 9'b101001001;
assign micromat[51][84] = 9'b100000000;
assign micromat[51][85] = 9'b100100100;
assign micromat[51][86] = 9'b111111111;
assign micromat[51][87] = 9'b111111111;
assign micromat[51][88] = 9'b111111111;
assign micromat[51][89] = 9'b111111111;
assign micromat[51][90] = 9'b111111111;
assign micromat[51][91] = 9'b111111111;
assign micromat[51][92] = 9'b111111111;
assign micromat[51][93] = 9'b111111111;
assign micromat[51][94] = 9'b111111111;
assign micromat[51][95] = 9'b111111111;
assign micromat[51][96] = 9'b111111111;
assign micromat[51][97] = 9'b111111111;
assign micromat[51][98] = 9'b111111111;
assign micromat[51][99] = 9'b111111111;
assign micromat[52][0] = 9'b111111111;
assign micromat[52][1] = 9'b111111111;
assign micromat[52][2] = 9'b111111111;
assign micromat[52][3] = 9'b111111111;
assign micromat[52][4] = 9'b111111111;
assign micromat[52][5] = 9'b111111111;
assign micromat[52][6] = 9'b111111111;
assign micromat[52][7] = 9'b111111111;
assign micromat[52][8] = 9'b111111111;
assign micromat[52][9] = 9'b111111111;
assign micromat[52][10] = 9'b111111111;
assign micromat[52][11] = 9'b111111111;
assign micromat[52][12] = 9'b111111111;
assign micromat[52][13] = 9'b111111111;
assign micromat[52][14] = 9'b100100100;
assign micromat[52][15] = 9'b100000000;
assign micromat[52][16] = 9'b101101101;
assign micromat[52][17] = 9'b111111111;
assign micromat[52][18] = 9'b111111111;
assign micromat[52][19] = 9'b111111111;
assign micromat[52][20] = 9'b111111111;
assign micromat[52][21] = 9'b100101000;
assign micromat[52][22] = 9'b100000000;
assign micromat[52][23] = 9'b100100100;
assign micromat[52][24] = 9'b101101101;
assign micromat[52][25] = 9'b101101101;
assign micromat[52][26] = 9'b101101101;
assign micromat[52][27] = 9'b101101101;
assign micromat[52][28] = 9'b101101101;
assign micromat[52][29] = 9'b101101101;
assign micromat[52][30] = 9'b101101101;
assign micromat[52][31] = 9'b101101101;
assign micromat[52][32] = 9'b101101101;
assign micromat[52][33] = 9'b101101101;
assign micromat[52][34] = 9'b101101101;
assign micromat[52][35] = 9'b101101101;
assign micromat[52][36] = 9'b101101101;
assign micromat[52][37] = 9'b101101101;
assign micromat[52][38] = 9'b101101101;
assign micromat[52][39] = 9'b101101101;
assign micromat[52][40] = 9'b101101101;
assign micromat[52][41] = 9'b101101101;
assign micromat[52][42] = 9'b101101101;
assign micromat[52][43] = 9'b101101101;
assign micromat[52][44] = 9'b101101101;
assign micromat[52][45] = 9'b101101101;
assign micromat[52][46] = 9'b101101101;
assign micromat[52][47] = 9'b101101101;
assign micromat[52][48] = 9'b101101101;
assign micromat[52][49] = 9'b101101101;
assign micromat[52][50] = 9'b101101101;
assign micromat[52][51] = 9'b101101101;
assign micromat[52][52] = 9'b101101101;
assign micromat[52][53] = 9'b101101101;
assign micromat[52][54] = 9'b101101101;
assign micromat[52][55] = 9'b101101101;
assign micromat[52][56] = 9'b101101101;
assign micromat[52][57] = 9'b110010001;
assign micromat[52][58] = 9'b110110110;
assign micromat[52][59] = 9'b101001001;
assign micromat[52][60] = 9'b100000000;
assign micromat[52][61] = 9'b100000000;
assign micromat[52][62] = 9'b110111111;
assign micromat[52][63] = 9'b111111111;
assign micromat[52][64] = 9'b110110111;
assign micromat[52][65] = 9'b110110111;
assign micromat[52][66] = 9'b101101101;
assign micromat[52][67] = 9'b100000000;
assign micromat[52][68] = 9'b100000000;
assign micromat[52][69] = 9'b111111111;
assign micromat[52][70] = 9'b111111111;
assign micromat[52][71] = 9'b110110111;
assign micromat[52][72] = 9'b101101101;
assign micromat[52][73] = 9'b101101101;
assign micromat[52][74] = 9'b101001001;
assign micromat[52][75] = 9'b101001001;
assign micromat[52][76] = 9'b101001001;
assign micromat[52][77] = 9'b101001001;
assign micromat[52][78] = 9'b101001001;
assign micromat[52][79] = 9'b101101101;
assign micromat[52][80] = 9'b101101101;
assign micromat[52][81] = 9'b110010110;
assign micromat[52][82] = 9'b110111111;
assign micromat[52][83] = 9'b101001001;
assign micromat[52][84] = 9'b100000000;
assign micromat[52][85] = 9'b100100100;
assign micromat[52][86] = 9'b111111111;
assign micromat[52][87] = 9'b111111111;
assign micromat[52][88] = 9'b111111111;
assign micromat[52][89] = 9'b111111111;
assign micromat[52][90] = 9'b111111111;
assign micromat[52][91] = 9'b111111111;
assign micromat[52][92] = 9'b111111111;
assign micromat[52][93] = 9'b111111111;
assign micromat[52][94] = 9'b111111111;
assign micromat[52][95] = 9'b111111111;
assign micromat[52][96] = 9'b111111111;
assign micromat[52][97] = 9'b111111111;
assign micromat[52][98] = 9'b111111111;
assign micromat[52][99] = 9'b111111111;
assign micromat[53][0] = 9'b111111111;
assign micromat[53][1] = 9'b111111111;
assign micromat[53][2] = 9'b111111111;
assign micromat[53][3] = 9'b111111111;
assign micromat[53][4] = 9'b111111111;
assign micromat[53][5] = 9'b111111111;
assign micromat[53][6] = 9'b111111111;
assign micromat[53][7] = 9'b111111111;
assign micromat[53][8] = 9'b111111111;
assign micromat[53][9] = 9'b111111111;
assign micromat[53][10] = 9'b111111111;
assign micromat[53][11] = 9'b111111111;
assign micromat[53][12] = 9'b111111111;
assign micromat[53][13] = 9'b111111111;
assign micromat[53][14] = 9'b100100100;
assign micromat[53][15] = 9'b100000000;
assign micromat[53][16] = 9'b101101101;
assign micromat[53][17] = 9'b111111111;
assign micromat[53][18] = 9'b111111111;
assign micromat[53][19] = 9'b111111111;
assign micromat[53][20] = 9'b111111111;
assign micromat[53][21] = 9'b100101000;
assign micromat[53][22] = 9'b100000000;
assign micromat[53][23] = 9'b100100100;
assign micromat[53][24] = 9'b101101101;
assign micromat[53][25] = 9'b101101101;
assign micromat[53][26] = 9'b101101101;
assign micromat[53][27] = 9'b101101101;
assign micromat[53][28] = 9'b101101101;
assign micromat[53][29] = 9'b101101101;
assign micromat[53][30] = 9'b101101101;
assign micromat[53][31] = 9'b101101101;
assign micromat[53][32] = 9'b101101101;
assign micromat[53][33] = 9'b101101101;
assign micromat[53][34] = 9'b101101101;
assign micromat[53][35] = 9'b101101101;
assign micromat[53][36] = 9'b101101101;
assign micromat[53][37] = 9'b101101101;
assign micromat[53][38] = 9'b101101101;
assign micromat[53][39] = 9'b101101101;
assign micromat[53][40] = 9'b101101101;
assign micromat[53][41] = 9'b101101101;
assign micromat[53][42] = 9'b101101101;
assign micromat[53][43] = 9'b101101101;
assign micromat[53][44] = 9'b101101101;
assign micromat[53][45] = 9'b101101101;
assign micromat[53][46] = 9'b101101101;
assign micromat[53][47] = 9'b101101101;
assign micromat[53][48] = 9'b101101101;
assign micromat[53][49] = 9'b101101101;
assign micromat[53][50] = 9'b101101101;
assign micromat[53][51] = 9'b101101101;
assign micromat[53][52] = 9'b101101101;
assign micromat[53][53] = 9'b101101101;
assign micromat[53][54] = 9'b101101101;
assign micromat[53][55] = 9'b101101101;
assign micromat[53][56] = 9'b101101101;
assign micromat[53][57] = 9'b110010001;
assign micromat[53][58] = 9'b110110110;
assign micromat[53][59] = 9'b101001001;
assign micromat[53][60] = 9'b100000000;
assign micromat[53][61] = 9'b100000000;
assign micromat[53][62] = 9'b110111111;
assign micromat[53][63] = 9'b111111111;
assign micromat[53][64] = 9'b110110111;
assign micromat[53][65] = 9'b110110111;
assign micromat[53][66] = 9'b101101101;
assign micromat[53][67] = 9'b100000000;
assign micromat[53][68] = 9'b100000000;
assign micromat[53][69] = 9'b111111111;
assign micromat[53][70] = 9'b111111111;
assign micromat[53][71] = 9'b111111111;
assign micromat[53][72] = 9'b111111111;
assign micromat[53][73] = 9'b110111111;
assign micromat[53][74] = 9'b100000000;
assign micromat[53][75] = 9'b100000000;
assign micromat[53][76] = 9'b100000000;
assign micromat[53][77] = 9'b100000000;
assign micromat[53][78] = 9'b100100100;
assign micromat[53][79] = 9'b111111111;
assign micromat[53][80] = 9'b111111111;
assign micromat[53][81] = 9'b110110111;
assign micromat[53][82] = 9'b110111111;
assign micromat[53][83] = 9'b101001001;
assign micromat[53][84] = 9'b100000000;
assign micromat[53][85] = 9'b100100100;
assign micromat[53][86] = 9'b111111111;
assign micromat[53][87] = 9'b111111111;
assign micromat[53][88] = 9'b111111111;
assign micromat[53][89] = 9'b111111111;
assign micromat[53][90] = 9'b111111111;
assign micromat[53][91] = 9'b111111111;
assign micromat[53][92] = 9'b111111111;
assign micromat[53][93] = 9'b111111111;
assign micromat[53][94] = 9'b111111111;
assign micromat[53][95] = 9'b111111111;
assign micromat[53][96] = 9'b111111111;
assign micromat[53][97] = 9'b111111111;
assign micromat[53][98] = 9'b111111111;
assign micromat[53][99] = 9'b111111111;
assign micromat[54][0] = 9'b111111111;
assign micromat[54][1] = 9'b111111111;
assign micromat[54][2] = 9'b111111111;
assign micromat[54][3] = 9'b111111111;
assign micromat[54][4] = 9'b111111111;
assign micromat[54][5] = 9'b111111111;
assign micromat[54][6] = 9'b111111111;
assign micromat[54][7] = 9'b111111111;
assign micromat[54][8] = 9'b111111111;
assign micromat[54][9] = 9'b111111111;
assign micromat[54][10] = 9'b111111111;
assign micromat[54][11] = 9'b111111111;
assign micromat[54][12] = 9'b111111111;
assign micromat[54][13] = 9'b111111111;
assign micromat[54][14] = 9'b100100100;
assign micromat[54][15] = 9'b100000000;
assign micromat[54][16] = 9'b101101101;
assign micromat[54][17] = 9'b111111111;
assign micromat[54][18] = 9'b111111111;
assign micromat[54][19] = 9'b111111111;
assign micromat[54][20] = 9'b111111111;
assign micromat[54][21] = 9'b100101000;
assign micromat[54][22] = 9'b100000000;
assign micromat[54][23] = 9'b100100100;
assign micromat[54][24] = 9'b101101101;
assign micromat[54][25] = 9'b101101101;
assign micromat[54][26] = 9'b101101101;
assign micromat[54][27] = 9'b101101101;
assign micromat[54][28] = 9'b101101101;
assign micromat[54][29] = 9'b101101101;
assign micromat[54][30] = 9'b101101101;
assign micromat[54][31] = 9'b101101101;
assign micromat[54][32] = 9'b101101101;
assign micromat[54][33] = 9'b101101101;
assign micromat[54][34] = 9'b101101101;
assign micromat[54][35] = 9'b101101101;
assign micromat[54][36] = 9'b101101101;
assign micromat[54][37] = 9'b101101101;
assign micromat[54][38] = 9'b101101101;
assign micromat[54][39] = 9'b101101101;
assign micromat[54][40] = 9'b101101101;
assign micromat[54][41] = 9'b101101101;
assign micromat[54][42] = 9'b101101101;
assign micromat[54][43] = 9'b101101101;
assign micromat[54][44] = 9'b101101101;
assign micromat[54][45] = 9'b101101101;
assign micromat[54][46] = 9'b101101101;
assign micromat[54][47] = 9'b101101101;
assign micromat[54][48] = 9'b101101101;
assign micromat[54][49] = 9'b101101101;
assign micromat[54][50] = 9'b101101101;
assign micromat[54][51] = 9'b101101101;
assign micromat[54][52] = 9'b101101101;
assign micromat[54][53] = 9'b101101101;
assign micromat[54][54] = 9'b101101101;
assign micromat[54][55] = 9'b101101101;
assign micromat[54][56] = 9'b101101101;
assign micromat[54][57] = 9'b110010001;
assign micromat[54][58] = 9'b110110110;
assign micromat[54][59] = 9'b101001001;
assign micromat[54][60] = 9'b100000000;
assign micromat[54][61] = 9'b100000000;
assign micromat[54][62] = 9'b110111111;
assign micromat[54][63] = 9'b111111111;
assign micromat[54][64] = 9'b110110111;
assign micromat[54][65] = 9'b110110111;
assign micromat[54][66] = 9'b101101101;
assign micromat[54][67] = 9'b100000000;
assign micromat[54][68] = 9'b100000000;
assign micromat[54][69] = 9'b111111111;
assign micromat[54][70] = 9'b111111111;
assign micromat[54][71] = 9'b111111111;
assign micromat[54][72] = 9'b111111111;
assign micromat[54][73] = 9'b110110111;
assign micromat[54][74] = 9'b100100100;
assign micromat[54][75] = 9'b100100100;
assign micromat[54][76] = 9'b100100100;
assign micromat[54][77] = 9'b100100100;
assign micromat[54][78] = 9'b101001001;
assign micromat[54][79] = 9'b111111111;
assign micromat[54][80] = 9'b111111111;
assign micromat[54][81] = 9'b110110111;
assign micromat[54][82] = 9'b110111111;
assign micromat[54][83] = 9'b101001001;
assign micromat[54][84] = 9'b100000000;
assign micromat[54][85] = 9'b100100100;
assign micromat[54][86] = 9'b111111111;
assign micromat[54][87] = 9'b111111111;
assign micromat[54][88] = 9'b111111111;
assign micromat[54][89] = 9'b111111111;
assign micromat[54][90] = 9'b111111111;
assign micromat[54][91] = 9'b111111111;
assign micromat[54][92] = 9'b111111111;
assign micromat[54][93] = 9'b111111111;
assign micromat[54][94] = 9'b111111111;
assign micromat[54][95] = 9'b111111111;
assign micromat[54][96] = 9'b111111111;
assign micromat[54][97] = 9'b111111111;
assign micromat[54][98] = 9'b111111111;
assign micromat[54][99] = 9'b111111111;
assign micromat[55][0] = 9'b111111111;
assign micromat[55][1] = 9'b111111111;
assign micromat[55][2] = 9'b111111111;
assign micromat[55][3] = 9'b111111111;
assign micromat[55][4] = 9'b111111111;
assign micromat[55][5] = 9'b111111111;
assign micromat[55][6] = 9'b111111111;
assign micromat[55][7] = 9'b111111111;
assign micromat[55][8] = 9'b111111111;
assign micromat[55][9] = 9'b111111111;
assign micromat[55][10] = 9'b111111111;
assign micromat[55][11] = 9'b111111111;
assign micromat[55][12] = 9'b111111111;
assign micromat[55][13] = 9'b111111111;
assign micromat[55][14] = 9'b100100100;
assign micromat[55][15] = 9'b100000000;
assign micromat[55][16] = 9'b101101101;
assign micromat[55][17] = 9'b111111111;
assign micromat[55][18] = 9'b111111111;
assign micromat[55][19] = 9'b111111111;
assign micromat[55][20] = 9'b111111111;
assign micromat[55][21] = 9'b100101000;
assign micromat[55][22] = 9'b100000000;
assign micromat[55][23] = 9'b100100100;
assign micromat[55][24] = 9'b101101101;
assign micromat[55][25] = 9'b101101101;
assign micromat[55][26] = 9'b101101101;
assign micromat[55][27] = 9'b101101101;
assign micromat[55][28] = 9'b101101101;
assign micromat[55][29] = 9'b101101101;
assign micromat[55][30] = 9'b101101101;
assign micromat[55][31] = 9'b101101101;
assign micromat[55][32] = 9'b101101101;
assign micromat[55][33] = 9'b101101101;
assign micromat[55][34] = 9'b101101101;
assign micromat[55][35] = 9'b101101101;
assign micromat[55][36] = 9'b101101101;
assign micromat[55][37] = 9'b101101101;
assign micromat[55][38] = 9'b101101101;
assign micromat[55][39] = 9'b101101101;
assign micromat[55][40] = 9'b101101101;
assign micromat[55][41] = 9'b101101101;
assign micromat[55][42] = 9'b101101101;
assign micromat[55][43] = 9'b101101101;
assign micromat[55][44] = 9'b101101101;
assign micromat[55][45] = 9'b101101101;
assign micromat[55][46] = 9'b101101101;
assign micromat[55][47] = 9'b101101101;
assign micromat[55][48] = 9'b101101101;
assign micromat[55][49] = 9'b101101101;
assign micromat[55][50] = 9'b101101101;
assign micromat[55][51] = 9'b101101101;
assign micromat[55][52] = 9'b101101101;
assign micromat[55][53] = 9'b101101101;
assign micromat[55][54] = 9'b101101101;
assign micromat[55][55] = 9'b101101101;
assign micromat[55][56] = 9'b101101101;
assign micromat[55][57] = 9'b110010001;
assign micromat[55][58] = 9'b110110110;
assign micromat[55][59] = 9'b101001001;
assign micromat[55][60] = 9'b100000000;
assign micromat[55][61] = 9'b100000000;
assign micromat[55][62] = 9'b110111111;
assign micromat[55][63] = 9'b111111111;
assign micromat[55][64] = 9'b110110111;
assign micromat[55][65] = 9'b110110111;
assign micromat[55][66] = 9'b101101101;
assign micromat[55][67] = 9'b100000000;
assign micromat[55][68] = 9'b100000000;
assign micromat[55][69] = 9'b111111111;
assign micromat[55][70] = 9'b111111111;
assign micromat[55][71] = 9'b111111111;
assign micromat[55][72] = 9'b111111111;
assign micromat[55][73] = 9'b111111111;
assign micromat[55][74] = 9'b111111111;
assign micromat[55][75] = 9'b111111111;
assign micromat[55][76] = 9'b111111111;
assign micromat[55][77] = 9'b111111111;
assign micromat[55][78] = 9'b111111111;
assign micromat[55][79] = 9'b111111111;
assign micromat[55][80] = 9'b111111111;
assign micromat[55][81] = 9'b110110111;
assign micromat[55][82] = 9'b110111111;
assign micromat[55][83] = 9'b101001001;
assign micromat[55][84] = 9'b100000000;
assign micromat[55][85] = 9'b100100100;
assign micromat[55][86] = 9'b111111111;
assign micromat[55][87] = 9'b111111111;
assign micromat[55][88] = 9'b111111111;
assign micromat[55][89] = 9'b111111111;
assign micromat[55][90] = 9'b111111111;
assign micromat[55][91] = 9'b111111111;
assign micromat[55][92] = 9'b111111111;
assign micromat[55][93] = 9'b111111111;
assign micromat[55][94] = 9'b111111111;
assign micromat[55][95] = 9'b111111111;
assign micromat[55][96] = 9'b111111111;
assign micromat[55][97] = 9'b111111111;
assign micromat[55][98] = 9'b111111111;
assign micromat[55][99] = 9'b111111111;
assign micromat[56][0] = 9'b111111111;
assign micromat[56][1] = 9'b111111111;
assign micromat[56][2] = 9'b111111111;
assign micromat[56][3] = 9'b111111111;
assign micromat[56][4] = 9'b111111111;
assign micromat[56][5] = 9'b111111111;
assign micromat[56][6] = 9'b111111111;
assign micromat[56][7] = 9'b111111111;
assign micromat[56][8] = 9'b111111111;
assign micromat[56][9] = 9'b111111111;
assign micromat[56][10] = 9'b111111111;
assign micromat[56][11] = 9'b111111111;
assign micromat[56][12] = 9'b111111111;
assign micromat[56][13] = 9'b111111111;
assign micromat[56][14] = 9'b100100100;
assign micromat[56][15] = 9'b100000000;
assign micromat[56][16] = 9'b101101101;
assign micromat[56][17] = 9'b111111111;
assign micromat[56][18] = 9'b111111111;
assign micromat[56][19] = 9'b111111111;
assign micromat[56][20] = 9'b111111111;
assign micromat[56][21] = 9'b100101000;
assign micromat[56][22] = 9'b100000000;
assign micromat[56][23] = 9'b100100100;
assign micromat[56][24] = 9'b101101101;
assign micromat[56][25] = 9'b101101101;
assign micromat[56][26] = 9'b101101101;
assign micromat[56][27] = 9'b101101101;
assign micromat[56][28] = 9'b101101101;
assign micromat[56][29] = 9'b101101101;
assign micromat[56][30] = 9'b101101101;
assign micromat[56][31] = 9'b101101101;
assign micromat[56][32] = 9'b101101101;
assign micromat[56][33] = 9'b101101101;
assign micromat[56][34] = 9'b101101101;
assign micromat[56][35] = 9'b101101101;
assign micromat[56][36] = 9'b101101101;
assign micromat[56][37] = 9'b101101101;
assign micromat[56][38] = 9'b101101101;
assign micromat[56][39] = 9'b101101101;
assign micromat[56][40] = 9'b101101101;
assign micromat[56][41] = 9'b101101101;
assign micromat[56][42] = 9'b101101101;
assign micromat[56][43] = 9'b101101101;
assign micromat[56][44] = 9'b101101101;
assign micromat[56][45] = 9'b101101101;
assign micromat[56][46] = 9'b101101101;
assign micromat[56][47] = 9'b101101101;
assign micromat[56][48] = 9'b101101101;
assign micromat[56][49] = 9'b101101101;
assign micromat[56][50] = 9'b101101101;
assign micromat[56][51] = 9'b101101101;
assign micromat[56][52] = 9'b101101101;
assign micromat[56][53] = 9'b101101101;
assign micromat[56][54] = 9'b101101101;
assign micromat[56][55] = 9'b101101101;
assign micromat[56][56] = 9'b101101101;
assign micromat[56][57] = 9'b110010001;
assign micromat[56][58] = 9'b110110110;
assign micromat[56][59] = 9'b101001001;
assign micromat[56][60] = 9'b100000000;
assign micromat[56][61] = 9'b100000000;
assign micromat[56][62] = 9'b110111111;
assign micromat[56][63] = 9'b111111111;
assign micromat[56][64] = 9'b110110111;
assign micromat[56][65] = 9'b110110111;
assign micromat[56][66] = 9'b101101101;
assign micromat[56][67] = 9'b100000000;
assign micromat[56][68] = 9'b100000000;
assign micromat[56][69] = 9'b111111111;
assign micromat[56][70] = 9'b111111111;
assign micromat[56][71] = 9'b111111111;
assign micromat[56][72] = 9'b111111111;
assign micromat[56][73] = 9'b111111111;
assign micromat[56][74] = 9'b111111111;
assign micromat[56][75] = 9'b111111111;
assign micromat[56][76] = 9'b111111111;
assign micromat[56][77] = 9'b111111111;
assign micromat[56][78] = 9'b111111111;
assign micromat[56][79] = 9'b111111111;
assign micromat[56][80] = 9'b111111111;
assign micromat[56][81] = 9'b110110111;
assign micromat[56][82] = 9'b110111111;
assign micromat[56][83] = 9'b101001001;
assign micromat[56][84] = 9'b100000000;
assign micromat[56][85] = 9'b100100100;
assign micromat[56][86] = 9'b111111111;
assign micromat[56][87] = 9'b111111111;
assign micromat[56][88] = 9'b111111111;
assign micromat[56][89] = 9'b111111111;
assign micromat[56][90] = 9'b111111111;
assign micromat[56][91] = 9'b111111111;
assign micromat[56][92] = 9'b111111111;
assign micromat[56][93] = 9'b111111111;
assign micromat[56][94] = 9'b111111111;
assign micromat[56][95] = 9'b111111111;
assign micromat[56][96] = 9'b111111111;
assign micromat[56][97] = 9'b111111111;
assign micromat[56][98] = 9'b111111111;
assign micromat[56][99] = 9'b111111111;
assign micromat[57][0] = 9'b111111111;
assign micromat[57][1] = 9'b111111111;
assign micromat[57][2] = 9'b111111111;
assign micromat[57][3] = 9'b111111111;
assign micromat[57][4] = 9'b111111111;
assign micromat[57][5] = 9'b111111111;
assign micromat[57][6] = 9'b111111111;
assign micromat[57][7] = 9'b111111111;
assign micromat[57][8] = 9'b111111111;
assign micromat[57][9] = 9'b111111111;
assign micromat[57][10] = 9'b111111111;
assign micromat[57][11] = 9'b111111111;
assign micromat[57][12] = 9'b111111111;
assign micromat[57][13] = 9'b111111111;
assign micromat[57][14] = 9'b100100100;
assign micromat[57][15] = 9'b100000000;
assign micromat[57][16] = 9'b101101101;
assign micromat[57][17] = 9'b111111111;
assign micromat[57][18] = 9'b111111111;
assign micromat[57][19] = 9'b111111111;
assign micromat[57][20] = 9'b111111111;
assign micromat[57][21] = 9'b100101000;
assign micromat[57][22] = 9'b100000000;
assign micromat[57][23] = 9'b100100100;
assign micromat[57][24] = 9'b101101101;
assign micromat[57][25] = 9'b101101101;
assign micromat[57][26] = 9'b100100100;
assign micromat[57][27] = 9'b100000000;
assign micromat[57][28] = 9'b100000000;
assign micromat[57][29] = 9'b100000000;
assign micromat[57][30] = 9'b100000000;
assign micromat[57][31] = 9'b100000000;
assign micromat[57][32] = 9'b100000000;
assign micromat[57][33] = 9'b100000000;
assign micromat[57][34] = 9'b100000000;
assign micromat[57][35] = 9'b100000000;
assign micromat[57][36] = 9'b100000000;
assign micromat[57][37] = 9'b100000000;
assign micromat[57][38] = 9'b100000000;
assign micromat[57][39] = 9'b100000000;
assign micromat[57][40] = 9'b100000000;
assign micromat[57][41] = 9'b100000000;
assign micromat[57][42] = 9'b100000000;
assign micromat[57][43] = 9'b100000000;
assign micromat[57][44] = 9'b100000000;
assign micromat[57][45] = 9'b100000000;
assign micromat[57][46] = 9'b100000000;
assign micromat[57][47] = 9'b100000000;
assign micromat[57][48] = 9'b100000000;
assign micromat[57][49] = 9'b100000000;
assign micromat[57][50] = 9'b100000000;
assign micromat[57][51] = 9'b100000000;
assign micromat[57][52] = 9'b100000000;
assign micromat[57][53] = 9'b100000000;
assign micromat[57][54] = 9'b100000000;
assign micromat[57][55] = 9'b100000000;
assign micromat[57][56] = 9'b100000000;
assign micromat[57][57] = 9'b101101101;
assign micromat[57][58] = 9'b110110110;
assign micromat[57][59] = 9'b101001001;
assign micromat[57][60] = 9'b100000000;
assign micromat[57][61] = 9'b100000000;
assign micromat[57][62] = 9'b110111111;
assign micromat[57][63] = 9'b111111111;
assign micromat[57][64] = 9'b110110111;
assign micromat[57][65] = 9'b110110111;
assign micromat[57][66] = 9'b101101101;
assign micromat[57][67] = 9'b100000000;
assign micromat[57][68] = 9'b100000000;
assign micromat[57][69] = 9'b111111111;
assign micromat[57][70] = 9'b111111111;
assign micromat[57][71] = 9'b111111111;
assign micromat[57][72] = 9'b111111111;
assign micromat[57][73] = 9'b110110111;
assign micromat[57][74] = 9'b100100100;
assign micromat[57][75] = 9'b100100100;
assign micromat[57][76] = 9'b100100100;
assign micromat[57][77] = 9'b100100100;
assign micromat[57][78] = 9'b101001001;
assign micromat[57][79] = 9'b111111111;
assign micromat[57][80] = 9'b111111111;
assign micromat[57][81] = 9'b110110111;
assign micromat[57][82] = 9'b110111111;
assign micromat[57][83] = 9'b101001001;
assign micromat[57][84] = 9'b100000000;
assign micromat[57][85] = 9'b100100100;
assign micromat[57][86] = 9'b111111111;
assign micromat[57][87] = 9'b111111111;
assign micromat[57][88] = 9'b111111111;
assign micromat[57][89] = 9'b111111111;
assign micromat[57][90] = 9'b111111111;
assign micromat[57][91] = 9'b111111111;
assign micromat[57][92] = 9'b111111111;
assign micromat[57][93] = 9'b111111111;
assign micromat[57][94] = 9'b111111111;
assign micromat[57][95] = 9'b111111111;
assign micromat[57][96] = 9'b111111111;
assign micromat[57][97] = 9'b111111111;
assign micromat[57][98] = 9'b111111111;
assign micromat[57][99] = 9'b111111111;
assign micromat[58][0] = 9'b111111111;
assign micromat[58][1] = 9'b111111111;
assign micromat[58][2] = 9'b111111111;
assign micromat[58][3] = 9'b111111111;
assign micromat[58][4] = 9'b111111111;
assign micromat[58][5] = 9'b111111111;
assign micromat[58][6] = 9'b111111111;
assign micromat[58][7] = 9'b111111111;
assign micromat[58][8] = 9'b111111111;
assign micromat[58][9] = 9'b111111111;
assign micromat[58][10] = 9'b111111111;
assign micromat[58][11] = 9'b111111111;
assign micromat[58][12] = 9'b111111111;
assign micromat[58][13] = 9'b111111111;
assign micromat[58][14] = 9'b100100100;
assign micromat[58][15] = 9'b100000000;
assign micromat[58][16] = 9'b101101101;
assign micromat[58][17] = 9'b111111111;
assign micromat[58][18] = 9'b111111111;
assign micromat[58][19] = 9'b111111111;
assign micromat[58][20] = 9'b111111111;
assign micromat[58][21] = 9'b100101000;
assign micromat[58][22] = 9'b100000000;
assign micromat[58][23] = 9'b100100100;
assign micromat[58][24] = 9'b101101101;
assign micromat[58][25] = 9'b101101101;
assign micromat[58][26] = 9'b100000000;
assign micromat[58][27] = 9'b100000000;
assign micromat[58][28] = 9'b100000000;
assign micromat[58][29] = 9'b100000000;
assign micromat[58][30] = 9'b100000000;
assign micromat[58][31] = 9'b100000000;
assign micromat[58][32] = 9'b100000000;
assign micromat[58][33] = 9'b100000000;
assign micromat[58][34] = 9'b100000000;
assign micromat[58][35] = 9'b100000000;
assign micromat[58][36] = 9'b100000000;
assign micromat[58][37] = 9'b100000000;
assign micromat[58][38] = 9'b100000000;
assign micromat[58][39] = 9'b100000000;
assign micromat[58][40] = 9'b100000000;
assign micromat[58][41] = 9'b100000000;
assign micromat[58][42] = 9'b100000000;
assign micromat[58][43] = 9'b100000000;
assign micromat[58][44] = 9'b100000000;
assign micromat[58][45] = 9'b100000000;
assign micromat[58][46] = 9'b100000000;
assign micromat[58][47] = 9'b100000000;
assign micromat[58][48] = 9'b100000000;
assign micromat[58][49] = 9'b100000000;
assign micromat[58][50] = 9'b100000000;
assign micromat[58][51] = 9'b100000000;
assign micromat[58][52] = 9'b100000000;
assign micromat[58][53] = 9'b100000000;
assign micromat[58][54] = 9'b100000000;
assign micromat[58][55] = 9'b100000000;
assign micromat[58][56] = 9'b100000000;
assign micromat[58][57] = 9'b101101101;
assign micromat[58][58] = 9'b110110110;
assign micromat[58][59] = 9'b101001001;
assign micromat[58][60] = 9'b100000000;
assign micromat[58][61] = 9'b100000000;
assign micromat[58][62] = 9'b110111111;
assign micromat[58][63] = 9'b111111111;
assign micromat[58][64] = 9'b110110111;
assign micromat[58][65] = 9'b110110111;
assign micromat[58][66] = 9'b101101101;
assign micromat[58][67] = 9'b100000000;
assign micromat[58][68] = 9'b100000000;
assign micromat[58][69] = 9'b111111111;
assign micromat[58][70] = 9'b111111111;
assign micromat[58][71] = 9'b111111111;
assign micromat[58][72] = 9'b111111111;
assign micromat[58][73] = 9'b110111111;
assign micromat[58][74] = 9'b100000000;
assign micromat[58][75] = 9'b100000000;
assign micromat[58][76] = 9'b100000000;
assign micromat[58][77] = 9'b100000000;
assign micromat[58][78] = 9'b100100100;
assign micromat[58][79] = 9'b111111111;
assign micromat[58][80] = 9'b111111111;
assign micromat[58][81] = 9'b110110111;
assign micromat[58][82] = 9'b110111111;
assign micromat[58][83] = 9'b101001001;
assign micromat[58][84] = 9'b100000000;
assign micromat[58][85] = 9'b100100100;
assign micromat[58][86] = 9'b111111111;
assign micromat[58][87] = 9'b111111111;
assign micromat[58][88] = 9'b111111111;
assign micromat[58][89] = 9'b111111111;
assign micromat[58][90] = 9'b111111111;
assign micromat[58][91] = 9'b111111111;
assign micromat[58][92] = 9'b111111111;
assign micromat[58][93] = 9'b111111111;
assign micromat[58][94] = 9'b111111111;
assign micromat[58][95] = 9'b111111111;
assign micromat[58][96] = 9'b111111111;
assign micromat[58][97] = 9'b111111111;
assign micromat[58][98] = 9'b111111111;
assign micromat[58][99] = 9'b111111111;
assign micromat[59][0] = 9'b111111111;
assign micromat[59][1] = 9'b111111111;
assign micromat[59][2] = 9'b111111111;
assign micromat[59][3] = 9'b111111111;
assign micromat[59][4] = 9'b111111111;
assign micromat[59][5] = 9'b111111111;
assign micromat[59][6] = 9'b111111111;
assign micromat[59][7] = 9'b111111111;
assign micromat[59][8] = 9'b111111111;
assign micromat[59][9] = 9'b111111111;
assign micromat[59][10] = 9'b111111111;
assign micromat[59][11] = 9'b111111111;
assign micromat[59][12] = 9'b111111111;
assign micromat[59][13] = 9'b111111111;
assign micromat[59][14] = 9'b100100100;
assign micromat[59][15] = 9'b100000000;
assign micromat[59][16] = 9'b101101101;
assign micromat[59][17] = 9'b111111111;
assign micromat[59][18] = 9'b111111111;
assign micromat[59][19] = 9'b111111111;
assign micromat[59][20] = 9'b111111111;
assign micromat[59][21] = 9'b100101000;
assign micromat[59][22] = 9'b100000000;
assign micromat[59][23] = 9'b100100100;
assign micromat[59][24] = 9'b101101101;
assign micromat[59][25] = 9'b101101101;
assign micromat[59][26] = 9'b101001001;
assign micromat[59][27] = 9'b101001000;
assign micromat[59][28] = 9'b101001000;
assign micromat[59][29] = 9'b101001000;
assign micromat[59][30] = 9'b101001000;
assign micromat[59][31] = 9'b101001000;
assign micromat[59][32] = 9'b101001000;
assign micromat[59][33] = 9'b101001000;
assign micromat[59][34] = 9'b101001000;
assign micromat[59][35] = 9'b101001000;
assign micromat[59][36] = 9'b101001000;
assign micromat[59][37] = 9'b101001000;
assign micromat[59][38] = 9'b101001000;
assign micromat[59][39] = 9'b101001000;
assign micromat[59][40] = 9'b101001000;
assign micromat[59][41] = 9'b101001000;
assign micromat[59][42] = 9'b101001000;
assign micromat[59][43] = 9'b101001000;
assign micromat[59][44] = 9'b101001000;
assign micromat[59][45] = 9'b101001000;
assign micromat[59][46] = 9'b101001000;
assign micromat[59][47] = 9'b101001000;
assign micromat[59][48] = 9'b101001000;
assign micromat[59][49] = 9'b101001000;
assign micromat[59][50] = 9'b101001000;
assign micromat[59][51] = 9'b101001000;
assign micromat[59][52] = 9'b101001000;
assign micromat[59][53] = 9'b101001000;
assign micromat[59][54] = 9'b101001000;
assign micromat[59][55] = 9'b101001000;
assign micromat[59][56] = 9'b101001000;
assign micromat[59][57] = 9'b110010001;
assign micromat[59][58] = 9'b110110110;
assign micromat[59][59] = 9'b101001001;
assign micromat[59][60] = 9'b100000000;
assign micromat[59][61] = 9'b100000000;
assign micromat[59][62] = 9'b110111111;
assign micromat[59][63] = 9'b111111111;
assign micromat[59][64] = 9'b110110111;
assign micromat[59][65] = 9'b110110111;
assign micromat[59][66] = 9'b101101101;
assign micromat[59][67] = 9'b100000000;
assign micromat[59][68] = 9'b100000000;
assign micromat[59][69] = 9'b111111111;
assign micromat[59][70] = 9'b111111111;
assign micromat[59][71] = 9'b110110110;
assign micromat[59][72] = 9'b101101101;
assign micromat[59][73] = 9'b101101101;
assign micromat[59][74] = 9'b101101101;
assign micromat[59][75] = 9'b101101101;
assign micromat[59][76] = 9'b101001001;
assign micromat[59][77] = 9'b101001001;
assign micromat[59][78] = 9'b101001101;
assign micromat[59][79] = 9'b101101101;
assign micromat[59][80] = 9'b101101101;
assign micromat[59][81] = 9'b110010010;
assign micromat[59][82] = 9'b110111111;
assign micromat[59][83] = 9'b101001001;
assign micromat[59][84] = 9'b100000000;
assign micromat[59][85] = 9'b100100100;
assign micromat[59][86] = 9'b111111111;
assign micromat[59][87] = 9'b111111111;
assign micromat[59][88] = 9'b111111111;
assign micromat[59][89] = 9'b111111111;
assign micromat[59][90] = 9'b111111111;
assign micromat[59][91] = 9'b111111111;
assign micromat[59][92] = 9'b111111111;
assign micromat[59][93] = 9'b111111111;
assign micromat[59][94] = 9'b111111111;
assign micromat[59][95] = 9'b111111111;
assign micromat[59][96] = 9'b111111111;
assign micromat[59][97] = 9'b111111111;
assign micromat[59][98] = 9'b111111111;
assign micromat[59][99] = 9'b111111111;
assign micromat[60][0] = 9'b111111111;
assign micromat[60][1] = 9'b111111111;
assign micromat[60][2] = 9'b111111111;
assign micromat[60][3] = 9'b111111111;
assign micromat[60][4] = 9'b111111111;
assign micromat[60][5] = 9'b111111111;
assign micromat[60][6] = 9'b111111111;
assign micromat[60][7] = 9'b111111111;
assign micromat[60][8] = 9'b111111111;
assign micromat[60][9] = 9'b111111111;
assign micromat[60][10] = 9'b111111111;
assign micromat[60][11] = 9'b111111111;
assign micromat[60][12] = 9'b111111111;
assign micromat[60][13] = 9'b111111111;
assign micromat[60][14] = 9'b100100100;
assign micromat[60][15] = 9'b100000000;
assign micromat[60][16] = 9'b101101101;
assign micromat[60][17] = 9'b111111111;
assign micromat[60][18] = 9'b111111111;
assign micromat[60][19] = 9'b111111111;
assign micromat[60][20] = 9'b111111111;
assign micromat[60][21] = 9'b100101000;
assign micromat[60][22] = 9'b100000000;
assign micromat[60][23] = 9'b100100100;
assign micromat[60][24] = 9'b101101101;
assign micromat[60][25] = 9'b101101101;
assign micromat[60][26] = 9'b110010010;
assign micromat[60][27] = 9'b110110110;
assign micromat[60][28] = 9'b110110110;
assign micromat[60][29] = 9'b110110110;
assign micromat[60][30] = 9'b110110110;
assign micromat[60][31] = 9'b110110110;
assign micromat[60][32] = 9'b110110110;
assign micromat[60][33] = 9'b110110110;
assign micromat[60][34] = 9'b110110110;
assign micromat[60][35] = 9'b110110110;
assign micromat[60][36] = 9'b110110110;
assign micromat[60][37] = 9'b110110110;
assign micromat[60][38] = 9'b110110110;
assign micromat[60][39] = 9'b110110110;
assign micromat[60][40] = 9'b110110110;
assign micromat[60][41] = 9'b110110110;
assign micromat[60][42] = 9'b110110110;
assign micromat[60][43] = 9'b110110110;
assign micromat[60][44] = 9'b110110110;
assign micromat[60][45] = 9'b110110110;
assign micromat[60][46] = 9'b110110110;
assign micromat[60][47] = 9'b110110110;
assign micromat[60][48] = 9'b110110110;
assign micromat[60][49] = 9'b110110110;
assign micromat[60][50] = 9'b110110110;
assign micromat[60][51] = 9'b110110110;
assign micromat[60][52] = 9'b110110110;
assign micromat[60][53] = 9'b110110110;
assign micromat[60][54] = 9'b110110110;
assign micromat[60][55] = 9'b110110110;
assign micromat[60][56] = 9'b110110110;
assign micromat[60][57] = 9'b110010010;
assign micromat[60][58] = 9'b110110110;
assign micromat[60][59] = 9'b101001001;
assign micromat[60][60] = 9'b100000000;
assign micromat[60][61] = 9'b100000000;
assign micromat[60][62] = 9'b110111111;
assign micromat[60][63] = 9'b111111111;
assign micromat[60][64] = 9'b110110111;
assign micromat[60][65] = 9'b110110111;
assign micromat[60][66] = 9'b101101101;
assign micromat[60][67] = 9'b100000000;
assign micromat[60][68] = 9'b100000000;
assign micromat[60][69] = 9'b111111111;
assign micromat[60][70] = 9'b111111111;
assign micromat[60][71] = 9'b101101101;
assign micromat[60][72] = 9'b100000000;
assign micromat[60][73] = 9'b100000000;
assign micromat[60][74] = 9'b111111111;
assign micromat[60][75] = 9'b111111111;
assign micromat[60][76] = 9'b111111111;
assign micromat[60][77] = 9'b111111111;
assign micromat[60][78] = 9'b110010010;
assign micromat[60][79] = 9'b100000000;
assign micromat[60][80] = 9'b100000000;
assign micromat[60][81] = 9'b110010010;
assign micromat[60][82] = 9'b111111111;
assign micromat[60][83] = 9'b101001001;
assign micromat[60][84] = 9'b100000000;
assign micromat[60][85] = 9'b100100100;
assign micromat[60][86] = 9'b111111111;
assign micromat[60][87] = 9'b111111111;
assign micromat[60][88] = 9'b111111111;
assign micromat[60][89] = 9'b111111111;
assign micromat[60][90] = 9'b111111111;
assign micromat[60][91] = 9'b111111111;
assign micromat[60][92] = 9'b111111111;
assign micromat[60][93] = 9'b111111111;
assign micromat[60][94] = 9'b111111111;
assign micromat[60][95] = 9'b111111111;
assign micromat[60][96] = 9'b111111111;
assign micromat[60][97] = 9'b111111111;
assign micromat[60][98] = 9'b111111111;
assign micromat[60][99] = 9'b111111111;
assign micromat[61][0] = 9'b111111111;
assign micromat[61][1] = 9'b111111111;
assign micromat[61][2] = 9'b111111111;
assign micromat[61][3] = 9'b111111111;
assign micromat[61][4] = 9'b111111111;
assign micromat[61][5] = 9'b111111111;
assign micromat[61][6] = 9'b111111111;
assign micromat[61][7] = 9'b111111111;
assign micromat[61][8] = 9'b111111111;
assign micromat[61][9] = 9'b111111111;
assign micromat[61][10] = 9'b111111111;
assign micromat[61][11] = 9'b111111111;
assign micromat[61][12] = 9'b111111111;
assign micromat[61][13] = 9'b111111111;
assign micromat[61][14] = 9'b100100100;
assign micromat[61][15] = 9'b100000000;
assign micromat[61][16] = 9'b101101101;
assign micromat[61][17] = 9'b111111111;
assign micromat[61][18] = 9'b111111111;
assign micromat[61][19] = 9'b111111111;
assign micromat[61][20] = 9'b111111111;
assign micromat[61][21] = 9'b100101000;
assign micromat[61][22] = 9'b100000000;
assign micromat[61][23] = 9'b100100100;
assign micromat[61][24] = 9'b101101101;
assign micromat[61][25] = 9'b101101101;
assign micromat[61][26] = 9'b110010001;
assign micromat[61][27] = 9'b110010001;
assign micromat[61][28] = 9'b110010001;
assign micromat[61][29] = 9'b110010001;
assign micromat[61][30] = 9'b110010001;
assign micromat[61][31] = 9'b110010001;
assign micromat[61][32] = 9'b110010001;
assign micromat[61][33] = 9'b110010001;
assign micromat[61][34] = 9'b110010001;
assign micromat[61][35] = 9'b110010001;
assign micromat[61][36] = 9'b110010001;
assign micromat[61][37] = 9'b110010001;
assign micromat[61][38] = 9'b110010001;
assign micromat[61][39] = 9'b110010001;
assign micromat[61][40] = 9'b110010001;
assign micromat[61][41] = 9'b110010001;
assign micromat[61][42] = 9'b110010001;
assign micromat[61][43] = 9'b110010001;
assign micromat[61][44] = 9'b110010001;
assign micromat[61][45] = 9'b110010001;
assign micromat[61][46] = 9'b110010001;
assign micromat[61][47] = 9'b110010001;
assign micromat[61][48] = 9'b110010001;
assign micromat[61][49] = 9'b110010001;
assign micromat[61][50] = 9'b110010001;
assign micromat[61][51] = 9'b110010001;
assign micromat[61][52] = 9'b110010001;
assign micromat[61][53] = 9'b110010001;
assign micromat[61][54] = 9'b110010001;
assign micromat[61][55] = 9'b110010001;
assign micromat[61][56] = 9'b110010001;
assign micromat[61][57] = 9'b110010001;
assign micromat[61][58] = 9'b110010001;
assign micromat[61][59] = 9'b101001001;
assign micromat[61][60] = 9'b100000000;
assign micromat[61][61] = 9'b100000000;
assign micromat[61][62] = 9'b110111111;
assign micromat[61][63] = 9'b111111111;
assign micromat[61][64] = 9'b110110111;
assign micromat[61][65] = 9'b110110111;
assign micromat[61][66] = 9'b101101101;
assign micromat[61][67] = 9'b100000000;
assign micromat[61][68] = 9'b100000000;
assign micromat[61][69] = 9'b111111111;
assign micromat[61][70] = 9'b111111111;
assign micromat[61][71] = 9'b101101101;
assign micromat[61][72] = 9'b100000000;
assign micromat[61][73] = 9'b100000100;
assign micromat[61][74] = 9'b111111111;
assign micromat[61][75] = 9'b111111111;
assign micromat[61][76] = 9'b111111111;
assign micromat[61][77] = 9'b111111111;
assign micromat[61][78] = 9'b110010001;
assign micromat[61][79] = 9'b100000000;
assign micromat[61][80] = 9'b100000000;
assign micromat[61][81] = 9'b110010010;
assign micromat[61][82] = 9'b111111111;
assign micromat[61][83] = 9'b101001001;
assign micromat[61][84] = 9'b100000000;
assign micromat[61][85] = 9'b100100100;
assign micromat[61][86] = 9'b111111111;
assign micromat[61][87] = 9'b111111111;
assign micromat[61][88] = 9'b111111111;
assign micromat[61][89] = 9'b111111111;
assign micromat[61][90] = 9'b111111111;
assign micromat[61][91] = 9'b111111111;
assign micromat[61][92] = 9'b111111111;
assign micromat[61][93] = 9'b111111111;
assign micromat[61][94] = 9'b111111111;
assign micromat[61][95] = 9'b111111111;
assign micromat[61][96] = 9'b111111111;
assign micromat[61][97] = 9'b111111111;
assign micromat[61][98] = 9'b111111111;
assign micromat[61][99] = 9'b111111111;
assign micromat[62][0] = 9'b111111111;
assign micromat[62][1] = 9'b111111111;
assign micromat[62][2] = 9'b111111111;
assign micromat[62][3] = 9'b111111111;
assign micromat[62][4] = 9'b111111111;
assign micromat[62][5] = 9'b111111111;
assign micromat[62][6] = 9'b111111111;
assign micromat[62][7] = 9'b111111111;
assign micromat[62][8] = 9'b111111111;
assign micromat[62][9] = 9'b111111111;
assign micromat[62][10] = 9'b111111111;
assign micromat[62][11] = 9'b111111111;
assign micromat[62][12] = 9'b111111111;
assign micromat[62][13] = 9'b111111111;
assign micromat[62][14] = 9'b100100100;
assign micromat[62][15] = 9'b100000000;
assign micromat[62][16] = 9'b101101101;
assign micromat[62][17] = 9'b111111111;
assign micromat[62][18] = 9'b111111111;
assign micromat[62][19] = 9'b111111111;
assign micromat[62][20] = 9'b111111111;
assign micromat[62][21] = 9'b100101000;
assign micromat[62][22] = 9'b100000000;
assign micromat[62][23] = 9'b100000000;
assign micromat[62][24] = 9'b100000000;
assign micromat[62][25] = 9'b100000000;
assign micromat[62][26] = 9'b100000000;
assign micromat[62][27] = 9'b100000000;
assign micromat[62][28] = 9'b100000000;
assign micromat[62][29] = 9'b100000000;
assign micromat[62][30] = 9'b100000000;
assign micromat[62][31] = 9'b100000000;
assign micromat[62][32] = 9'b100000000;
assign micromat[62][33] = 9'b100000000;
assign micromat[62][34] = 9'b100000000;
assign micromat[62][35] = 9'b100000000;
assign micromat[62][36] = 9'b100000000;
assign micromat[62][37] = 9'b100000000;
assign micromat[62][38] = 9'b100000000;
assign micromat[62][39] = 9'b100000000;
assign micromat[62][40] = 9'b100000000;
assign micromat[62][41] = 9'b100000000;
assign micromat[62][42] = 9'b100000000;
assign micromat[62][43] = 9'b100000000;
assign micromat[62][44] = 9'b100000000;
assign micromat[62][45] = 9'b100000000;
assign micromat[62][46] = 9'b100000000;
assign micromat[62][47] = 9'b100000000;
assign micromat[62][48] = 9'b100000000;
assign micromat[62][49] = 9'b100000000;
assign micromat[62][50] = 9'b100000000;
assign micromat[62][51] = 9'b100000000;
assign micromat[62][52] = 9'b100000000;
assign micromat[62][53] = 9'b100000000;
assign micromat[62][54] = 9'b100000000;
assign micromat[62][55] = 9'b100000000;
assign micromat[62][56] = 9'b100000000;
assign micromat[62][57] = 9'b100000000;
assign micromat[62][58] = 9'b100000000;
assign micromat[62][59] = 9'b100000000;
assign micromat[62][60] = 9'b100000000;
assign micromat[62][61] = 9'b100000000;
assign micromat[62][62] = 9'b110111111;
assign micromat[62][63] = 9'b111111111;
assign micromat[62][64] = 9'b110110111;
assign micromat[62][65] = 9'b110110111;
assign micromat[62][66] = 9'b101101101;
assign micromat[62][67] = 9'b100000000;
assign micromat[62][68] = 9'b100000000;
assign micromat[62][69] = 9'b111111111;
assign micromat[62][70] = 9'b111111111;
assign micromat[62][71] = 9'b101101101;
assign micromat[62][72] = 9'b100000000;
assign micromat[62][73] = 9'b100000000;
assign micromat[62][74] = 9'b111111111;
assign micromat[62][75] = 9'b111111111;
assign micromat[62][76] = 9'b110110111;
assign micromat[62][77] = 9'b110110111;
assign micromat[62][78] = 9'b101101101;
assign micromat[62][79] = 9'b100000000;
assign micromat[62][80] = 9'b100000000;
assign micromat[62][81] = 9'b110010010;
assign micromat[62][82] = 9'b111111111;
assign micromat[62][83] = 9'b101001001;
assign micromat[62][84] = 9'b100000000;
assign micromat[62][85] = 9'b100100100;
assign micromat[62][86] = 9'b111111111;
assign micromat[62][87] = 9'b111111111;
assign micromat[62][88] = 9'b111111111;
assign micromat[62][89] = 9'b111111111;
assign micromat[62][90] = 9'b111111111;
assign micromat[62][91] = 9'b111111111;
assign micromat[62][92] = 9'b111111111;
assign micromat[62][93] = 9'b111111111;
assign micromat[62][94] = 9'b111111111;
assign micromat[62][95] = 9'b111111111;
assign micromat[62][96] = 9'b111111111;
assign micromat[62][97] = 9'b111111111;
assign micromat[62][98] = 9'b111111111;
assign micromat[62][99] = 9'b111111111;
assign micromat[63][0] = 9'b111111111;
assign micromat[63][1] = 9'b111111111;
assign micromat[63][2] = 9'b111111111;
assign micromat[63][3] = 9'b111111111;
assign micromat[63][4] = 9'b111111111;
assign micromat[63][5] = 9'b111111111;
assign micromat[63][6] = 9'b111111111;
assign micromat[63][7] = 9'b111111111;
assign micromat[63][8] = 9'b111111111;
assign micromat[63][9] = 9'b111111111;
assign micromat[63][10] = 9'b111111111;
assign micromat[63][11] = 9'b111111111;
assign micromat[63][12] = 9'b111111111;
assign micromat[63][13] = 9'b111111111;
assign micromat[63][14] = 9'b100100100;
assign micromat[63][15] = 9'b100000000;
assign micromat[63][16] = 9'b101101101;
assign micromat[63][17] = 9'b111111111;
assign micromat[63][18] = 9'b111111111;
assign micromat[63][19] = 9'b111111111;
assign micromat[63][20] = 9'b111111111;
assign micromat[63][21] = 9'b100100100;
assign micromat[63][22] = 9'b100000000;
assign micromat[63][23] = 9'b100000000;
assign micromat[63][24] = 9'b100000000;
assign micromat[63][25] = 9'b100000000;
assign micromat[63][26] = 9'b100000000;
assign micromat[63][27] = 9'b100000000;
assign micromat[63][28] = 9'b100000000;
assign micromat[63][29] = 9'b100000000;
assign micromat[63][30] = 9'b100000000;
assign micromat[63][31] = 9'b100000000;
assign micromat[63][32] = 9'b100000000;
assign micromat[63][33] = 9'b100000000;
assign micromat[63][34] = 9'b100000000;
assign micromat[63][35] = 9'b100000000;
assign micromat[63][36] = 9'b100000000;
assign micromat[63][37] = 9'b100000000;
assign micromat[63][38] = 9'b100000000;
assign micromat[63][39] = 9'b100000000;
assign micromat[63][40] = 9'b100000000;
assign micromat[63][41] = 9'b100000000;
assign micromat[63][42] = 9'b100000000;
assign micromat[63][43] = 9'b100000000;
assign micromat[63][44] = 9'b100000000;
assign micromat[63][45] = 9'b100000000;
assign micromat[63][46] = 9'b100000000;
assign micromat[63][47] = 9'b100000000;
assign micromat[63][48] = 9'b100000000;
assign micromat[63][49] = 9'b100000000;
assign micromat[63][50] = 9'b100000000;
assign micromat[63][51] = 9'b100000000;
assign micromat[63][52] = 9'b100000000;
assign micromat[63][53] = 9'b100000000;
assign micromat[63][54] = 9'b100000000;
assign micromat[63][55] = 9'b100000000;
assign micromat[63][56] = 9'b100000000;
assign micromat[63][57] = 9'b100000000;
assign micromat[63][58] = 9'b100000000;
assign micromat[63][59] = 9'b100000000;
assign micromat[63][60] = 9'b100000000;
assign micromat[63][61] = 9'b100000000;
assign micromat[63][62] = 9'b110111111;
assign micromat[63][63] = 9'b111111111;
assign micromat[63][64] = 9'b110110111;
assign micromat[63][65] = 9'b110110111;
assign micromat[63][66] = 9'b101101101;
assign micromat[63][67] = 9'b100000000;
assign micromat[63][68] = 9'b100000000;
assign micromat[63][69] = 9'b111111111;
assign micromat[63][70] = 9'b111111111;
assign micromat[63][71] = 9'b101101101;
assign micromat[63][72] = 9'b100000000;
assign micromat[63][73] = 9'b100000000;
assign micromat[63][74] = 9'b111111111;
assign micromat[63][75] = 9'b111111111;
assign micromat[63][76] = 9'b111111111;
assign micromat[63][77] = 9'b111111111;
assign micromat[63][78] = 9'b101101101;
assign micromat[63][79] = 9'b100000000;
assign micromat[63][80] = 9'b100000000;
assign micromat[63][81] = 9'b110010010;
assign micromat[63][82] = 9'b111111111;
assign micromat[63][83] = 9'b101001001;
assign micromat[63][84] = 9'b100000000;
assign micromat[63][85] = 9'b100100100;
assign micromat[63][86] = 9'b111111111;
assign micromat[63][87] = 9'b111111111;
assign micromat[63][88] = 9'b111111111;
assign micromat[63][89] = 9'b111111111;
assign micromat[63][90] = 9'b111111111;
assign micromat[63][91] = 9'b111111111;
assign micromat[63][92] = 9'b111111111;
assign micromat[63][93] = 9'b111111111;
assign micromat[63][94] = 9'b111111111;
assign micromat[63][95] = 9'b111111111;
assign micromat[63][96] = 9'b111111111;
assign micromat[63][97] = 9'b111111111;
assign micromat[63][98] = 9'b111111111;
assign micromat[63][99] = 9'b111111111;
assign micromat[64][0] = 9'b111111111;
assign micromat[64][1] = 9'b111111111;
assign micromat[64][2] = 9'b111111111;
assign micromat[64][3] = 9'b111111111;
assign micromat[64][4] = 9'b111111111;
assign micromat[64][5] = 9'b111111111;
assign micromat[64][6] = 9'b111111111;
assign micromat[64][7] = 9'b111111111;
assign micromat[64][8] = 9'b111111111;
assign micromat[64][9] = 9'b111111111;
assign micromat[64][10] = 9'b111111111;
assign micromat[64][11] = 9'b111111111;
assign micromat[64][12] = 9'b111111111;
assign micromat[64][13] = 9'b111111111;
assign micromat[64][14] = 9'b100100100;
assign micromat[64][15] = 9'b100000000;
assign micromat[64][16] = 9'b101101101;
assign micromat[64][17] = 9'b111111111;
assign micromat[64][18] = 9'b111111111;
assign micromat[64][19] = 9'b111111111;
assign micromat[64][20] = 9'b111111111;
assign micromat[64][21] = 9'b110010010;
assign micromat[64][22] = 9'b101101101;
assign micromat[64][23] = 9'b101110001;
assign micromat[64][24] = 9'b101110001;
assign micromat[64][25] = 9'b101110001;
assign micromat[64][26] = 9'b101110001;
assign micromat[64][27] = 9'b101110001;
assign micromat[64][28] = 9'b101110001;
assign micromat[64][29] = 9'b101110001;
assign micromat[64][30] = 9'b101110001;
assign micromat[64][31] = 9'b101110001;
assign micromat[64][32] = 9'b101110001;
assign micromat[64][33] = 9'b101110001;
assign micromat[64][34] = 9'b101110001;
assign micromat[64][35] = 9'b101110001;
assign micromat[64][36] = 9'b101110001;
assign micromat[64][37] = 9'b101110001;
assign micromat[64][38] = 9'b101110001;
assign micromat[64][39] = 9'b101110001;
assign micromat[64][40] = 9'b101110001;
assign micromat[64][41] = 9'b101110001;
assign micromat[64][42] = 9'b101110001;
assign micromat[64][43] = 9'b101110001;
assign micromat[64][44] = 9'b101110001;
assign micromat[64][45] = 9'b101110001;
assign micromat[64][46] = 9'b101110001;
assign micromat[64][47] = 9'b101110001;
assign micromat[64][48] = 9'b101110001;
assign micromat[64][49] = 9'b101110001;
assign micromat[64][50] = 9'b101110001;
assign micromat[64][51] = 9'b101110001;
assign micromat[64][52] = 9'b101110001;
assign micromat[64][53] = 9'b101110001;
assign micromat[64][54] = 9'b101110001;
assign micromat[64][55] = 9'b101110001;
assign micromat[64][56] = 9'b101110001;
assign micromat[64][57] = 9'b101110001;
assign micromat[64][58] = 9'b101110001;
assign micromat[64][59] = 9'b101110001;
assign micromat[64][60] = 9'b101110001;
assign micromat[64][61] = 9'b101110001;
assign micromat[64][62] = 9'b111111111;
assign micromat[64][63] = 9'b111111111;
assign micromat[64][64] = 9'b110110111;
assign micromat[64][65] = 9'b110110111;
assign micromat[64][66] = 9'b101101101;
assign micromat[64][67] = 9'b100000000;
assign micromat[64][68] = 9'b100000000;
assign micromat[64][69] = 9'b111111111;
assign micromat[64][70] = 9'b111111111;
assign micromat[64][71] = 9'b110110111;
assign micromat[64][72] = 9'b101110001;
assign micromat[64][73] = 9'b101101101;
assign micromat[64][74] = 9'b101001001;
assign micromat[64][75] = 9'b101001001;
assign micromat[64][76] = 9'b100101000;
assign micromat[64][77] = 9'b100100100;
assign micromat[64][78] = 9'b101001001;
assign micromat[64][79] = 9'b110010001;
assign micromat[64][80] = 9'b101110001;
assign micromat[64][81] = 9'b110010110;
assign micromat[64][82] = 9'b110111111;
assign micromat[64][83] = 9'b101001001;
assign micromat[64][84] = 9'b100000000;
assign micromat[64][85] = 9'b100100100;
assign micromat[64][86] = 9'b111111111;
assign micromat[64][87] = 9'b111111111;
assign micromat[64][88] = 9'b111111111;
assign micromat[64][89] = 9'b111111111;
assign micromat[64][90] = 9'b111111111;
assign micromat[64][91] = 9'b111111111;
assign micromat[64][92] = 9'b111111111;
assign micromat[64][93] = 9'b111111111;
assign micromat[64][94] = 9'b111111111;
assign micromat[64][95] = 9'b111111111;
assign micromat[64][96] = 9'b111111111;
assign micromat[64][97] = 9'b111111111;
assign micromat[64][98] = 9'b111111111;
assign micromat[64][99] = 9'b111111111;
assign micromat[65][0] = 9'b111111111;
assign micromat[65][1] = 9'b111111111;
assign micromat[65][2] = 9'b111111111;
assign micromat[65][3] = 9'b111111111;
assign micromat[65][4] = 9'b111111111;
assign micromat[65][5] = 9'b111111111;
assign micromat[65][6] = 9'b111111111;
assign micromat[65][7] = 9'b111111111;
assign micromat[65][8] = 9'b111111111;
assign micromat[65][9] = 9'b111111111;
assign micromat[65][10] = 9'b111111111;
assign micromat[65][11] = 9'b111111111;
assign micromat[65][12] = 9'b111111111;
assign micromat[65][13] = 9'b111111111;
assign micromat[65][14] = 9'b100100100;
assign micromat[65][15] = 9'b100000000;
assign micromat[65][16] = 9'b101101101;
assign micromat[65][17] = 9'b111111111;
assign micromat[65][18] = 9'b111111111;
assign micromat[65][19] = 9'b111111111;
assign micromat[65][20] = 9'b111111111;
assign micromat[65][21] = 9'b111111111;
assign micromat[65][22] = 9'b111111111;
assign micromat[65][23] = 9'b111111111;
assign micromat[65][24] = 9'b111111111;
assign micromat[65][25] = 9'b111111111;
assign micromat[65][26] = 9'b111111111;
assign micromat[65][27] = 9'b111111111;
assign micromat[65][28] = 9'b111111111;
assign micromat[65][29] = 9'b111111111;
assign micromat[65][30] = 9'b111111111;
assign micromat[65][31] = 9'b111111111;
assign micromat[65][32] = 9'b111111111;
assign micromat[65][33] = 9'b111111111;
assign micromat[65][34] = 9'b111111111;
assign micromat[65][35] = 9'b111111111;
assign micromat[65][36] = 9'b111111111;
assign micromat[65][37] = 9'b111111111;
assign micromat[65][38] = 9'b111111111;
assign micromat[65][39] = 9'b111111111;
assign micromat[65][40] = 9'b111111111;
assign micromat[65][41] = 9'b111111111;
assign micromat[65][42] = 9'b111111111;
assign micromat[65][43] = 9'b111111111;
assign micromat[65][44] = 9'b111111111;
assign micromat[65][45] = 9'b111111111;
assign micromat[65][46] = 9'b111111111;
assign micromat[65][47] = 9'b111111111;
assign micromat[65][48] = 9'b111111111;
assign micromat[65][49] = 9'b111111111;
assign micromat[65][50] = 9'b111111111;
assign micromat[65][51] = 9'b111111111;
assign micromat[65][52] = 9'b111111111;
assign micromat[65][53] = 9'b111111111;
assign micromat[65][54] = 9'b111111111;
assign micromat[65][55] = 9'b111111111;
assign micromat[65][56] = 9'b111111111;
assign micromat[65][57] = 9'b111111111;
assign micromat[65][58] = 9'b111111111;
assign micromat[65][59] = 9'b111111111;
assign micromat[65][60] = 9'b111111111;
assign micromat[65][61] = 9'b111111111;
assign micromat[65][62] = 9'b111111111;
assign micromat[65][63] = 9'b111111111;
assign micromat[65][64] = 9'b110110111;
assign micromat[65][65] = 9'b110110111;
assign micromat[65][66] = 9'b101101101;
assign micromat[65][67] = 9'b100000000;
assign micromat[65][68] = 9'b100000000;
assign micromat[65][69] = 9'b111111111;
assign micromat[65][70] = 9'b111111111;
assign micromat[65][71] = 9'b111111111;
assign micromat[65][72] = 9'b111111111;
assign micromat[65][73] = 9'b110111111;
assign micromat[65][74] = 9'b100000000;
assign micromat[65][75] = 9'b100000000;
assign micromat[65][76] = 9'b100000000;
assign micromat[65][77] = 9'b100000000;
assign micromat[65][78] = 9'b100100100;
assign micromat[65][79] = 9'b111111111;
assign micromat[65][80] = 9'b111111111;
assign micromat[65][81] = 9'b110110111;
assign micromat[65][82] = 9'b110111111;
assign micromat[65][83] = 9'b101001001;
assign micromat[65][84] = 9'b100000000;
assign micromat[65][85] = 9'b100100100;
assign micromat[65][86] = 9'b111111111;
assign micromat[65][87] = 9'b111111111;
assign micromat[65][88] = 9'b111111111;
assign micromat[65][89] = 9'b111111111;
assign micromat[65][90] = 9'b111111111;
assign micromat[65][91] = 9'b111111111;
assign micromat[65][92] = 9'b111111111;
assign micromat[65][93] = 9'b111111111;
assign micromat[65][94] = 9'b111111111;
assign micromat[65][95] = 9'b111111111;
assign micromat[65][96] = 9'b111111111;
assign micromat[65][97] = 9'b111111111;
assign micromat[65][98] = 9'b111111111;
assign micromat[65][99] = 9'b111111111;
assign micromat[66][0] = 9'b111111111;
assign micromat[66][1] = 9'b111111111;
assign micromat[66][2] = 9'b111111111;
assign micromat[66][3] = 9'b111111111;
assign micromat[66][4] = 9'b111111111;
assign micromat[66][5] = 9'b111111111;
assign micromat[66][6] = 9'b111111111;
assign micromat[66][7] = 9'b111111111;
assign micromat[66][8] = 9'b111111111;
assign micromat[66][9] = 9'b111111111;
assign micromat[66][10] = 9'b111111111;
assign micromat[66][11] = 9'b111111111;
assign micromat[66][12] = 9'b111111111;
assign micromat[66][13] = 9'b111111111;
assign micromat[66][14] = 9'b100100100;
assign micromat[66][15] = 9'b100000000;
assign micromat[66][16] = 9'b101101101;
assign micromat[66][17] = 9'b111111111;
assign micromat[66][18] = 9'b111111111;
assign micromat[66][19] = 9'b110111111;
assign micromat[66][20] = 9'b110111111;
assign micromat[66][21] = 9'b110111111;
assign micromat[66][22] = 9'b110111111;
assign micromat[66][23] = 9'b110111111;
assign micromat[66][24] = 9'b110111111;
assign micromat[66][25] = 9'b110111111;
assign micromat[66][26] = 9'b110111111;
assign micromat[66][27] = 9'b110111111;
assign micromat[66][28] = 9'b110111111;
assign micromat[66][29] = 9'b110111111;
assign micromat[66][30] = 9'b110111111;
assign micromat[66][31] = 9'b110111111;
assign micromat[66][32] = 9'b110111111;
assign micromat[66][33] = 9'b110111111;
assign micromat[66][34] = 9'b110111111;
assign micromat[66][35] = 9'b110111111;
assign micromat[66][36] = 9'b110111111;
assign micromat[66][37] = 9'b110111111;
assign micromat[66][38] = 9'b110111111;
assign micromat[66][39] = 9'b110111111;
assign micromat[66][40] = 9'b110111111;
assign micromat[66][41] = 9'b110111111;
assign micromat[66][42] = 9'b110111111;
assign micromat[66][43] = 9'b110111111;
assign micromat[66][44] = 9'b110111111;
assign micromat[66][45] = 9'b110111111;
assign micromat[66][46] = 9'b110111111;
assign micromat[66][47] = 9'b110111111;
assign micromat[66][48] = 9'b110111111;
assign micromat[66][49] = 9'b110111111;
assign micromat[66][50] = 9'b110111111;
assign micromat[66][51] = 9'b110111111;
assign micromat[66][52] = 9'b110111111;
assign micromat[66][53] = 9'b110111111;
assign micromat[66][54] = 9'b110111111;
assign micromat[66][55] = 9'b110111111;
assign micromat[66][56] = 9'b110111111;
assign micromat[66][57] = 9'b110111111;
assign micromat[66][58] = 9'b110111111;
assign micromat[66][59] = 9'b110111111;
assign micromat[66][60] = 9'b110111111;
assign micromat[66][61] = 9'b110111111;
assign micromat[66][62] = 9'b110111111;
assign micromat[66][63] = 9'b110111111;
assign micromat[66][64] = 9'b110110111;
assign micromat[66][65] = 9'b110110111;
assign micromat[66][66] = 9'b101101101;
assign micromat[66][67] = 9'b100000000;
assign micromat[66][68] = 9'b100000000;
assign micromat[66][69] = 9'b110111111;
assign micromat[66][70] = 9'b111111111;
assign micromat[66][71] = 9'b111111111;
assign micromat[66][72] = 9'b111111111;
assign micromat[66][73] = 9'b110110111;
assign micromat[66][74] = 9'b100100100;
assign micromat[66][75] = 9'b100100100;
assign micromat[66][76] = 9'b100100100;
assign micromat[66][77] = 9'b100100100;
assign micromat[66][78] = 9'b101001001;
assign micromat[66][79] = 9'b111111111;
assign micromat[66][80] = 9'b110111111;
assign micromat[66][81] = 9'b110110111;
assign micromat[66][82] = 9'b110111111;
assign micromat[66][83] = 9'b101001001;
assign micromat[66][84] = 9'b100000000;
assign micromat[66][85] = 9'b100100100;
assign micromat[66][86] = 9'b111111111;
assign micromat[66][87] = 9'b111111111;
assign micromat[66][88] = 9'b111111111;
assign micromat[66][89] = 9'b111111111;
assign micromat[66][90] = 9'b111111111;
assign micromat[66][91] = 9'b111111111;
assign micromat[66][92] = 9'b111111111;
assign micromat[66][93] = 9'b111111111;
assign micromat[66][94] = 9'b111111111;
assign micromat[66][95] = 9'b111111111;
assign micromat[66][96] = 9'b111111111;
assign micromat[66][97] = 9'b111111111;
assign micromat[66][98] = 9'b111111111;
assign micromat[66][99] = 9'b111111111;
assign micromat[67][0] = 9'b111111111;
assign micromat[67][1] = 9'b111111111;
assign micromat[67][2] = 9'b111111111;
assign micromat[67][3] = 9'b111111111;
assign micromat[67][4] = 9'b111111111;
assign micromat[67][5] = 9'b111111111;
assign micromat[67][6] = 9'b111111111;
assign micromat[67][7] = 9'b111111111;
assign micromat[67][8] = 9'b111111111;
assign micromat[67][9] = 9'b111111111;
assign micromat[67][10] = 9'b111111111;
assign micromat[67][11] = 9'b111111111;
assign micromat[67][12] = 9'b111111111;
assign micromat[67][13] = 9'b111111111;
assign micromat[67][14] = 9'b100100100;
assign micromat[67][15] = 9'b100000000;
assign micromat[67][16] = 9'b101001101;
assign micromat[67][17] = 9'b111111111;
assign micromat[67][18] = 9'b110111111;
assign micromat[67][19] = 9'b110110111;
assign micromat[67][20] = 9'b110110111;
assign micromat[67][21] = 9'b110110111;
assign micromat[67][22] = 9'b110110111;
assign micromat[67][23] = 9'b110110111;
assign micromat[67][24] = 9'b110110111;
assign micromat[67][25] = 9'b110110111;
assign micromat[67][26] = 9'b110110111;
assign micromat[67][27] = 9'b110110111;
assign micromat[67][28] = 9'b110110111;
assign micromat[67][29] = 9'b110110111;
assign micromat[67][30] = 9'b110110111;
assign micromat[67][31] = 9'b110110111;
assign micromat[67][32] = 9'b110110111;
assign micromat[67][33] = 9'b110110111;
assign micromat[67][34] = 9'b110110111;
assign micromat[67][35] = 9'b110110111;
assign micromat[67][36] = 9'b110110111;
assign micromat[67][37] = 9'b110110111;
assign micromat[67][38] = 9'b110110111;
assign micromat[67][39] = 9'b110110111;
assign micromat[67][40] = 9'b110110111;
assign micromat[67][41] = 9'b110110111;
assign micromat[67][42] = 9'b110110111;
assign micromat[67][43] = 9'b110110111;
assign micromat[67][44] = 9'b110110111;
assign micromat[67][45] = 9'b110110111;
assign micromat[67][46] = 9'b110110111;
assign micromat[67][47] = 9'b110110111;
assign micromat[67][48] = 9'b110110111;
assign micromat[67][49] = 9'b110110111;
assign micromat[67][50] = 9'b110110111;
assign micromat[67][51] = 9'b110110111;
assign micromat[67][52] = 9'b110110111;
assign micromat[67][53] = 9'b110110111;
assign micromat[67][54] = 9'b110110111;
assign micromat[67][55] = 9'b110110111;
assign micromat[67][56] = 9'b110110111;
assign micromat[67][57] = 9'b110110111;
assign micromat[67][58] = 9'b110110111;
assign micromat[67][59] = 9'b110110111;
assign micromat[67][60] = 9'b110110111;
assign micromat[67][61] = 9'b110110111;
assign micromat[67][62] = 9'b110110111;
assign micromat[67][63] = 9'b110110111;
assign micromat[67][64] = 9'b110110111;
assign micromat[67][65] = 9'b110111111;
assign micromat[67][66] = 9'b101101101;
assign micromat[67][67] = 9'b100000000;
assign micromat[67][68] = 9'b100000000;
assign micromat[67][69] = 9'b110010110;
assign micromat[67][70] = 9'b111111111;
assign micromat[67][71] = 9'b110111111;
assign micromat[67][72] = 9'b110010110;
assign micromat[67][73] = 9'b110110111;
assign micromat[67][74] = 9'b110111111;
assign micromat[67][75] = 9'b110111111;
assign micromat[67][76] = 9'b110111111;
assign micromat[67][77] = 9'b110111111;
assign micromat[67][78] = 9'b110110111;
assign micromat[67][79] = 9'b110010111;
assign micromat[67][80] = 9'b110110111;
assign micromat[67][81] = 9'b110110111;
assign micromat[67][82] = 9'b110111111;
assign micromat[67][83] = 9'b101001001;
assign micromat[67][84] = 9'b100000000;
assign micromat[67][85] = 9'b100100100;
assign micromat[67][86] = 9'b111111111;
assign micromat[67][87] = 9'b111111111;
assign micromat[67][88] = 9'b111111111;
assign micromat[67][89] = 9'b111111111;
assign micromat[67][90] = 9'b111111111;
assign micromat[67][91] = 9'b111111111;
assign micromat[67][92] = 9'b111111111;
assign micromat[67][93] = 9'b111111111;
assign micromat[67][94] = 9'b111111111;
assign micromat[67][95] = 9'b111111111;
assign micromat[67][96] = 9'b111111111;
assign micromat[67][97] = 9'b111111111;
assign micromat[67][98] = 9'b111111111;
assign micromat[67][99] = 9'b111111111;
assign micromat[68][0] = 9'b111111111;
assign micromat[68][1] = 9'b111111111;
assign micromat[68][2] = 9'b111111111;
assign micromat[68][3] = 9'b111111111;
assign micromat[68][4] = 9'b111111111;
assign micromat[68][5] = 9'b111111111;
assign micromat[68][6] = 9'b111111111;
assign micromat[68][7] = 9'b111111111;
assign micromat[68][8] = 9'b111111111;
assign micromat[68][9] = 9'b111111111;
assign micromat[68][10] = 9'b111111111;
assign micromat[68][11] = 9'b111111111;
assign micromat[68][12] = 9'b111111111;
assign micromat[68][13] = 9'b111111111;
assign micromat[68][14] = 9'b100100100;
assign micromat[68][15] = 9'b100000000;
assign micromat[68][16] = 9'b101001101;
assign micromat[68][17] = 9'b111111111;
assign micromat[68][18] = 9'b111111111;
assign micromat[68][19] = 9'b110110111;
assign micromat[68][20] = 9'b110110111;
assign micromat[68][21] = 9'b110110111;
assign micromat[68][22] = 9'b110110111;
assign micromat[68][23] = 9'b110110111;
assign micromat[68][24] = 9'b110110111;
assign micromat[68][25] = 9'b110110111;
assign micromat[68][26] = 9'b110110111;
assign micromat[68][27] = 9'b110110111;
assign micromat[68][28] = 9'b110110111;
assign micromat[68][29] = 9'b110110111;
assign micromat[68][30] = 9'b110110111;
assign micromat[68][31] = 9'b110110111;
assign micromat[68][32] = 9'b110110111;
assign micromat[68][33] = 9'b110110111;
assign micromat[68][34] = 9'b110110111;
assign micromat[68][35] = 9'b110110111;
assign micromat[68][36] = 9'b110110111;
assign micromat[68][37] = 9'b110110111;
assign micromat[68][38] = 9'b110110111;
assign micromat[68][39] = 9'b110110111;
assign micromat[68][40] = 9'b110110111;
assign micromat[68][41] = 9'b110110111;
assign micromat[68][42] = 9'b110110111;
assign micromat[68][43] = 9'b110110111;
assign micromat[68][44] = 9'b110110111;
assign micromat[68][45] = 9'b110110111;
assign micromat[68][46] = 9'b110110111;
assign micromat[68][47] = 9'b110110111;
assign micromat[68][48] = 9'b110110111;
assign micromat[68][49] = 9'b110110111;
assign micromat[68][50] = 9'b110110111;
assign micromat[68][51] = 9'b110110111;
assign micromat[68][52] = 9'b110110111;
assign micromat[68][53] = 9'b110110111;
assign micromat[68][54] = 9'b110110111;
assign micromat[68][55] = 9'b110110111;
assign micromat[68][56] = 9'b110110111;
assign micromat[68][57] = 9'b110110111;
assign micromat[68][58] = 9'b110110111;
assign micromat[68][59] = 9'b110110111;
assign micromat[68][60] = 9'b110110111;
assign micromat[68][61] = 9'b110110111;
assign micromat[68][62] = 9'b110110111;
assign micromat[68][63] = 9'b110110111;
assign micromat[68][64] = 9'b110110111;
assign micromat[68][65] = 9'b110111111;
assign micromat[68][66] = 9'b101101101;
assign micromat[68][67] = 9'b100000000;
assign micromat[68][68] = 9'b100000000;
assign micromat[68][69] = 9'b110010110;
assign micromat[68][70] = 9'b111111111;
assign micromat[68][71] = 9'b110111111;
assign micromat[68][72] = 9'b110110111;
assign micromat[68][73] = 9'b110110111;
assign micromat[68][74] = 9'b110110111;
assign micromat[68][75] = 9'b110110111;
assign micromat[68][76] = 9'b110110111;
assign micromat[68][77] = 9'b110110111;
assign micromat[68][78] = 9'b110110111;
assign micromat[68][79] = 9'b110110111;
assign micromat[68][80] = 9'b110110111;
assign micromat[68][81] = 9'b110110111;
assign micromat[68][82] = 9'b110111111;
assign micromat[68][83] = 9'b101001001;
assign micromat[68][84] = 9'b100000000;
assign micromat[68][85] = 9'b100100100;
assign micromat[68][86] = 9'b111111111;
assign micromat[68][87] = 9'b111111111;
assign micromat[68][88] = 9'b111111111;
assign micromat[68][89] = 9'b111111111;
assign micromat[68][90] = 9'b111111111;
assign micromat[68][91] = 9'b111111111;
assign micromat[68][92] = 9'b111111111;
assign micromat[68][93] = 9'b111111111;
assign micromat[68][94] = 9'b111111111;
assign micromat[68][95] = 9'b111111111;
assign micromat[68][96] = 9'b111111111;
assign micromat[68][97] = 9'b111111111;
assign micromat[68][98] = 9'b111111111;
assign micromat[68][99] = 9'b111111111;
assign micromat[69][0] = 9'b111111111;
assign micromat[69][1] = 9'b111111111;
assign micromat[69][2] = 9'b111111111;
assign micromat[69][3] = 9'b111111111;
assign micromat[69][4] = 9'b111111111;
assign micromat[69][5] = 9'b111111111;
assign micromat[69][6] = 9'b111111111;
assign micromat[69][7] = 9'b111111111;
assign micromat[69][8] = 9'b111111111;
assign micromat[69][9] = 9'b111111111;
assign micromat[69][10] = 9'b111111111;
assign micromat[69][11] = 9'b111111111;
assign micromat[69][12] = 9'b111111111;
assign micromat[69][13] = 9'b111111111;
assign micromat[69][14] = 9'b111111111;
assign micromat[69][15] = 9'b111111111;
assign micromat[69][16] = 9'b101101101;
assign micromat[69][17] = 9'b100100100;
assign micromat[69][18] = 9'b100100100;
assign micromat[69][19] = 9'b100000000;
assign micromat[69][20] = 9'b100000000;
assign micromat[69][21] = 9'b100000000;
assign micromat[69][22] = 9'b100000000;
assign micromat[69][23] = 9'b100000000;
assign micromat[69][24] = 9'b100000000;
assign micromat[69][25] = 9'b100000000;
assign micromat[69][26] = 9'b100000000;
assign micromat[69][27] = 9'b100000000;
assign micromat[69][28] = 9'b100000000;
assign micromat[69][29] = 9'b100000000;
assign micromat[69][30] = 9'b100000000;
assign micromat[69][31] = 9'b100000000;
assign micromat[69][32] = 9'b100000000;
assign micromat[69][33] = 9'b100000000;
assign micromat[69][34] = 9'b100000000;
assign micromat[69][35] = 9'b100000000;
assign micromat[69][36] = 9'b100000000;
assign micromat[69][37] = 9'b100000000;
assign micromat[69][38] = 9'b100000000;
assign micromat[69][39] = 9'b100000000;
assign micromat[69][40] = 9'b100000000;
assign micromat[69][41] = 9'b100000000;
assign micromat[69][42] = 9'b100000000;
assign micromat[69][43] = 9'b100000000;
assign micromat[69][44] = 9'b100000000;
assign micromat[69][45] = 9'b100000000;
assign micromat[69][46] = 9'b100000000;
assign micromat[69][47] = 9'b100000000;
assign micromat[69][48] = 9'b100000000;
assign micromat[69][49] = 9'b100000000;
assign micromat[69][50] = 9'b100000000;
assign micromat[69][51] = 9'b100000000;
assign micromat[69][52] = 9'b100000000;
assign micromat[69][53] = 9'b100000000;
assign micromat[69][54] = 9'b100000000;
assign micromat[69][55] = 9'b100000000;
assign micromat[69][56] = 9'b100000000;
assign micromat[69][57] = 9'b100000000;
assign micromat[69][58] = 9'b100000000;
assign micromat[69][59] = 9'b100000000;
assign micromat[69][60] = 9'b100000000;
assign micromat[69][61] = 9'b100000000;
assign micromat[69][62] = 9'b100000000;
assign micromat[69][63] = 9'b100000000;
assign micromat[69][64] = 9'b100000000;
assign micromat[69][65] = 9'b100100100;
assign micromat[69][66] = 9'b100000000;
assign micromat[69][67] = 9'b100000000;
assign micromat[69][68] = 9'b100000000;
assign micromat[69][69] = 9'b100000000;
assign micromat[69][70] = 9'b100100100;
assign micromat[69][71] = 9'b100100100;
assign micromat[69][72] = 9'b100000000;
assign micromat[69][73] = 9'b100000000;
assign micromat[69][74] = 9'b100000000;
assign micromat[69][75] = 9'b100000000;
assign micromat[69][76] = 9'b100000000;
assign micromat[69][77] = 9'b100000000;
assign micromat[69][78] = 9'b100000000;
assign micromat[69][79] = 9'b100000000;
assign micromat[69][80] = 9'b100000000;
assign micromat[69][81] = 9'b100000000;
assign micromat[69][82] = 9'b100000000;
assign micromat[69][83] = 9'b101101101;
assign micromat[69][84] = 9'b111111111;
assign micromat[69][85] = 9'b111111111;
assign micromat[69][86] = 9'b111111111;
assign micromat[69][87] = 9'b111111111;
assign micromat[69][88] = 9'b111111111;
assign micromat[69][89] = 9'b111111111;
assign micromat[69][90] = 9'b111111111;
assign micromat[69][91] = 9'b111111111;
assign micromat[69][92] = 9'b111111111;
assign micromat[69][93] = 9'b111111111;
assign micromat[69][94] = 9'b111111111;
assign micromat[69][95] = 9'b111111111;
assign micromat[69][96] = 9'b111111111;
assign micromat[69][97] = 9'b111111111;
assign micromat[69][98] = 9'b111111111;
assign micromat[69][99] = 9'b111111111;
assign micromat[70][0] = 9'b111111111;
assign micromat[70][1] = 9'b111111111;
assign micromat[70][2] = 9'b111111111;
assign micromat[70][3] = 9'b111111111;
assign micromat[70][4] = 9'b111111111;
assign micromat[70][5] = 9'b111111111;
assign micromat[70][6] = 9'b111111111;
assign micromat[70][7] = 9'b111111111;
assign micromat[70][8] = 9'b111111111;
assign micromat[70][9] = 9'b111111111;
assign micromat[70][10] = 9'b111111111;
assign micromat[70][11] = 9'b111111111;
assign micromat[70][12] = 9'b111111111;
assign micromat[70][13] = 9'b111111111;
assign micromat[70][14] = 9'b111111111;
assign micromat[70][15] = 9'b111111111;
assign micromat[70][16] = 9'b101101101;
assign micromat[70][17] = 9'b100000000;
assign micromat[70][18] = 9'b100000000;
assign micromat[70][19] = 9'b100000000;
assign micromat[70][20] = 9'b100000000;
assign micromat[70][21] = 9'b100000000;
assign micromat[70][22] = 9'b100000000;
assign micromat[70][23] = 9'b100000000;
assign micromat[70][24] = 9'b100000000;
assign micromat[70][25] = 9'b100000000;
assign micromat[70][26] = 9'b100000000;
assign micromat[70][27] = 9'b100000000;
assign micromat[70][28] = 9'b100000000;
assign micromat[70][29] = 9'b100000000;
assign micromat[70][30] = 9'b100000000;
assign micromat[70][31] = 9'b100000000;
assign micromat[70][32] = 9'b100000000;
assign micromat[70][33] = 9'b100000000;
assign micromat[70][34] = 9'b100000000;
assign micromat[70][35] = 9'b100000000;
assign micromat[70][36] = 9'b100000000;
assign micromat[70][37] = 9'b100000000;
assign micromat[70][38] = 9'b100000000;
assign micromat[70][39] = 9'b100000000;
assign micromat[70][40] = 9'b100000000;
assign micromat[70][41] = 9'b100000000;
assign micromat[70][42] = 9'b100000000;
assign micromat[70][43] = 9'b100000000;
assign micromat[70][44] = 9'b100000000;
assign micromat[70][45] = 9'b100000000;
assign micromat[70][46] = 9'b100000000;
assign micromat[70][47] = 9'b100000000;
assign micromat[70][48] = 9'b100000000;
assign micromat[70][49] = 9'b100000000;
assign micromat[70][50] = 9'b100000000;
assign micromat[70][51] = 9'b100000000;
assign micromat[70][52] = 9'b100000000;
assign micromat[70][53] = 9'b100000000;
assign micromat[70][54] = 9'b100000000;
assign micromat[70][55] = 9'b100000000;
assign micromat[70][56] = 9'b100000000;
assign micromat[70][57] = 9'b100000000;
assign micromat[70][58] = 9'b100000000;
assign micromat[70][59] = 9'b100000000;
assign micromat[70][60] = 9'b100000000;
assign micromat[70][61] = 9'b100000000;
assign micromat[70][62] = 9'b100000000;
assign micromat[70][63] = 9'b100000000;
assign micromat[70][64] = 9'b100000000;
assign micromat[70][65] = 9'b100000000;
assign micromat[70][66] = 9'b100000000;
assign micromat[70][67] = 9'b100000000;
assign micromat[70][68] = 9'b100000000;
assign micromat[70][69] = 9'b100000000;
assign micromat[70][70] = 9'b100000000;
assign micromat[70][71] = 9'b100000000;
assign micromat[70][72] = 9'b100000000;
assign micromat[70][73] = 9'b100000000;
assign micromat[70][74] = 9'b100000000;
assign micromat[70][75] = 9'b100000000;
assign micromat[70][76] = 9'b100000000;
assign micromat[70][77] = 9'b100000000;
assign micromat[70][78] = 9'b100000000;
assign micromat[70][79] = 9'b100000000;
assign micromat[70][80] = 9'b100000000;
assign micromat[70][81] = 9'b100000000;
assign micromat[70][82] = 9'b100000000;
assign micromat[70][83] = 9'b101101101;
assign micromat[70][84] = 9'b111111111;
assign micromat[70][85] = 9'b111111111;
assign micromat[70][86] = 9'b111111111;
assign micromat[70][87] = 9'b111111111;
assign micromat[70][88] = 9'b111111111;
assign micromat[70][89] = 9'b111111111;
assign micromat[70][90] = 9'b111111111;
assign micromat[70][91] = 9'b111111111;
assign micromat[70][92] = 9'b111111111;
assign micromat[70][93] = 9'b111111111;
assign micromat[70][94] = 9'b111111111;
assign micromat[70][95] = 9'b111111111;
assign micromat[70][96] = 9'b111111111;
assign micromat[70][97] = 9'b111111111;
assign micromat[70][98] = 9'b111111111;
assign micromat[70][99] = 9'b111111111;
assign micromat[71][0] = 9'b111111111;
assign micromat[71][1] = 9'b111111111;
assign micromat[71][2] = 9'b111111111;
assign micromat[71][3] = 9'b111111111;
assign micromat[71][4] = 9'b111111111;
assign micromat[71][5] = 9'b111111111;
assign micromat[71][6] = 9'b111111111;
assign micromat[71][7] = 9'b111111111;
assign micromat[71][8] = 9'b111111111;
assign micromat[71][9] = 9'b111111111;
assign micromat[71][10] = 9'b111111111;
assign micromat[71][11] = 9'b111111111;
assign micromat[71][12] = 9'b111111111;
assign micromat[71][13] = 9'b111111111;
assign micromat[71][14] = 9'b111111111;
assign micromat[71][15] = 9'b111111111;
assign micromat[71][16] = 9'b110110110;
assign micromat[71][17] = 9'b101101101;
assign micromat[71][18] = 9'b101101101;
assign micromat[71][19] = 9'b101101101;
assign micromat[71][20] = 9'b101101101;
assign micromat[71][21] = 9'b101101101;
assign micromat[71][22] = 9'b101101101;
assign micromat[71][23] = 9'b101101101;
assign micromat[71][24] = 9'b101101101;
assign micromat[71][25] = 9'b101101101;
assign micromat[71][26] = 9'b101101101;
assign micromat[71][27] = 9'b101101101;
assign micromat[71][28] = 9'b101101101;
assign micromat[71][29] = 9'b101101101;
assign micromat[71][30] = 9'b101101101;
assign micromat[71][31] = 9'b101101101;
assign micromat[71][32] = 9'b101101101;
assign micromat[71][33] = 9'b101101101;
assign micromat[71][34] = 9'b101101101;
assign micromat[71][35] = 9'b101101101;
assign micromat[71][36] = 9'b101101101;
assign micromat[71][37] = 9'b101101101;
assign micromat[71][38] = 9'b101101101;
assign micromat[71][39] = 9'b101101101;
assign micromat[71][40] = 9'b101101101;
assign micromat[71][41] = 9'b101101101;
assign micromat[71][42] = 9'b101101101;
assign micromat[71][43] = 9'b101101101;
assign micromat[71][44] = 9'b101101101;
assign micromat[71][45] = 9'b101101101;
assign micromat[71][46] = 9'b101101101;
assign micromat[71][47] = 9'b101101101;
assign micromat[71][48] = 9'b101101101;
assign micromat[71][49] = 9'b101101101;
assign micromat[71][50] = 9'b101101101;
assign micromat[71][51] = 9'b101101101;
assign micromat[71][52] = 9'b101101101;
assign micromat[71][53] = 9'b101101101;
assign micromat[71][54] = 9'b101101101;
assign micromat[71][55] = 9'b101101101;
assign micromat[71][56] = 9'b101101101;
assign micromat[71][57] = 9'b101101101;
assign micromat[71][58] = 9'b101101101;
assign micromat[71][59] = 9'b101101101;
assign micromat[71][60] = 9'b101101101;
assign micromat[71][61] = 9'b101101101;
assign micromat[71][62] = 9'b101101101;
assign micromat[71][63] = 9'b101101101;
assign micromat[71][64] = 9'b101101101;
assign micromat[71][65] = 9'b101101101;
assign micromat[71][66] = 9'b101101101;
assign micromat[71][67] = 9'b101101101;
assign micromat[71][68] = 9'b101101101;
assign micromat[71][69] = 9'b101101101;
assign micromat[71][70] = 9'b101101101;
assign micromat[71][71] = 9'b101101101;
assign micromat[71][72] = 9'b101101101;
assign micromat[71][73] = 9'b101101101;
assign micromat[71][74] = 9'b101101101;
assign micromat[71][75] = 9'b101101101;
assign micromat[71][76] = 9'b101101101;
assign micromat[71][77] = 9'b101101101;
assign micromat[71][78] = 9'b101101101;
assign micromat[71][79] = 9'b101101101;
assign micromat[71][80] = 9'b101101101;
assign micromat[71][81] = 9'b101101101;
assign micromat[71][82] = 9'b101101101;
assign micromat[71][83] = 9'b110110110;
assign micromat[71][84] = 9'b111111111;
assign micromat[71][85] = 9'b111111111;
assign micromat[71][86] = 9'b111111111;
assign micromat[71][87] = 9'b111111111;
assign micromat[71][88] = 9'b111111111;
assign micromat[71][89] = 9'b111111111;
assign micromat[71][90] = 9'b111111111;
assign micromat[71][91] = 9'b111111111;
assign micromat[71][92] = 9'b111111111;
assign micromat[71][93] = 9'b111111111;
assign micromat[71][94] = 9'b111111111;
assign micromat[71][95] = 9'b111111111;
assign micromat[71][96] = 9'b111111111;
assign micromat[71][97] = 9'b111111111;
assign micromat[71][98] = 9'b111111111;
assign micromat[71][99] = 9'b111111111;
assign micromat[72][0] = 9'b111111111;
assign micromat[72][1] = 9'b111111111;
assign micromat[72][2] = 9'b111111111;
assign micromat[72][3] = 9'b111111111;
assign micromat[72][4] = 9'b111111111;
assign micromat[72][5] = 9'b111111111;
assign micromat[72][6] = 9'b111111111;
assign micromat[72][7] = 9'b111111111;
assign micromat[72][8] = 9'b111111111;
assign micromat[72][9] = 9'b111111111;
assign micromat[72][10] = 9'b111111111;
assign micromat[72][11] = 9'b111111111;
assign micromat[72][12] = 9'b111111111;
assign micromat[72][13] = 9'b111111111;
assign micromat[72][14] = 9'b111111111;
assign micromat[72][15] = 9'b111111111;
assign micromat[72][16] = 9'b111111111;
assign micromat[72][17] = 9'b111111111;
assign micromat[72][18] = 9'b111111111;
assign micromat[72][19] = 9'b111111111;
assign micromat[72][20] = 9'b111111111;
assign micromat[72][21] = 9'b111111111;
assign micromat[72][22] = 9'b111111111;
assign micromat[72][23] = 9'b111111111;
assign micromat[72][24] = 9'b111111111;
assign micromat[72][25] = 9'b111111111;
assign micromat[72][26] = 9'b111111111;
assign micromat[72][27] = 9'b111111111;
assign micromat[72][28] = 9'b111111111;
assign micromat[72][29] = 9'b111111111;
assign micromat[72][30] = 9'b111111111;
assign micromat[72][31] = 9'b111111111;
assign micromat[72][32] = 9'b111111111;
assign micromat[72][33] = 9'b111111111;
assign micromat[72][34] = 9'b111111111;
assign micromat[72][35] = 9'b111111111;
assign micromat[72][36] = 9'b111111111;
assign micromat[72][37] = 9'b111111111;
assign micromat[72][38] = 9'b111111111;
assign micromat[72][39] = 9'b111111111;
assign micromat[72][40] = 9'b111111111;
assign micromat[72][41] = 9'b111111111;
assign micromat[72][42] = 9'b111111111;
assign micromat[72][43] = 9'b111111111;
assign micromat[72][44] = 9'b111111111;
assign micromat[72][45] = 9'b111111111;
assign micromat[72][46] = 9'b111111111;
assign micromat[72][47] = 9'b111111111;
assign micromat[72][48] = 9'b111111111;
assign micromat[72][49] = 9'b111111111;
assign micromat[72][50] = 9'b111111111;
assign micromat[72][51] = 9'b111111111;
assign micromat[72][52] = 9'b111111111;
assign micromat[72][53] = 9'b111111111;
assign micromat[72][54] = 9'b111111111;
assign micromat[72][55] = 9'b111111111;
assign micromat[72][56] = 9'b111111111;
assign micromat[72][57] = 9'b111111111;
assign micromat[72][58] = 9'b111111111;
assign micromat[72][59] = 9'b111111111;
assign micromat[72][60] = 9'b111111111;
assign micromat[72][61] = 9'b111111111;
assign micromat[72][62] = 9'b111111111;
assign micromat[72][63] = 9'b111111111;
assign micromat[72][64] = 9'b111111111;
assign micromat[72][65] = 9'b111111111;
assign micromat[72][66] = 9'b111111111;
assign micromat[72][67] = 9'b111111111;
assign micromat[72][68] = 9'b111111111;
assign micromat[72][69] = 9'b111111111;
assign micromat[72][70] = 9'b111111111;
assign micromat[72][71] = 9'b111111111;
assign micromat[72][72] = 9'b111111111;
assign micromat[72][73] = 9'b111111111;
assign micromat[72][74] = 9'b111111111;
assign micromat[72][75] = 9'b111111111;
assign micromat[72][76] = 9'b111111111;
assign micromat[72][77] = 9'b111111111;
assign micromat[72][78] = 9'b111111111;
assign micromat[72][79] = 9'b111111111;
assign micromat[72][80] = 9'b111111111;
assign micromat[72][81] = 9'b111111111;
assign micromat[72][82] = 9'b111111111;
assign micromat[72][83] = 9'b111111111;
assign micromat[72][84] = 9'b111111111;
assign micromat[72][85] = 9'b111111111;
assign micromat[72][86] = 9'b111111111;
assign micromat[72][87] = 9'b111111111;
assign micromat[72][88] = 9'b111111111;
assign micromat[72][89] = 9'b111111111;
assign micromat[72][90] = 9'b111111111;
assign micromat[72][91] = 9'b111111111;
assign micromat[72][92] = 9'b111111111;
assign micromat[72][93] = 9'b111111111;
assign micromat[72][94] = 9'b111111111;
assign micromat[72][95] = 9'b111111111;
assign micromat[72][96] = 9'b111111111;
assign micromat[72][97] = 9'b111111111;
assign micromat[72][98] = 9'b111111111;
assign micromat[72][99] = 9'b111111111;
assign micromat[73][0] = 9'b111111111;
assign micromat[73][1] = 9'b111111111;
assign micromat[73][2] = 9'b111111111;
assign micromat[73][3] = 9'b111111111;
assign micromat[73][4] = 9'b111111111;
assign micromat[73][5] = 9'b111111111;
assign micromat[73][6] = 9'b111111111;
assign micromat[73][7] = 9'b111111111;
assign micromat[73][8] = 9'b111111111;
assign micromat[73][9] = 9'b111111111;
assign micromat[73][10] = 9'b111111111;
assign micromat[73][11] = 9'b111111111;
assign micromat[73][12] = 9'b111111111;
assign micromat[73][13] = 9'b111111111;
assign micromat[73][14] = 9'b111111111;
assign micromat[73][15] = 9'b111111111;
assign micromat[73][16] = 9'b111111111;
assign micromat[73][17] = 9'b111111111;
assign micromat[73][18] = 9'b111111111;
assign micromat[73][19] = 9'b111111111;
assign micromat[73][20] = 9'b111111111;
assign micromat[73][21] = 9'b111111111;
assign micromat[73][22] = 9'b111111111;
assign micromat[73][23] = 9'b111111111;
assign micromat[73][24] = 9'b111111111;
assign micromat[73][25] = 9'b111111111;
assign micromat[73][26] = 9'b111111111;
assign micromat[73][27] = 9'b111111111;
assign micromat[73][28] = 9'b111111111;
assign micromat[73][29] = 9'b111111111;
assign micromat[73][30] = 9'b111111111;
assign micromat[73][31] = 9'b111111111;
assign micromat[73][32] = 9'b111111111;
assign micromat[73][33] = 9'b111111111;
assign micromat[73][34] = 9'b111111111;
assign micromat[73][35] = 9'b111111111;
assign micromat[73][36] = 9'b111111111;
assign micromat[73][37] = 9'b111111111;
assign micromat[73][38] = 9'b111111111;
assign micromat[73][39] = 9'b111111111;
assign micromat[73][40] = 9'b111111111;
assign micromat[73][41] = 9'b111111111;
assign micromat[73][42] = 9'b111111111;
assign micromat[73][43] = 9'b111111111;
assign micromat[73][44] = 9'b111111111;
assign micromat[73][45] = 9'b111111111;
assign micromat[73][46] = 9'b111111111;
assign micromat[73][47] = 9'b111111111;
assign micromat[73][48] = 9'b111111111;
assign micromat[73][49] = 9'b111111111;
assign micromat[73][50] = 9'b111111111;
assign micromat[73][51] = 9'b111111111;
assign micromat[73][52] = 9'b111111111;
assign micromat[73][53] = 9'b111111111;
assign micromat[73][54] = 9'b111111111;
assign micromat[73][55] = 9'b111111111;
assign micromat[73][56] = 9'b111111111;
assign micromat[73][57] = 9'b111111111;
assign micromat[73][58] = 9'b111111111;
assign micromat[73][59] = 9'b111111111;
assign micromat[73][60] = 9'b111111111;
assign micromat[73][61] = 9'b111111111;
assign micromat[73][62] = 9'b111111111;
assign micromat[73][63] = 9'b111111111;
assign micromat[73][64] = 9'b111111111;
assign micromat[73][65] = 9'b111111111;
assign micromat[73][66] = 9'b111111111;
assign micromat[73][67] = 9'b111111111;
assign micromat[73][68] = 9'b111111111;
assign micromat[73][69] = 9'b111111111;
assign micromat[73][70] = 9'b111111111;
assign micromat[73][71] = 9'b111111111;
assign micromat[73][72] = 9'b111111111;
assign micromat[73][73] = 9'b111111111;
assign micromat[73][74] = 9'b111111111;
assign micromat[73][75] = 9'b111111111;
assign micromat[73][76] = 9'b111111111;
assign micromat[73][77] = 9'b111111111;
assign micromat[73][78] = 9'b111111111;
assign micromat[73][79] = 9'b111111111;
assign micromat[73][80] = 9'b111111111;
assign micromat[73][81] = 9'b111111111;
assign micromat[73][82] = 9'b111111111;
assign micromat[73][83] = 9'b111111111;
assign micromat[73][84] = 9'b111111111;
assign micromat[73][85] = 9'b111111111;
assign micromat[73][86] = 9'b111111111;
assign micromat[73][87] = 9'b111111111;
assign micromat[73][88] = 9'b111111111;
assign micromat[73][89] = 9'b111111111;
assign micromat[73][90] = 9'b111111111;
assign micromat[73][91] = 9'b111111111;
assign micromat[73][92] = 9'b111111111;
assign micromat[73][93] = 9'b111111111;
assign micromat[73][94] = 9'b111111111;
assign micromat[73][95] = 9'b111111111;
assign micromat[73][96] = 9'b111111111;
assign micromat[73][97] = 9'b111111111;
assign micromat[73][98] = 9'b111111111;
assign micromat[73][99] = 9'b111111111;
assign micromat[74][0] = 9'b111111111;
assign micromat[74][1] = 9'b111111111;
assign micromat[74][2] = 9'b111111111;
assign micromat[74][3] = 9'b111111111;
assign micromat[74][4] = 9'b111111111;
assign micromat[74][5] = 9'b111111111;
assign micromat[74][6] = 9'b111111111;
assign micromat[74][7] = 9'b111111111;
assign micromat[74][8] = 9'b111111111;
assign micromat[74][9] = 9'b111111111;
assign micromat[74][10] = 9'b111111111;
assign micromat[74][11] = 9'b111111111;
assign micromat[74][12] = 9'b111111111;
assign micromat[74][13] = 9'b111111111;
assign micromat[74][14] = 9'b111111111;
assign micromat[74][15] = 9'b111111111;
assign micromat[74][16] = 9'b111111111;
assign micromat[74][17] = 9'b111111111;
assign micromat[74][18] = 9'b111111111;
assign micromat[74][19] = 9'b111111111;
assign micromat[74][20] = 9'b111111111;
assign micromat[74][21] = 9'b111111111;
assign micromat[74][22] = 9'b111111111;
assign micromat[74][23] = 9'b111111111;
assign micromat[74][24] = 9'b111111111;
assign micromat[74][25] = 9'b111111111;
assign micromat[74][26] = 9'b111111111;
assign micromat[74][27] = 9'b111111111;
assign micromat[74][28] = 9'b111111111;
assign micromat[74][29] = 9'b111111111;
assign micromat[74][30] = 9'b111111111;
assign micromat[74][31] = 9'b111111111;
assign micromat[74][32] = 9'b111111111;
assign micromat[74][33] = 9'b111111111;
assign micromat[74][34] = 9'b111111111;
assign micromat[74][35] = 9'b111111111;
assign micromat[74][36] = 9'b111111111;
assign micromat[74][37] = 9'b111111111;
assign micromat[74][38] = 9'b111111111;
assign micromat[74][39] = 9'b111111111;
assign micromat[74][40] = 9'b111111111;
assign micromat[74][41] = 9'b111111111;
assign micromat[74][42] = 9'b111111111;
assign micromat[74][43] = 9'b111111111;
assign micromat[74][44] = 9'b111111111;
assign micromat[74][45] = 9'b111111111;
assign micromat[74][46] = 9'b111111111;
assign micromat[74][47] = 9'b111111111;
assign micromat[74][48] = 9'b111111111;
assign micromat[74][49] = 9'b111111111;
assign micromat[74][50] = 9'b111111111;
assign micromat[74][51] = 9'b111111111;
assign micromat[74][52] = 9'b111111111;
assign micromat[74][53] = 9'b111111111;
assign micromat[74][54] = 9'b111111111;
assign micromat[74][55] = 9'b111111111;
assign micromat[74][56] = 9'b111111111;
assign micromat[74][57] = 9'b111111111;
assign micromat[74][58] = 9'b111111111;
assign micromat[74][59] = 9'b111111111;
assign micromat[74][60] = 9'b111111111;
assign micromat[74][61] = 9'b111111111;
assign micromat[74][62] = 9'b111111111;
assign micromat[74][63] = 9'b111111111;
assign micromat[74][64] = 9'b111111111;
assign micromat[74][65] = 9'b111111111;
assign micromat[74][66] = 9'b111111111;
assign micromat[74][67] = 9'b111111111;
assign micromat[74][68] = 9'b111111111;
assign micromat[74][69] = 9'b111111111;
assign micromat[74][70] = 9'b111111111;
assign micromat[74][71] = 9'b111111111;
assign micromat[74][72] = 9'b111111111;
assign micromat[74][73] = 9'b111111111;
assign micromat[74][74] = 9'b111111111;
assign micromat[74][75] = 9'b111111111;
assign micromat[74][76] = 9'b111111111;
assign micromat[74][77] = 9'b111111111;
assign micromat[74][78] = 9'b111111111;
assign micromat[74][79] = 9'b111111111;
assign micromat[74][80] = 9'b111111111;
assign micromat[74][81] = 9'b111111111;
assign micromat[74][82] = 9'b111111111;
assign micromat[74][83] = 9'b111111111;
assign micromat[74][84] = 9'b111111111;
assign micromat[74][85] = 9'b111111111;
assign micromat[74][86] = 9'b111111111;
assign micromat[74][87] = 9'b111111111;
assign micromat[74][88] = 9'b111111111;
assign micromat[74][89] = 9'b111111111;
assign micromat[74][90] = 9'b111111111;
assign micromat[74][91] = 9'b111111111;
assign micromat[74][92] = 9'b111111111;
assign micromat[74][93] = 9'b111111111;
assign micromat[74][94] = 9'b111111111;
assign micromat[74][95] = 9'b111111111;
assign micromat[74][96] = 9'b111111111;
assign micromat[74][97] = 9'b111111111;
assign micromat[74][98] = 9'b111111111;
assign micromat[74][99] = 9'b111111111;
assign micromat[75][0] = 9'b111111111;
assign micromat[75][1] = 9'b111111111;
assign micromat[75][2] = 9'b111111111;
assign micromat[75][3] = 9'b111111111;
assign micromat[75][4] = 9'b111111111;
assign micromat[75][5] = 9'b111111111;
assign micromat[75][6] = 9'b111111111;
assign micromat[75][7] = 9'b111111111;
assign micromat[75][8] = 9'b111111111;
assign micromat[75][9] = 9'b111111111;
assign micromat[75][10] = 9'b111111111;
assign micromat[75][11] = 9'b111111111;
assign micromat[75][12] = 9'b111111111;
assign micromat[75][13] = 9'b111111111;
assign micromat[75][14] = 9'b111111111;
assign micromat[75][15] = 9'b111111111;
assign micromat[75][16] = 9'b111111111;
assign micromat[75][17] = 9'b111111111;
assign micromat[75][18] = 9'b111111111;
assign micromat[75][19] = 9'b111111111;
assign micromat[75][20] = 9'b111111111;
assign micromat[75][21] = 9'b111111111;
assign micromat[75][22] = 9'b111111111;
assign micromat[75][23] = 9'b111111111;
assign micromat[75][24] = 9'b111111111;
assign micromat[75][25] = 9'b111111111;
assign micromat[75][26] = 9'b111111111;
assign micromat[75][27] = 9'b111111111;
assign micromat[75][28] = 9'b111111111;
assign micromat[75][29] = 9'b111111111;
assign micromat[75][30] = 9'b111111111;
assign micromat[75][31] = 9'b111111111;
assign micromat[75][32] = 9'b111111111;
assign micromat[75][33] = 9'b111111111;
assign micromat[75][34] = 9'b111111111;
assign micromat[75][35] = 9'b111111111;
assign micromat[75][36] = 9'b111111111;
assign micromat[75][37] = 9'b111111111;
assign micromat[75][38] = 9'b111111111;
assign micromat[75][39] = 9'b111111111;
assign micromat[75][40] = 9'b111111111;
assign micromat[75][41] = 9'b111111111;
assign micromat[75][42] = 9'b111111111;
assign micromat[75][43] = 9'b111111111;
assign micromat[75][44] = 9'b111111111;
assign micromat[75][45] = 9'b111111111;
assign micromat[75][46] = 9'b111111111;
assign micromat[75][47] = 9'b111111111;
assign micromat[75][48] = 9'b111111111;
assign micromat[75][49] = 9'b111111111;
assign micromat[75][50] = 9'b111111111;
assign micromat[75][51] = 9'b111111111;
assign micromat[75][52] = 9'b111111111;
assign micromat[75][53] = 9'b111111111;
assign micromat[75][54] = 9'b111111111;
assign micromat[75][55] = 9'b111111111;
assign micromat[75][56] = 9'b111111111;
assign micromat[75][57] = 9'b111111111;
assign micromat[75][58] = 9'b111111111;
assign micromat[75][59] = 9'b111111111;
assign micromat[75][60] = 9'b111111111;
assign micromat[75][61] = 9'b111111111;
assign micromat[75][62] = 9'b111111111;
assign micromat[75][63] = 9'b111111111;
assign micromat[75][64] = 9'b111111111;
assign micromat[75][65] = 9'b111111111;
assign micromat[75][66] = 9'b111111111;
assign micromat[75][67] = 9'b111111111;
assign micromat[75][68] = 9'b111111111;
assign micromat[75][69] = 9'b111111111;
assign micromat[75][70] = 9'b111111111;
assign micromat[75][71] = 9'b111111111;
assign micromat[75][72] = 9'b111111111;
assign micromat[75][73] = 9'b111111111;
assign micromat[75][74] = 9'b111111111;
assign micromat[75][75] = 9'b111111111;
assign micromat[75][76] = 9'b111111111;
assign micromat[75][77] = 9'b111111111;
assign micromat[75][78] = 9'b111111111;
assign micromat[75][79] = 9'b111111111;
assign micromat[75][80] = 9'b111111111;
assign micromat[75][81] = 9'b111111111;
assign micromat[75][82] = 9'b111111111;
assign micromat[75][83] = 9'b111111111;
assign micromat[75][84] = 9'b111111111;
assign micromat[75][85] = 9'b111111111;
assign micromat[75][86] = 9'b111111111;
assign micromat[75][87] = 9'b111111111;
assign micromat[75][88] = 9'b111111111;
assign micromat[75][89] = 9'b111111111;
assign micromat[75][90] = 9'b111111111;
assign micromat[75][91] = 9'b111111111;
assign micromat[75][92] = 9'b111111111;
assign micromat[75][93] = 9'b111111111;
assign micromat[75][94] = 9'b111111111;
assign micromat[75][95] = 9'b111111111;
assign micromat[75][96] = 9'b111111111;
assign micromat[75][97] = 9'b111111111;
assign micromat[75][98] = 9'b111111111;
assign micromat[75][99] = 9'b111111111;
assign micromat[76][0] = 9'b111111111;
assign micromat[76][1] = 9'b111111111;
assign micromat[76][2] = 9'b111111111;
assign micromat[76][3] = 9'b111111111;
assign micromat[76][4] = 9'b111111111;
assign micromat[76][5] = 9'b111111111;
assign micromat[76][6] = 9'b111111111;
assign micromat[76][7] = 9'b111111111;
assign micromat[76][8] = 9'b111111111;
assign micromat[76][9] = 9'b111111111;
assign micromat[76][10] = 9'b111111111;
assign micromat[76][11] = 9'b111111111;
assign micromat[76][12] = 9'b111111111;
assign micromat[76][13] = 9'b111111111;
assign micromat[76][14] = 9'b111111111;
assign micromat[76][15] = 9'b111111111;
assign micromat[76][16] = 9'b111111111;
assign micromat[76][17] = 9'b111111111;
assign micromat[76][18] = 9'b111111111;
assign micromat[76][19] = 9'b111111111;
assign micromat[76][20] = 9'b111111111;
assign micromat[76][21] = 9'b111111111;
assign micromat[76][22] = 9'b111111111;
assign micromat[76][23] = 9'b111111111;
assign micromat[76][24] = 9'b111111111;
assign micromat[76][25] = 9'b111111111;
assign micromat[76][26] = 9'b111111111;
assign micromat[76][27] = 9'b111111111;
assign micromat[76][28] = 9'b111111111;
assign micromat[76][29] = 9'b111111111;
assign micromat[76][30] = 9'b111111111;
assign micromat[76][31] = 9'b111111111;
assign micromat[76][32] = 9'b111111111;
assign micromat[76][33] = 9'b111111111;
assign micromat[76][34] = 9'b111111111;
assign micromat[76][35] = 9'b111111111;
assign micromat[76][36] = 9'b111111111;
assign micromat[76][37] = 9'b111111111;
assign micromat[76][38] = 9'b111111111;
assign micromat[76][39] = 9'b111111111;
assign micromat[76][40] = 9'b111111111;
assign micromat[76][41] = 9'b111111111;
assign micromat[76][42] = 9'b111111111;
assign micromat[76][43] = 9'b111111111;
assign micromat[76][44] = 9'b111111111;
assign micromat[76][45] = 9'b111111111;
assign micromat[76][46] = 9'b111111111;
assign micromat[76][47] = 9'b111111111;
assign micromat[76][48] = 9'b111111111;
assign micromat[76][49] = 9'b111111111;
assign micromat[76][50] = 9'b111111111;
assign micromat[76][51] = 9'b111111111;
assign micromat[76][52] = 9'b111111111;
assign micromat[76][53] = 9'b111111111;
assign micromat[76][54] = 9'b111111111;
assign micromat[76][55] = 9'b111111111;
assign micromat[76][56] = 9'b111111111;
assign micromat[76][57] = 9'b111111111;
assign micromat[76][58] = 9'b111111111;
assign micromat[76][59] = 9'b111111111;
assign micromat[76][60] = 9'b111111111;
assign micromat[76][61] = 9'b111111111;
assign micromat[76][62] = 9'b111111111;
assign micromat[76][63] = 9'b111111111;
assign micromat[76][64] = 9'b111111111;
assign micromat[76][65] = 9'b111111111;
assign micromat[76][66] = 9'b111111111;
assign micromat[76][67] = 9'b111111111;
assign micromat[76][68] = 9'b111111111;
assign micromat[76][69] = 9'b111111111;
assign micromat[76][70] = 9'b111111111;
assign micromat[76][71] = 9'b111111111;
assign micromat[76][72] = 9'b111111111;
assign micromat[76][73] = 9'b111111111;
assign micromat[76][74] = 9'b111111111;
assign micromat[76][75] = 9'b111111111;
assign micromat[76][76] = 9'b111111111;
assign micromat[76][77] = 9'b111111111;
assign micromat[76][78] = 9'b111111111;
assign micromat[76][79] = 9'b111111111;
assign micromat[76][80] = 9'b111111111;
assign micromat[76][81] = 9'b111111111;
assign micromat[76][82] = 9'b111111111;
assign micromat[76][83] = 9'b111111111;
assign micromat[76][84] = 9'b111111111;
assign micromat[76][85] = 9'b111111111;
assign micromat[76][86] = 9'b111111111;
assign micromat[76][87] = 9'b111111111;
assign micromat[76][88] = 9'b111111111;
assign micromat[76][89] = 9'b111111111;
assign micromat[76][90] = 9'b111111111;
assign micromat[76][91] = 9'b111111111;
assign micromat[76][92] = 9'b111111111;
assign micromat[76][93] = 9'b111111111;
assign micromat[76][94] = 9'b111111111;
assign micromat[76][95] = 9'b111111111;
assign micromat[76][96] = 9'b111111111;
assign micromat[76][97] = 9'b111111111;
assign micromat[76][98] = 9'b111111111;
assign micromat[76][99] = 9'b111111111;
assign micromat[77][0] = 9'b111111111;
assign micromat[77][1] = 9'b111111111;
assign micromat[77][2] = 9'b111111111;
assign micromat[77][3] = 9'b111111111;
assign micromat[77][4] = 9'b111111111;
assign micromat[77][5] = 9'b111111111;
assign micromat[77][6] = 9'b111111111;
assign micromat[77][7] = 9'b111111111;
assign micromat[77][8] = 9'b111111111;
assign micromat[77][9] = 9'b111111111;
assign micromat[77][10] = 9'b111111111;
assign micromat[77][11] = 9'b111111111;
assign micromat[77][12] = 9'b111111111;
assign micromat[77][13] = 9'b111111111;
assign micromat[77][14] = 9'b111111111;
assign micromat[77][15] = 9'b111111111;
assign micromat[77][16] = 9'b111111111;
assign micromat[77][17] = 9'b111111111;
assign micromat[77][18] = 9'b111111111;
assign micromat[77][19] = 9'b111111111;
assign micromat[77][20] = 9'b111111111;
assign micromat[77][21] = 9'b111111111;
assign micromat[77][22] = 9'b111111111;
assign micromat[77][23] = 9'b111111111;
assign micromat[77][24] = 9'b111111111;
assign micromat[77][25] = 9'b111111111;
assign micromat[77][26] = 9'b111111111;
assign micromat[77][27] = 9'b111111111;
assign micromat[77][28] = 9'b111111111;
assign micromat[77][29] = 9'b111111111;
assign micromat[77][30] = 9'b111111111;
assign micromat[77][31] = 9'b111111111;
assign micromat[77][32] = 9'b111111111;
assign micromat[77][33] = 9'b111111111;
assign micromat[77][34] = 9'b111111111;
assign micromat[77][35] = 9'b111111111;
assign micromat[77][36] = 9'b111111111;
assign micromat[77][37] = 9'b111111111;
assign micromat[77][38] = 9'b111111111;
assign micromat[77][39] = 9'b111111111;
assign micromat[77][40] = 9'b111111111;
assign micromat[77][41] = 9'b111111111;
assign micromat[77][42] = 9'b111111111;
assign micromat[77][43] = 9'b111111111;
assign micromat[77][44] = 9'b111111111;
assign micromat[77][45] = 9'b111111111;
assign micromat[77][46] = 9'b111111111;
assign micromat[77][47] = 9'b111111111;
assign micromat[77][48] = 9'b111111111;
assign micromat[77][49] = 9'b111111111;
assign micromat[77][50] = 9'b111111111;
assign micromat[77][51] = 9'b111111111;
assign micromat[77][52] = 9'b111111111;
assign micromat[77][53] = 9'b111111111;
assign micromat[77][54] = 9'b111111111;
assign micromat[77][55] = 9'b111111111;
assign micromat[77][56] = 9'b111111111;
assign micromat[77][57] = 9'b111111111;
assign micromat[77][58] = 9'b111111111;
assign micromat[77][59] = 9'b111111111;
assign micromat[77][60] = 9'b111111111;
assign micromat[77][61] = 9'b111111111;
assign micromat[77][62] = 9'b111111111;
assign micromat[77][63] = 9'b111111111;
assign micromat[77][64] = 9'b111111111;
assign micromat[77][65] = 9'b111111111;
assign micromat[77][66] = 9'b111111111;
assign micromat[77][67] = 9'b111111111;
assign micromat[77][68] = 9'b111111111;
assign micromat[77][69] = 9'b111111111;
assign micromat[77][70] = 9'b111111111;
assign micromat[77][71] = 9'b111111111;
assign micromat[77][72] = 9'b111111111;
assign micromat[77][73] = 9'b111111111;
assign micromat[77][74] = 9'b111111111;
assign micromat[77][75] = 9'b111111111;
assign micromat[77][76] = 9'b111111111;
assign micromat[77][77] = 9'b111111111;
assign micromat[77][78] = 9'b111111111;
assign micromat[77][79] = 9'b111111111;
assign micromat[77][80] = 9'b111111111;
assign micromat[77][81] = 9'b111111111;
assign micromat[77][82] = 9'b111111111;
assign micromat[77][83] = 9'b111111111;
assign micromat[77][84] = 9'b111111111;
assign micromat[77][85] = 9'b111111111;
assign micromat[77][86] = 9'b111111111;
assign micromat[77][87] = 9'b111111111;
assign micromat[77][88] = 9'b111111111;
assign micromat[77][89] = 9'b111111111;
assign micromat[77][90] = 9'b111111111;
assign micromat[77][91] = 9'b111111111;
assign micromat[77][92] = 9'b111111111;
assign micromat[77][93] = 9'b111111111;
assign micromat[77][94] = 9'b111111111;
assign micromat[77][95] = 9'b111111111;
assign micromat[77][96] = 9'b111111111;
assign micromat[77][97] = 9'b111111111;
assign micromat[77][98] = 9'b111111111;
assign micromat[77][99] = 9'b111111111;
assign micromat[78][0] = 9'b111111111;
assign micromat[78][1] = 9'b111111111;
assign micromat[78][2] = 9'b111111111;
assign micromat[78][3] = 9'b111111111;
assign micromat[78][4] = 9'b111111111;
assign micromat[78][5] = 9'b111111111;
assign micromat[78][6] = 9'b111111111;
assign micromat[78][7] = 9'b111111111;
assign micromat[78][8] = 9'b111111111;
assign micromat[78][9] = 9'b111111111;
assign micromat[78][10] = 9'b111111111;
assign micromat[78][11] = 9'b111111111;
assign micromat[78][12] = 9'b111111111;
assign micromat[78][13] = 9'b111111111;
assign micromat[78][14] = 9'b111111111;
assign micromat[78][15] = 9'b111111111;
assign micromat[78][16] = 9'b111111111;
assign micromat[78][17] = 9'b111111111;
assign micromat[78][18] = 9'b111111111;
assign micromat[78][19] = 9'b111111111;
assign micromat[78][20] = 9'b111111111;
assign micromat[78][21] = 9'b111111111;
assign micromat[78][22] = 9'b111111111;
assign micromat[78][23] = 9'b111111111;
assign micromat[78][24] = 9'b111111111;
assign micromat[78][25] = 9'b111111111;
assign micromat[78][26] = 9'b111111111;
assign micromat[78][27] = 9'b111111111;
assign micromat[78][28] = 9'b111111111;
assign micromat[78][29] = 9'b111111111;
assign micromat[78][30] = 9'b111111111;
assign micromat[78][31] = 9'b111111111;
assign micromat[78][32] = 9'b111111111;
assign micromat[78][33] = 9'b111111111;
assign micromat[78][34] = 9'b111111111;
assign micromat[78][35] = 9'b111111111;
assign micromat[78][36] = 9'b111111111;
assign micromat[78][37] = 9'b111111111;
assign micromat[78][38] = 9'b111111111;
assign micromat[78][39] = 9'b111111111;
assign micromat[78][40] = 9'b111111111;
assign micromat[78][41] = 9'b111111111;
assign micromat[78][42] = 9'b111111111;
assign micromat[78][43] = 9'b111111111;
assign micromat[78][44] = 9'b111111111;
assign micromat[78][45] = 9'b111111111;
assign micromat[78][46] = 9'b111111111;
assign micromat[78][47] = 9'b111111111;
assign micromat[78][48] = 9'b111111111;
assign micromat[78][49] = 9'b111111111;
assign micromat[78][50] = 9'b111111111;
assign micromat[78][51] = 9'b111111111;
assign micromat[78][52] = 9'b111111111;
assign micromat[78][53] = 9'b111111111;
assign micromat[78][54] = 9'b111111111;
assign micromat[78][55] = 9'b111111111;
assign micromat[78][56] = 9'b111111111;
assign micromat[78][57] = 9'b111111111;
assign micromat[78][58] = 9'b111111111;
assign micromat[78][59] = 9'b111111111;
assign micromat[78][60] = 9'b111111111;
assign micromat[78][61] = 9'b111111111;
assign micromat[78][62] = 9'b111111111;
assign micromat[78][63] = 9'b111111111;
assign micromat[78][64] = 9'b111111111;
assign micromat[78][65] = 9'b111111111;
assign micromat[78][66] = 9'b111111111;
assign micromat[78][67] = 9'b111111111;
assign micromat[78][68] = 9'b111111111;
assign micromat[78][69] = 9'b111111111;
assign micromat[78][70] = 9'b111111111;
assign micromat[78][71] = 9'b111111111;
assign micromat[78][72] = 9'b111111111;
assign micromat[78][73] = 9'b111111111;
assign micromat[78][74] = 9'b111111111;
assign micromat[78][75] = 9'b111111111;
assign micromat[78][76] = 9'b111111111;
assign micromat[78][77] = 9'b111111111;
assign micromat[78][78] = 9'b111111111;
assign micromat[78][79] = 9'b111111111;
assign micromat[78][80] = 9'b111111111;
assign micromat[78][81] = 9'b111111111;
assign micromat[78][82] = 9'b111111111;
assign micromat[78][83] = 9'b111111111;
assign micromat[78][84] = 9'b111111111;
assign micromat[78][85] = 9'b111111111;
assign micromat[78][86] = 9'b111111111;
assign micromat[78][87] = 9'b111111111;
assign micromat[78][88] = 9'b111111111;
assign micromat[78][89] = 9'b111111111;
assign micromat[78][90] = 9'b111111111;
assign micromat[78][91] = 9'b111111111;
assign micromat[78][92] = 9'b111111111;
assign micromat[78][93] = 9'b111111111;
assign micromat[78][94] = 9'b111111111;
assign micromat[78][95] = 9'b111111111;
assign micromat[78][96] = 9'b111111111;
assign micromat[78][97] = 9'b111111111;
assign micromat[78][98] = 9'b111111111;
assign micromat[78][99] = 9'b111111111;
assign micromat[79][0] = 9'b111111111;
assign micromat[79][1] = 9'b111111111;
assign micromat[79][2] = 9'b111111111;
assign micromat[79][3] = 9'b111111111;
assign micromat[79][4] = 9'b111111111;
assign micromat[79][5] = 9'b111111111;
assign micromat[79][6] = 9'b111111111;
assign micromat[79][7] = 9'b111111111;
assign micromat[79][8] = 9'b111111111;
assign micromat[79][9] = 9'b111111111;
assign micromat[79][10] = 9'b111111111;
assign micromat[79][11] = 9'b111111111;
assign micromat[79][12] = 9'b111111111;
assign micromat[79][13] = 9'b111111111;
assign micromat[79][14] = 9'b111111111;
assign micromat[79][15] = 9'b111111111;
assign micromat[79][16] = 9'b111111111;
assign micromat[79][17] = 9'b111111111;
assign micromat[79][18] = 9'b111111111;
assign micromat[79][19] = 9'b111111111;
assign micromat[79][20] = 9'b111111111;
assign micromat[79][21] = 9'b111111111;
assign micromat[79][22] = 9'b111111111;
assign micromat[79][23] = 9'b111111111;
assign micromat[79][24] = 9'b111111111;
assign micromat[79][25] = 9'b111111111;
assign micromat[79][26] = 9'b111111111;
assign micromat[79][27] = 9'b111111111;
assign micromat[79][28] = 9'b111111111;
assign micromat[79][29] = 9'b111111111;
assign micromat[79][30] = 9'b111111111;
assign micromat[79][31] = 9'b111111111;
assign micromat[79][32] = 9'b111111111;
assign micromat[79][33] = 9'b111111111;
assign micromat[79][34] = 9'b111111111;
assign micromat[79][35] = 9'b111111111;
assign micromat[79][36] = 9'b111111111;
assign micromat[79][37] = 9'b111111111;
assign micromat[79][38] = 9'b111111111;
assign micromat[79][39] = 9'b111111111;
assign micromat[79][40] = 9'b111111111;
assign micromat[79][41] = 9'b111111111;
assign micromat[79][42] = 9'b111111111;
assign micromat[79][43] = 9'b111111111;
assign micromat[79][44] = 9'b111111111;
assign micromat[79][45] = 9'b111111111;
assign micromat[79][46] = 9'b111111111;
assign micromat[79][47] = 9'b111111111;
assign micromat[79][48] = 9'b111111111;
assign micromat[79][49] = 9'b111111111;
assign micromat[79][50] = 9'b111111111;
assign micromat[79][51] = 9'b111111111;
assign micromat[79][52] = 9'b111111111;
assign micromat[79][53] = 9'b111111111;
assign micromat[79][54] = 9'b111111111;
assign micromat[79][55] = 9'b111111111;
assign micromat[79][56] = 9'b111111111;
assign micromat[79][57] = 9'b111111111;
assign micromat[79][58] = 9'b111111111;
assign micromat[79][59] = 9'b111111111;
assign micromat[79][60] = 9'b111111111;
assign micromat[79][61] = 9'b111111111;
assign micromat[79][62] = 9'b111111111;
assign micromat[79][63] = 9'b111111111;
assign micromat[79][64] = 9'b111111111;
assign micromat[79][65] = 9'b111111111;
assign micromat[79][66] = 9'b111111111;
assign micromat[79][67] = 9'b111111111;
assign micromat[79][68] = 9'b111111111;
assign micromat[79][69] = 9'b111111111;
assign micromat[79][70] = 9'b111111111;
assign micromat[79][71] = 9'b111111111;
assign micromat[79][72] = 9'b111111111;
assign micromat[79][73] = 9'b111111111;
assign micromat[79][74] = 9'b111111111;
assign micromat[79][75] = 9'b111111111;
assign micromat[79][76] = 9'b111111111;
assign micromat[79][77] = 9'b111111111;
assign micromat[79][78] = 9'b111111111;
assign micromat[79][79] = 9'b111111111;
assign micromat[79][80] = 9'b111111111;
assign micromat[79][81] = 9'b111111111;
assign micromat[79][82] = 9'b111111111;
assign micromat[79][83] = 9'b111111111;
assign micromat[79][84] = 9'b111111111;
assign micromat[79][85] = 9'b111111111;
assign micromat[79][86] = 9'b111111111;
assign micromat[79][87] = 9'b111111111;
assign micromat[79][88] = 9'b111111111;
assign micromat[79][89] = 9'b111111111;
assign micromat[79][90] = 9'b111111111;
assign micromat[79][91] = 9'b111111111;
assign micromat[79][92] = 9'b111111111;
assign micromat[79][93] = 9'b111111111;
assign micromat[79][94] = 9'b111111111;
assign micromat[79][95] = 9'b111111111;
assign micromat[79][96] = 9'b111111111;
assign micromat[79][97] = 9'b111111111;
assign micromat[79][98] = 9'b111111111;
assign micromat[79][99] = 9'b111111111;
assign micromat[80][0] = 9'b111111111;
assign micromat[80][1] = 9'b111111111;
assign micromat[80][2] = 9'b111111111;
assign micromat[80][3] = 9'b111111111;
assign micromat[80][4] = 9'b111111111;
assign micromat[80][5] = 9'b111111111;
assign micromat[80][6] = 9'b111111111;
assign micromat[80][7] = 9'b111111111;
assign micromat[80][8] = 9'b111111111;
assign micromat[80][9] = 9'b111111111;
assign micromat[80][10] = 9'b111111111;
assign micromat[80][11] = 9'b111111111;
assign micromat[80][12] = 9'b111111111;
assign micromat[80][13] = 9'b111111111;
assign micromat[80][14] = 9'b111111111;
assign micromat[80][15] = 9'b111111111;
assign micromat[80][16] = 9'b111111111;
assign micromat[80][17] = 9'b111111111;
assign micromat[80][18] = 9'b111111111;
assign micromat[80][19] = 9'b111111111;
assign micromat[80][20] = 9'b111111111;
assign micromat[80][21] = 9'b111111111;
assign micromat[80][22] = 9'b111111111;
assign micromat[80][23] = 9'b111111111;
assign micromat[80][24] = 9'b111111111;
assign micromat[80][25] = 9'b111111111;
assign micromat[80][26] = 9'b111111111;
assign micromat[80][27] = 9'b111111111;
assign micromat[80][28] = 9'b111111111;
assign micromat[80][29] = 9'b111111111;
assign micromat[80][30] = 9'b111111111;
assign micromat[80][31] = 9'b111111111;
assign micromat[80][32] = 9'b111111111;
assign micromat[80][33] = 9'b111111111;
assign micromat[80][34] = 9'b111111111;
assign micromat[80][35] = 9'b111111111;
assign micromat[80][36] = 9'b111111111;
assign micromat[80][37] = 9'b111111111;
assign micromat[80][38] = 9'b111111111;
assign micromat[80][39] = 9'b111111111;
assign micromat[80][40] = 9'b111111111;
assign micromat[80][41] = 9'b111111111;
assign micromat[80][42] = 9'b111111111;
assign micromat[80][43] = 9'b111111111;
assign micromat[80][44] = 9'b111111111;
assign micromat[80][45] = 9'b111111111;
assign micromat[80][46] = 9'b111111111;
assign micromat[80][47] = 9'b111111111;
assign micromat[80][48] = 9'b111111111;
assign micromat[80][49] = 9'b111111111;
assign micromat[80][50] = 9'b111111111;
assign micromat[80][51] = 9'b111111111;
assign micromat[80][52] = 9'b111111111;
assign micromat[80][53] = 9'b111111111;
assign micromat[80][54] = 9'b111111111;
assign micromat[80][55] = 9'b111111111;
assign micromat[80][56] = 9'b111111111;
assign micromat[80][57] = 9'b111111111;
assign micromat[80][58] = 9'b111111111;
assign micromat[80][59] = 9'b111111111;
assign micromat[80][60] = 9'b111111111;
assign micromat[80][61] = 9'b111111111;
assign micromat[80][62] = 9'b111111111;
assign micromat[80][63] = 9'b111111111;
assign micromat[80][64] = 9'b111111111;
assign micromat[80][65] = 9'b111111111;
assign micromat[80][66] = 9'b111111111;
assign micromat[80][67] = 9'b111111111;
assign micromat[80][68] = 9'b111111111;
assign micromat[80][69] = 9'b111111111;
assign micromat[80][70] = 9'b111111111;
assign micromat[80][71] = 9'b111111111;
assign micromat[80][72] = 9'b111111111;
assign micromat[80][73] = 9'b111111111;
assign micromat[80][74] = 9'b111111111;
assign micromat[80][75] = 9'b111111111;
assign micromat[80][76] = 9'b111111111;
assign micromat[80][77] = 9'b111111111;
assign micromat[80][78] = 9'b111111111;
assign micromat[80][79] = 9'b111111111;
assign micromat[80][80] = 9'b111111111;
assign micromat[80][81] = 9'b111111111;
assign micromat[80][82] = 9'b111111111;
assign micromat[80][83] = 9'b111111111;
assign micromat[80][84] = 9'b111111111;
assign micromat[80][85] = 9'b111111111;
assign micromat[80][86] = 9'b111111111;
assign micromat[80][87] = 9'b111111111;
assign micromat[80][88] = 9'b111111111;
assign micromat[80][89] = 9'b111111111;
assign micromat[80][90] = 9'b111111111;
assign micromat[80][91] = 9'b111111111;
assign micromat[80][92] = 9'b111111111;
assign micromat[80][93] = 9'b111111111;
assign micromat[80][94] = 9'b111111111;
assign micromat[80][95] = 9'b111111111;
assign micromat[80][96] = 9'b111111111;
assign micromat[80][97] = 9'b111111111;
assign micromat[80][98] = 9'b111111111;
assign micromat[80][99] = 9'b111111111;
assign micromat[81][0] = 9'b111111111;
assign micromat[81][1] = 9'b111111111;
assign micromat[81][2] = 9'b111111111;
assign micromat[81][3] = 9'b111111111;
assign micromat[81][4] = 9'b111111111;
assign micromat[81][5] = 9'b111111111;
assign micromat[81][6] = 9'b111111111;
assign micromat[81][7] = 9'b111111111;
assign micromat[81][8] = 9'b111111111;
assign micromat[81][9] = 9'b111111111;
assign micromat[81][10] = 9'b111111111;
assign micromat[81][11] = 9'b111111111;
assign micromat[81][12] = 9'b111111111;
assign micromat[81][13] = 9'b111111111;
assign micromat[81][14] = 9'b111111111;
assign micromat[81][15] = 9'b111111111;
assign micromat[81][16] = 9'b111111111;
assign micromat[81][17] = 9'b111111111;
assign micromat[81][18] = 9'b111111111;
assign micromat[81][19] = 9'b111111111;
assign micromat[81][20] = 9'b111111111;
assign micromat[81][21] = 9'b111111111;
assign micromat[81][22] = 9'b111111111;
assign micromat[81][23] = 9'b111111111;
assign micromat[81][24] = 9'b111111111;
assign micromat[81][25] = 9'b111111111;
assign micromat[81][26] = 9'b111111111;
assign micromat[81][27] = 9'b111111111;
assign micromat[81][28] = 9'b111111111;
assign micromat[81][29] = 9'b111111111;
assign micromat[81][30] = 9'b111111111;
assign micromat[81][31] = 9'b111111111;
assign micromat[81][32] = 9'b111111111;
assign micromat[81][33] = 9'b111111111;
assign micromat[81][34] = 9'b111111111;
assign micromat[81][35] = 9'b111111111;
assign micromat[81][36] = 9'b111111111;
assign micromat[81][37] = 9'b111111111;
assign micromat[81][38] = 9'b111111111;
assign micromat[81][39] = 9'b111111111;
assign micromat[81][40] = 9'b111111111;
assign micromat[81][41] = 9'b111111111;
assign micromat[81][42] = 9'b111111111;
assign micromat[81][43] = 9'b111111111;
assign micromat[81][44] = 9'b111111111;
assign micromat[81][45] = 9'b111111111;
assign micromat[81][46] = 9'b111111111;
assign micromat[81][47] = 9'b111111111;
assign micromat[81][48] = 9'b111111111;
assign micromat[81][49] = 9'b111111111;
assign micromat[81][50] = 9'b111111111;
assign micromat[81][51] = 9'b111111111;
assign micromat[81][52] = 9'b111111111;
assign micromat[81][53] = 9'b111111111;
assign micromat[81][54] = 9'b111111111;
assign micromat[81][55] = 9'b111111111;
assign micromat[81][56] = 9'b111111111;
assign micromat[81][57] = 9'b111111111;
assign micromat[81][58] = 9'b111111111;
assign micromat[81][59] = 9'b111111111;
assign micromat[81][60] = 9'b111111111;
assign micromat[81][61] = 9'b111111111;
assign micromat[81][62] = 9'b111111111;
assign micromat[81][63] = 9'b111111111;
assign micromat[81][64] = 9'b111111111;
assign micromat[81][65] = 9'b111111111;
assign micromat[81][66] = 9'b111111111;
assign micromat[81][67] = 9'b111111111;
assign micromat[81][68] = 9'b111111111;
assign micromat[81][69] = 9'b111111111;
assign micromat[81][70] = 9'b111111111;
assign micromat[81][71] = 9'b111111111;
assign micromat[81][72] = 9'b111111111;
assign micromat[81][73] = 9'b111111111;
assign micromat[81][74] = 9'b111111111;
assign micromat[81][75] = 9'b111111111;
assign micromat[81][76] = 9'b111111111;
assign micromat[81][77] = 9'b111111111;
assign micromat[81][78] = 9'b111111111;
assign micromat[81][79] = 9'b111111111;
assign micromat[81][80] = 9'b111111111;
assign micromat[81][81] = 9'b111111111;
assign micromat[81][82] = 9'b111111111;
assign micromat[81][83] = 9'b111111111;
assign micromat[81][84] = 9'b111111111;
assign micromat[81][85] = 9'b111111111;
assign micromat[81][86] = 9'b111111111;
assign micromat[81][87] = 9'b111111111;
assign micromat[81][88] = 9'b111111111;
assign micromat[81][89] = 9'b111111111;
assign micromat[81][90] = 9'b111111111;
assign micromat[81][91] = 9'b111111111;
assign micromat[81][92] = 9'b111111111;
assign micromat[81][93] = 9'b111111111;
assign micromat[81][94] = 9'b111111111;
assign micromat[81][95] = 9'b111111111;
assign micromat[81][96] = 9'b111111111;
assign micromat[81][97] = 9'b111111111;
assign micromat[81][98] = 9'b111111111;
assign micromat[81][99] = 9'b111111111;
assign micromat[82][0] = 9'b111111111;
assign micromat[82][1] = 9'b111111111;
assign micromat[82][2] = 9'b111111111;
assign micromat[82][3] = 9'b111111111;
assign micromat[82][4] = 9'b111111111;
assign micromat[82][5] = 9'b111111111;
assign micromat[82][6] = 9'b111111111;
assign micromat[82][7] = 9'b111111111;
assign micromat[82][8] = 9'b111111111;
assign micromat[82][9] = 9'b111111111;
assign micromat[82][10] = 9'b111111111;
assign micromat[82][11] = 9'b111111111;
assign micromat[82][12] = 9'b111111111;
assign micromat[82][13] = 9'b111111111;
assign micromat[82][14] = 9'b111111111;
assign micromat[82][15] = 9'b111111111;
assign micromat[82][16] = 9'b111111111;
assign micromat[82][17] = 9'b111111111;
assign micromat[82][18] = 9'b111111111;
assign micromat[82][19] = 9'b111111111;
assign micromat[82][20] = 9'b111111111;
assign micromat[82][21] = 9'b111111111;
assign micromat[82][22] = 9'b111111111;
assign micromat[82][23] = 9'b111111111;
assign micromat[82][24] = 9'b111111111;
assign micromat[82][25] = 9'b111111111;
assign micromat[82][26] = 9'b111111111;
assign micromat[82][27] = 9'b111111111;
assign micromat[82][28] = 9'b111111111;
assign micromat[82][29] = 9'b111111111;
assign micromat[82][30] = 9'b111111111;
assign micromat[82][31] = 9'b111111111;
assign micromat[82][32] = 9'b111111111;
assign micromat[82][33] = 9'b111111111;
assign micromat[82][34] = 9'b111111111;
assign micromat[82][35] = 9'b111111111;
assign micromat[82][36] = 9'b111111111;
assign micromat[82][37] = 9'b111111111;
assign micromat[82][38] = 9'b111111111;
assign micromat[82][39] = 9'b111111111;
assign micromat[82][40] = 9'b111111111;
assign micromat[82][41] = 9'b111111111;
assign micromat[82][42] = 9'b111111111;
assign micromat[82][43] = 9'b111111111;
assign micromat[82][44] = 9'b111111111;
assign micromat[82][45] = 9'b111111111;
assign micromat[82][46] = 9'b111111111;
assign micromat[82][47] = 9'b111111111;
assign micromat[82][48] = 9'b111111111;
assign micromat[82][49] = 9'b111111111;
assign micromat[82][50] = 9'b111111111;
assign micromat[82][51] = 9'b111111111;
assign micromat[82][52] = 9'b111111111;
assign micromat[82][53] = 9'b111111111;
assign micromat[82][54] = 9'b111111111;
assign micromat[82][55] = 9'b111111111;
assign micromat[82][56] = 9'b111111111;
assign micromat[82][57] = 9'b111111111;
assign micromat[82][58] = 9'b111111111;
assign micromat[82][59] = 9'b111111111;
assign micromat[82][60] = 9'b111111111;
assign micromat[82][61] = 9'b111111111;
assign micromat[82][62] = 9'b111111111;
assign micromat[82][63] = 9'b111111111;
assign micromat[82][64] = 9'b111111111;
assign micromat[82][65] = 9'b111111111;
assign micromat[82][66] = 9'b111111111;
assign micromat[82][67] = 9'b111111111;
assign micromat[82][68] = 9'b111111111;
assign micromat[82][69] = 9'b111111111;
assign micromat[82][70] = 9'b111111111;
assign micromat[82][71] = 9'b111111111;
assign micromat[82][72] = 9'b111111111;
assign micromat[82][73] = 9'b111111111;
assign micromat[82][74] = 9'b111111111;
assign micromat[82][75] = 9'b111111111;
assign micromat[82][76] = 9'b111111111;
assign micromat[82][77] = 9'b111111111;
assign micromat[82][78] = 9'b111111111;
assign micromat[82][79] = 9'b111111111;
assign micromat[82][80] = 9'b111111111;
assign micromat[82][81] = 9'b111111111;
assign micromat[82][82] = 9'b111111111;
assign micromat[82][83] = 9'b111111111;
assign micromat[82][84] = 9'b111111111;
assign micromat[82][85] = 9'b111111111;
assign micromat[82][86] = 9'b111111111;
assign micromat[82][87] = 9'b111111111;
assign micromat[82][88] = 9'b111111111;
assign micromat[82][89] = 9'b111111111;
assign micromat[82][90] = 9'b111111111;
assign micromat[82][91] = 9'b111111111;
assign micromat[82][92] = 9'b111111111;
assign micromat[82][93] = 9'b111111111;
assign micromat[82][94] = 9'b111111111;
assign micromat[82][95] = 9'b111111111;
assign micromat[82][96] = 9'b111111111;
assign micromat[82][97] = 9'b111111111;
assign micromat[82][98] = 9'b111111111;
assign micromat[82][99] = 9'b111111111;
assign micromat[83][0] = 9'b111111111;
assign micromat[83][1] = 9'b111111111;
assign micromat[83][2] = 9'b111111111;
assign micromat[83][3] = 9'b111111111;
assign micromat[83][4] = 9'b111111111;
assign micromat[83][5] = 9'b111111111;
assign micromat[83][6] = 9'b111111111;
assign micromat[83][7] = 9'b111111111;
assign micromat[83][8] = 9'b111111111;
assign micromat[83][9] = 9'b111111111;
assign micromat[83][10] = 9'b111111111;
assign micromat[83][11] = 9'b111111111;
assign micromat[83][12] = 9'b111111111;
assign micromat[83][13] = 9'b111111111;
assign micromat[83][14] = 9'b111111111;
assign micromat[83][15] = 9'b111111111;
assign micromat[83][16] = 9'b111111111;
assign micromat[83][17] = 9'b111111111;
assign micromat[83][18] = 9'b111111111;
assign micromat[83][19] = 9'b111111111;
assign micromat[83][20] = 9'b111111111;
assign micromat[83][21] = 9'b111111111;
assign micromat[83][22] = 9'b111111111;
assign micromat[83][23] = 9'b111111111;
assign micromat[83][24] = 9'b111111111;
assign micromat[83][25] = 9'b111111111;
assign micromat[83][26] = 9'b111111111;
assign micromat[83][27] = 9'b111111111;
assign micromat[83][28] = 9'b111111111;
assign micromat[83][29] = 9'b111111111;
assign micromat[83][30] = 9'b111111111;
assign micromat[83][31] = 9'b111111111;
assign micromat[83][32] = 9'b111111111;
assign micromat[83][33] = 9'b111111111;
assign micromat[83][34] = 9'b111111111;
assign micromat[83][35] = 9'b111111111;
assign micromat[83][36] = 9'b111111111;
assign micromat[83][37] = 9'b111111111;
assign micromat[83][38] = 9'b111111111;
assign micromat[83][39] = 9'b111111111;
assign micromat[83][40] = 9'b111111111;
assign micromat[83][41] = 9'b111111111;
assign micromat[83][42] = 9'b111111111;
assign micromat[83][43] = 9'b111111111;
assign micromat[83][44] = 9'b111111111;
assign micromat[83][45] = 9'b111111111;
assign micromat[83][46] = 9'b111111111;
assign micromat[83][47] = 9'b111111111;
assign micromat[83][48] = 9'b111111111;
assign micromat[83][49] = 9'b111111111;
assign micromat[83][50] = 9'b111111111;
assign micromat[83][51] = 9'b111111111;
assign micromat[83][52] = 9'b111111111;
assign micromat[83][53] = 9'b111111111;
assign micromat[83][54] = 9'b111111111;
assign micromat[83][55] = 9'b111111111;
assign micromat[83][56] = 9'b111111111;
assign micromat[83][57] = 9'b111111111;
assign micromat[83][58] = 9'b111111111;
assign micromat[83][59] = 9'b111111111;
assign micromat[83][60] = 9'b111111111;
assign micromat[83][61] = 9'b111111111;
assign micromat[83][62] = 9'b111111111;
assign micromat[83][63] = 9'b111111111;
assign micromat[83][64] = 9'b111111111;
assign micromat[83][65] = 9'b111111111;
assign micromat[83][66] = 9'b111111111;
assign micromat[83][67] = 9'b111111111;
assign micromat[83][68] = 9'b111111111;
assign micromat[83][69] = 9'b111111111;
assign micromat[83][70] = 9'b111111111;
assign micromat[83][71] = 9'b111111111;
assign micromat[83][72] = 9'b111111111;
assign micromat[83][73] = 9'b111111111;
assign micromat[83][74] = 9'b111111111;
assign micromat[83][75] = 9'b111111111;
assign micromat[83][76] = 9'b111111111;
assign micromat[83][77] = 9'b111111111;
assign micromat[83][78] = 9'b111111111;
assign micromat[83][79] = 9'b111111111;
assign micromat[83][80] = 9'b111111111;
assign micromat[83][81] = 9'b111111111;
assign micromat[83][82] = 9'b111111111;
assign micromat[83][83] = 9'b111111111;
assign micromat[83][84] = 9'b111111111;
assign micromat[83][85] = 9'b111111111;
assign micromat[83][86] = 9'b111111111;
assign micromat[83][87] = 9'b111111111;
assign micromat[83][88] = 9'b111111111;
assign micromat[83][89] = 9'b111111111;
assign micromat[83][90] = 9'b111111111;
assign micromat[83][91] = 9'b111111111;
assign micromat[83][92] = 9'b111111111;
assign micromat[83][93] = 9'b111111111;
assign micromat[83][94] = 9'b111111111;
assign micromat[83][95] = 9'b111111111;
assign micromat[83][96] = 9'b111111111;
assign micromat[83][97] = 9'b111111111;
assign micromat[83][98] = 9'b111111111;
assign micromat[83][99] = 9'b111111111;
assign micromat[84][0] = 9'b111111111;
assign micromat[84][1] = 9'b111111111;
assign micromat[84][2] = 9'b111111111;
assign micromat[84][3] = 9'b111111111;
assign micromat[84][4] = 9'b111111111;
assign micromat[84][5] = 9'b111111111;
assign micromat[84][6] = 9'b111111111;
assign micromat[84][7] = 9'b111111111;
assign micromat[84][8] = 9'b111111111;
assign micromat[84][9] = 9'b111111111;
assign micromat[84][10] = 9'b111111111;
assign micromat[84][11] = 9'b111111111;
assign micromat[84][12] = 9'b111111111;
assign micromat[84][13] = 9'b111111111;
assign micromat[84][14] = 9'b111111111;
assign micromat[84][15] = 9'b111111111;
assign micromat[84][16] = 9'b111111111;
assign micromat[84][17] = 9'b111111111;
assign micromat[84][18] = 9'b111111111;
assign micromat[84][19] = 9'b111111111;
assign micromat[84][20] = 9'b111111111;
assign micromat[84][21] = 9'b111111111;
assign micromat[84][22] = 9'b111111111;
assign micromat[84][23] = 9'b111111111;
assign micromat[84][24] = 9'b111111111;
assign micromat[84][25] = 9'b111111111;
assign micromat[84][26] = 9'b111111111;
assign micromat[84][27] = 9'b111111111;
assign micromat[84][28] = 9'b111111111;
assign micromat[84][29] = 9'b111111111;
assign micromat[84][30] = 9'b111111111;
assign micromat[84][31] = 9'b111111111;
assign micromat[84][32] = 9'b111111111;
assign micromat[84][33] = 9'b111111111;
assign micromat[84][34] = 9'b111111111;
assign micromat[84][35] = 9'b111111111;
assign micromat[84][36] = 9'b111111111;
assign micromat[84][37] = 9'b111111111;
assign micromat[84][38] = 9'b111111111;
assign micromat[84][39] = 9'b111111111;
assign micromat[84][40] = 9'b111111111;
assign micromat[84][41] = 9'b111111111;
assign micromat[84][42] = 9'b111111111;
assign micromat[84][43] = 9'b111111111;
assign micromat[84][44] = 9'b111111111;
assign micromat[84][45] = 9'b111111111;
assign micromat[84][46] = 9'b111111111;
assign micromat[84][47] = 9'b111111111;
assign micromat[84][48] = 9'b111111111;
assign micromat[84][49] = 9'b111111111;
assign micromat[84][50] = 9'b111111111;
assign micromat[84][51] = 9'b111111111;
assign micromat[84][52] = 9'b111111111;
assign micromat[84][53] = 9'b111111111;
assign micromat[84][54] = 9'b111111111;
assign micromat[84][55] = 9'b111111111;
assign micromat[84][56] = 9'b111111111;
assign micromat[84][57] = 9'b111111111;
assign micromat[84][58] = 9'b111111111;
assign micromat[84][59] = 9'b111111111;
assign micromat[84][60] = 9'b111111111;
assign micromat[84][61] = 9'b111111111;
assign micromat[84][62] = 9'b111111111;
assign micromat[84][63] = 9'b111111111;
assign micromat[84][64] = 9'b111111111;
assign micromat[84][65] = 9'b111111111;
assign micromat[84][66] = 9'b111111111;
assign micromat[84][67] = 9'b111111111;
assign micromat[84][68] = 9'b111111111;
assign micromat[84][69] = 9'b111111111;
assign micromat[84][70] = 9'b111111111;
assign micromat[84][71] = 9'b111111111;
assign micromat[84][72] = 9'b111111111;
assign micromat[84][73] = 9'b111111111;
assign micromat[84][74] = 9'b111111111;
assign micromat[84][75] = 9'b111111111;
assign micromat[84][76] = 9'b111111111;
assign micromat[84][77] = 9'b111111111;
assign micromat[84][78] = 9'b111111111;
assign micromat[84][79] = 9'b111111111;
assign micromat[84][80] = 9'b111111111;
assign micromat[84][81] = 9'b111111111;
assign micromat[84][82] = 9'b111111111;
assign micromat[84][83] = 9'b111111111;
assign micromat[84][84] = 9'b111111111;
assign micromat[84][85] = 9'b111111111;
assign micromat[84][86] = 9'b111111111;
assign micromat[84][87] = 9'b111111111;
assign micromat[84][88] = 9'b111111111;
assign micromat[84][89] = 9'b111111111;
assign micromat[84][90] = 9'b111111111;
assign micromat[84][91] = 9'b111111111;
assign micromat[84][92] = 9'b111111111;
assign micromat[84][93] = 9'b111111111;
assign micromat[84][94] = 9'b111111111;
assign micromat[84][95] = 9'b111111111;
assign micromat[84][96] = 9'b111111111;
assign micromat[84][97] = 9'b111111111;
assign micromat[84][98] = 9'b111111111;
assign micromat[84][99] = 9'b111111111;
assign micromat[85][0] = 9'b111111111;
assign micromat[85][1] = 9'b111111111;
assign micromat[85][2] = 9'b111111111;
assign micromat[85][3] = 9'b111111111;
assign micromat[85][4] = 9'b111111111;
assign micromat[85][5] = 9'b111111111;
assign micromat[85][6] = 9'b111111111;
assign micromat[85][7] = 9'b111111111;
assign micromat[85][8] = 9'b111111111;
assign micromat[85][9] = 9'b111111111;
assign micromat[85][10] = 9'b111111111;
assign micromat[85][11] = 9'b111111111;
assign micromat[85][12] = 9'b111111111;
assign micromat[85][13] = 9'b111111111;
assign micromat[85][14] = 9'b111111111;
assign micromat[85][15] = 9'b111111111;
assign micromat[85][16] = 9'b111111111;
assign micromat[85][17] = 9'b111111111;
assign micromat[85][18] = 9'b111111111;
assign micromat[85][19] = 9'b111111111;
assign micromat[85][20] = 9'b111111111;
assign micromat[85][21] = 9'b111111111;
assign micromat[85][22] = 9'b111111111;
assign micromat[85][23] = 9'b111111111;
assign micromat[85][24] = 9'b111111111;
assign micromat[85][25] = 9'b111111111;
assign micromat[85][26] = 9'b111111111;
assign micromat[85][27] = 9'b111111111;
assign micromat[85][28] = 9'b111111111;
assign micromat[85][29] = 9'b111111111;
assign micromat[85][30] = 9'b111111111;
assign micromat[85][31] = 9'b111111111;
assign micromat[85][32] = 9'b111111111;
assign micromat[85][33] = 9'b111111111;
assign micromat[85][34] = 9'b111111111;
assign micromat[85][35] = 9'b111111111;
assign micromat[85][36] = 9'b111111111;
assign micromat[85][37] = 9'b111111111;
assign micromat[85][38] = 9'b111111111;
assign micromat[85][39] = 9'b111111111;
assign micromat[85][40] = 9'b111111111;
assign micromat[85][41] = 9'b111111111;
assign micromat[85][42] = 9'b111111111;
assign micromat[85][43] = 9'b111111111;
assign micromat[85][44] = 9'b111111111;
assign micromat[85][45] = 9'b111111111;
assign micromat[85][46] = 9'b111111111;
assign micromat[85][47] = 9'b111111111;
assign micromat[85][48] = 9'b111111111;
assign micromat[85][49] = 9'b111111111;
assign micromat[85][50] = 9'b111111111;
assign micromat[85][51] = 9'b111111111;
assign micromat[85][52] = 9'b111111111;
assign micromat[85][53] = 9'b111111111;
assign micromat[85][54] = 9'b111111111;
assign micromat[85][55] = 9'b111111111;
assign micromat[85][56] = 9'b111111111;
assign micromat[85][57] = 9'b111111111;
assign micromat[85][58] = 9'b111111111;
assign micromat[85][59] = 9'b111111111;
assign micromat[85][60] = 9'b111111111;
assign micromat[85][61] = 9'b111111111;
assign micromat[85][62] = 9'b111111111;
assign micromat[85][63] = 9'b111111111;
assign micromat[85][64] = 9'b111111111;
assign micromat[85][65] = 9'b111111111;
assign micromat[85][66] = 9'b111111111;
assign micromat[85][67] = 9'b111111111;
assign micromat[85][68] = 9'b111111111;
assign micromat[85][69] = 9'b111111111;
assign micromat[85][70] = 9'b111111111;
assign micromat[85][71] = 9'b111111111;
assign micromat[85][72] = 9'b111111111;
assign micromat[85][73] = 9'b111111111;
assign micromat[85][74] = 9'b111111111;
assign micromat[85][75] = 9'b111111111;
assign micromat[85][76] = 9'b111111111;
assign micromat[85][77] = 9'b111111111;
assign micromat[85][78] = 9'b111111111;
assign micromat[85][79] = 9'b111111111;
assign micromat[85][80] = 9'b111111111;
assign micromat[85][81] = 9'b111111111;
assign micromat[85][82] = 9'b111111111;
assign micromat[85][83] = 9'b111111111;
assign micromat[85][84] = 9'b111111111;
assign micromat[85][85] = 9'b111111111;
assign micromat[85][86] = 9'b111111111;
assign micromat[85][87] = 9'b111111111;
assign micromat[85][88] = 9'b111111111;
assign micromat[85][89] = 9'b111111111;
assign micromat[85][90] = 9'b111111111;
assign micromat[85][91] = 9'b111111111;
assign micromat[85][92] = 9'b111111111;
assign micromat[85][93] = 9'b111111111;
assign micromat[85][94] = 9'b111111111;
assign micromat[85][95] = 9'b111111111;
assign micromat[85][96] = 9'b111111111;
assign micromat[85][97] = 9'b111111111;
assign micromat[85][98] = 9'b111111111;
assign micromat[85][99] = 9'b111111111;
assign micromat[86][0] = 9'b111111111;
assign micromat[86][1] = 9'b111111111;
assign micromat[86][2] = 9'b111111111;
assign micromat[86][3] = 9'b111111111;
assign micromat[86][4] = 9'b111111111;
assign micromat[86][5] = 9'b111111111;
assign micromat[86][6] = 9'b111111111;
assign micromat[86][7] = 9'b111111111;
assign micromat[86][8] = 9'b111111111;
assign micromat[86][9] = 9'b111111111;
assign micromat[86][10] = 9'b111111111;
assign micromat[86][11] = 9'b111111111;
assign micromat[86][12] = 9'b111111111;
assign micromat[86][13] = 9'b111111111;
assign micromat[86][14] = 9'b111111111;
assign micromat[86][15] = 9'b111111111;
assign micromat[86][16] = 9'b111111111;
assign micromat[86][17] = 9'b111111111;
assign micromat[86][18] = 9'b111111111;
assign micromat[86][19] = 9'b111111111;
assign micromat[86][20] = 9'b111111111;
assign micromat[86][21] = 9'b111111111;
assign micromat[86][22] = 9'b111111111;
assign micromat[86][23] = 9'b111111111;
assign micromat[86][24] = 9'b111111111;
assign micromat[86][25] = 9'b111111111;
assign micromat[86][26] = 9'b111111111;
assign micromat[86][27] = 9'b111111111;
assign micromat[86][28] = 9'b111111111;
assign micromat[86][29] = 9'b111111111;
assign micromat[86][30] = 9'b111111111;
assign micromat[86][31] = 9'b111111111;
assign micromat[86][32] = 9'b111111111;
assign micromat[86][33] = 9'b111111111;
assign micromat[86][34] = 9'b111111111;
assign micromat[86][35] = 9'b111111111;
assign micromat[86][36] = 9'b111111111;
assign micromat[86][37] = 9'b111111111;
assign micromat[86][38] = 9'b111111111;
assign micromat[86][39] = 9'b111111111;
assign micromat[86][40] = 9'b111111111;
assign micromat[86][41] = 9'b111111111;
assign micromat[86][42] = 9'b111111111;
assign micromat[86][43] = 9'b111111111;
assign micromat[86][44] = 9'b111111111;
assign micromat[86][45] = 9'b111111111;
assign micromat[86][46] = 9'b111111111;
assign micromat[86][47] = 9'b111111111;
assign micromat[86][48] = 9'b111111111;
assign micromat[86][49] = 9'b111111111;
assign micromat[86][50] = 9'b111111111;
assign micromat[86][51] = 9'b111111111;
assign micromat[86][52] = 9'b111111111;
assign micromat[86][53] = 9'b111111111;
assign micromat[86][54] = 9'b111111111;
assign micromat[86][55] = 9'b111111111;
assign micromat[86][56] = 9'b111111111;
assign micromat[86][57] = 9'b111111111;
assign micromat[86][58] = 9'b111111111;
assign micromat[86][59] = 9'b111111111;
assign micromat[86][60] = 9'b111111111;
assign micromat[86][61] = 9'b111111111;
assign micromat[86][62] = 9'b111111111;
assign micromat[86][63] = 9'b111111111;
assign micromat[86][64] = 9'b111111111;
assign micromat[86][65] = 9'b111111111;
assign micromat[86][66] = 9'b111111111;
assign micromat[86][67] = 9'b111111111;
assign micromat[86][68] = 9'b111111111;
assign micromat[86][69] = 9'b111111111;
assign micromat[86][70] = 9'b111111111;
assign micromat[86][71] = 9'b111111111;
assign micromat[86][72] = 9'b111111111;
assign micromat[86][73] = 9'b111111111;
assign micromat[86][74] = 9'b111111111;
assign micromat[86][75] = 9'b111111111;
assign micromat[86][76] = 9'b111111111;
assign micromat[86][77] = 9'b111111111;
assign micromat[86][78] = 9'b111111111;
assign micromat[86][79] = 9'b111111111;
assign micromat[86][80] = 9'b111111111;
assign micromat[86][81] = 9'b111111111;
assign micromat[86][82] = 9'b111111111;
assign micromat[86][83] = 9'b111111111;
assign micromat[86][84] = 9'b111111111;
assign micromat[86][85] = 9'b111111111;
assign micromat[86][86] = 9'b111111111;
assign micromat[86][87] = 9'b111111111;
assign micromat[86][88] = 9'b111111111;
assign micromat[86][89] = 9'b111111111;
assign micromat[86][90] = 9'b111111111;
assign micromat[86][91] = 9'b111111111;
assign micromat[86][92] = 9'b111111111;
assign micromat[86][93] = 9'b111111111;
assign micromat[86][94] = 9'b111111111;
assign micromat[86][95] = 9'b111111111;
assign micromat[86][96] = 9'b111111111;
assign micromat[86][97] = 9'b111111111;
assign micromat[86][98] = 9'b111111111;
assign micromat[86][99] = 9'b111111111;
assign micromat[87][0] = 9'b111111111;
assign micromat[87][1] = 9'b111111111;
assign micromat[87][2] = 9'b111111111;
assign micromat[87][3] = 9'b111111111;
assign micromat[87][4] = 9'b111111111;
assign micromat[87][5] = 9'b111111111;
assign micromat[87][6] = 9'b111111111;
assign micromat[87][7] = 9'b111111111;
assign micromat[87][8] = 9'b111111111;
assign micromat[87][9] = 9'b111111111;
assign micromat[87][10] = 9'b111111111;
assign micromat[87][11] = 9'b111111111;
assign micromat[87][12] = 9'b111111111;
assign micromat[87][13] = 9'b111111111;
assign micromat[87][14] = 9'b111111111;
assign micromat[87][15] = 9'b111111111;
assign micromat[87][16] = 9'b111111111;
assign micromat[87][17] = 9'b111111111;
assign micromat[87][18] = 9'b111111111;
assign micromat[87][19] = 9'b111111111;
assign micromat[87][20] = 9'b111111111;
assign micromat[87][21] = 9'b111111111;
assign micromat[87][22] = 9'b111111111;
assign micromat[87][23] = 9'b111111111;
assign micromat[87][24] = 9'b111111111;
assign micromat[87][25] = 9'b111111111;
assign micromat[87][26] = 9'b111111111;
assign micromat[87][27] = 9'b111111111;
assign micromat[87][28] = 9'b111111111;
assign micromat[87][29] = 9'b111111111;
assign micromat[87][30] = 9'b111111111;
assign micromat[87][31] = 9'b111111111;
assign micromat[87][32] = 9'b111111111;
assign micromat[87][33] = 9'b111111111;
assign micromat[87][34] = 9'b111111111;
assign micromat[87][35] = 9'b111111111;
assign micromat[87][36] = 9'b111111111;
assign micromat[87][37] = 9'b111111111;
assign micromat[87][38] = 9'b111111111;
assign micromat[87][39] = 9'b111111111;
assign micromat[87][40] = 9'b111111111;
assign micromat[87][41] = 9'b111111111;
assign micromat[87][42] = 9'b111111111;
assign micromat[87][43] = 9'b111111111;
assign micromat[87][44] = 9'b111111111;
assign micromat[87][45] = 9'b111111111;
assign micromat[87][46] = 9'b111111111;
assign micromat[87][47] = 9'b111111111;
assign micromat[87][48] = 9'b111111111;
assign micromat[87][49] = 9'b111111111;
assign micromat[87][50] = 9'b111111111;
assign micromat[87][51] = 9'b111111111;
assign micromat[87][52] = 9'b111111111;
assign micromat[87][53] = 9'b111111111;
assign micromat[87][54] = 9'b111111111;
assign micromat[87][55] = 9'b111111111;
assign micromat[87][56] = 9'b111111111;
assign micromat[87][57] = 9'b111111111;
assign micromat[87][58] = 9'b111111111;
assign micromat[87][59] = 9'b111111111;
assign micromat[87][60] = 9'b111111111;
assign micromat[87][61] = 9'b111111111;
assign micromat[87][62] = 9'b111111111;
assign micromat[87][63] = 9'b111111111;
assign micromat[87][64] = 9'b111111111;
assign micromat[87][65] = 9'b111111111;
assign micromat[87][66] = 9'b111111111;
assign micromat[87][67] = 9'b111111111;
assign micromat[87][68] = 9'b111111111;
assign micromat[87][69] = 9'b111111111;
assign micromat[87][70] = 9'b111111111;
assign micromat[87][71] = 9'b111111111;
assign micromat[87][72] = 9'b111111111;
assign micromat[87][73] = 9'b111111111;
assign micromat[87][74] = 9'b111111111;
assign micromat[87][75] = 9'b111111111;
assign micromat[87][76] = 9'b111111111;
assign micromat[87][77] = 9'b111111111;
assign micromat[87][78] = 9'b111111111;
assign micromat[87][79] = 9'b111111111;
assign micromat[87][80] = 9'b111111111;
assign micromat[87][81] = 9'b111111111;
assign micromat[87][82] = 9'b111111111;
assign micromat[87][83] = 9'b111111111;
assign micromat[87][84] = 9'b111111111;
assign micromat[87][85] = 9'b111111111;
assign micromat[87][86] = 9'b111111111;
assign micromat[87][87] = 9'b111111111;
assign micromat[87][88] = 9'b111111111;
assign micromat[87][89] = 9'b111111111;
assign micromat[87][90] = 9'b111111111;
assign micromat[87][91] = 9'b111111111;
assign micromat[87][92] = 9'b111111111;
assign micromat[87][93] = 9'b111111111;
assign micromat[87][94] = 9'b111111111;
assign micromat[87][95] = 9'b111111111;
assign micromat[87][96] = 9'b111111111;
assign micromat[87][97] = 9'b111111111;
assign micromat[87][98] = 9'b111111111;
assign micromat[87][99] = 9'b111111111;
assign micromat[88][0] = 9'b111111111;
assign micromat[88][1] = 9'b111111111;
assign micromat[88][2] = 9'b111111111;
assign micromat[88][3] = 9'b111111111;
assign micromat[88][4] = 9'b111111111;
assign micromat[88][5] = 9'b111111111;
assign micromat[88][6] = 9'b111111111;
assign micromat[88][7] = 9'b111111111;
assign micromat[88][8] = 9'b111111111;
assign micromat[88][9] = 9'b111111111;
assign micromat[88][10] = 9'b111111111;
assign micromat[88][11] = 9'b111111111;
assign micromat[88][12] = 9'b111111111;
assign micromat[88][13] = 9'b111111111;
assign micromat[88][14] = 9'b111111111;
assign micromat[88][15] = 9'b111111111;
assign micromat[88][16] = 9'b111111111;
assign micromat[88][17] = 9'b111111111;
assign micromat[88][18] = 9'b111111111;
assign micromat[88][19] = 9'b111111111;
assign micromat[88][20] = 9'b111111111;
assign micromat[88][21] = 9'b111111111;
assign micromat[88][22] = 9'b111111111;
assign micromat[88][23] = 9'b111111111;
assign micromat[88][24] = 9'b111111111;
assign micromat[88][25] = 9'b111111111;
assign micromat[88][26] = 9'b111111111;
assign micromat[88][27] = 9'b111111111;
assign micromat[88][28] = 9'b111111111;
assign micromat[88][29] = 9'b111111111;
assign micromat[88][30] = 9'b111111111;
assign micromat[88][31] = 9'b111111111;
assign micromat[88][32] = 9'b111111111;
assign micromat[88][33] = 9'b111111111;
assign micromat[88][34] = 9'b111111111;
assign micromat[88][35] = 9'b111111111;
assign micromat[88][36] = 9'b111111111;
assign micromat[88][37] = 9'b111111111;
assign micromat[88][38] = 9'b111111111;
assign micromat[88][39] = 9'b111111111;
assign micromat[88][40] = 9'b111111111;
assign micromat[88][41] = 9'b111111111;
assign micromat[88][42] = 9'b111111111;
assign micromat[88][43] = 9'b111111111;
assign micromat[88][44] = 9'b111111111;
assign micromat[88][45] = 9'b111111111;
assign micromat[88][46] = 9'b111111111;
assign micromat[88][47] = 9'b111111111;
assign micromat[88][48] = 9'b111111111;
assign micromat[88][49] = 9'b111111111;
assign micromat[88][50] = 9'b111111111;
assign micromat[88][51] = 9'b111111111;
assign micromat[88][52] = 9'b111111111;
assign micromat[88][53] = 9'b111111111;
assign micromat[88][54] = 9'b111111111;
assign micromat[88][55] = 9'b111111111;
assign micromat[88][56] = 9'b111111111;
assign micromat[88][57] = 9'b111111111;
assign micromat[88][58] = 9'b111111111;
assign micromat[88][59] = 9'b111111111;
assign micromat[88][60] = 9'b111111111;
assign micromat[88][61] = 9'b111111111;
assign micromat[88][62] = 9'b111111111;
assign micromat[88][63] = 9'b111111111;
assign micromat[88][64] = 9'b111111111;
assign micromat[88][65] = 9'b111111111;
assign micromat[88][66] = 9'b111111111;
assign micromat[88][67] = 9'b111111111;
assign micromat[88][68] = 9'b111111111;
assign micromat[88][69] = 9'b111111111;
assign micromat[88][70] = 9'b111111111;
assign micromat[88][71] = 9'b111111111;
assign micromat[88][72] = 9'b111111111;
assign micromat[88][73] = 9'b111111111;
assign micromat[88][74] = 9'b111111111;
assign micromat[88][75] = 9'b111111111;
assign micromat[88][76] = 9'b111111111;
assign micromat[88][77] = 9'b111111111;
assign micromat[88][78] = 9'b111111111;
assign micromat[88][79] = 9'b111111111;
assign micromat[88][80] = 9'b111111111;
assign micromat[88][81] = 9'b111111111;
assign micromat[88][82] = 9'b111111111;
assign micromat[88][83] = 9'b111111111;
assign micromat[88][84] = 9'b111111111;
assign micromat[88][85] = 9'b111111111;
assign micromat[88][86] = 9'b111111111;
assign micromat[88][87] = 9'b111111111;
assign micromat[88][88] = 9'b111111111;
assign micromat[88][89] = 9'b111111111;
assign micromat[88][90] = 9'b111111111;
assign micromat[88][91] = 9'b111111111;
assign micromat[88][92] = 9'b111111111;
assign micromat[88][93] = 9'b111111111;
assign micromat[88][94] = 9'b111111111;
assign micromat[88][95] = 9'b111111111;
assign micromat[88][96] = 9'b111111111;
assign micromat[88][97] = 9'b111111111;
assign micromat[88][98] = 9'b111111111;
assign micromat[88][99] = 9'b111111111;
assign micromat[89][0] = 9'b111111111;
assign micromat[89][1] = 9'b111111111;
assign micromat[89][2] = 9'b111111111;
assign micromat[89][3] = 9'b111111111;
assign micromat[89][4] = 9'b111111111;
assign micromat[89][5] = 9'b111111111;
assign micromat[89][6] = 9'b111111111;
assign micromat[89][7] = 9'b111111111;
assign micromat[89][8] = 9'b111111111;
assign micromat[89][9] = 9'b111111111;
assign micromat[89][10] = 9'b111111111;
assign micromat[89][11] = 9'b111111111;
assign micromat[89][12] = 9'b111111111;
assign micromat[89][13] = 9'b111111111;
assign micromat[89][14] = 9'b111111111;
assign micromat[89][15] = 9'b111111111;
assign micromat[89][16] = 9'b111111111;
assign micromat[89][17] = 9'b111111111;
assign micromat[89][18] = 9'b111111111;
assign micromat[89][19] = 9'b111111111;
assign micromat[89][20] = 9'b111111111;
assign micromat[89][21] = 9'b111111111;
assign micromat[89][22] = 9'b111111111;
assign micromat[89][23] = 9'b111111111;
assign micromat[89][24] = 9'b111111111;
assign micromat[89][25] = 9'b111111111;
assign micromat[89][26] = 9'b111111111;
assign micromat[89][27] = 9'b111111111;
assign micromat[89][28] = 9'b111111111;
assign micromat[89][29] = 9'b111111111;
assign micromat[89][30] = 9'b111111111;
assign micromat[89][31] = 9'b111111111;
assign micromat[89][32] = 9'b111111111;
assign micromat[89][33] = 9'b111111111;
assign micromat[89][34] = 9'b111111111;
assign micromat[89][35] = 9'b111111111;
assign micromat[89][36] = 9'b111111111;
assign micromat[89][37] = 9'b111111111;
assign micromat[89][38] = 9'b111111111;
assign micromat[89][39] = 9'b111111111;
assign micromat[89][40] = 9'b111111111;
assign micromat[89][41] = 9'b111111111;
assign micromat[89][42] = 9'b111111111;
assign micromat[89][43] = 9'b111111111;
assign micromat[89][44] = 9'b111111111;
assign micromat[89][45] = 9'b111111111;
assign micromat[89][46] = 9'b111111111;
assign micromat[89][47] = 9'b111111111;
assign micromat[89][48] = 9'b111111111;
assign micromat[89][49] = 9'b111111111;
assign micromat[89][50] = 9'b111111111;
assign micromat[89][51] = 9'b111111111;
assign micromat[89][52] = 9'b111111111;
assign micromat[89][53] = 9'b111111111;
assign micromat[89][54] = 9'b111111111;
assign micromat[89][55] = 9'b111111111;
assign micromat[89][56] = 9'b111111111;
assign micromat[89][57] = 9'b111111111;
assign micromat[89][58] = 9'b111111111;
assign micromat[89][59] = 9'b111111111;
assign micromat[89][60] = 9'b111111111;
assign micromat[89][61] = 9'b111111111;
assign micromat[89][62] = 9'b111111111;
assign micromat[89][63] = 9'b111111111;
assign micromat[89][64] = 9'b111111111;
assign micromat[89][65] = 9'b111111111;
assign micromat[89][66] = 9'b111111111;
assign micromat[89][67] = 9'b111111111;
assign micromat[89][68] = 9'b111111111;
assign micromat[89][69] = 9'b111111111;
assign micromat[89][70] = 9'b111111111;
assign micromat[89][71] = 9'b111111111;
assign micromat[89][72] = 9'b111111111;
assign micromat[89][73] = 9'b111111111;
assign micromat[89][74] = 9'b111111111;
assign micromat[89][75] = 9'b111111111;
assign micromat[89][76] = 9'b111111111;
assign micromat[89][77] = 9'b111111111;
assign micromat[89][78] = 9'b111111111;
assign micromat[89][79] = 9'b111111111;
assign micromat[89][80] = 9'b111111111;
assign micromat[89][81] = 9'b111111111;
assign micromat[89][82] = 9'b111111111;
assign micromat[89][83] = 9'b111111111;
assign micromat[89][84] = 9'b111111111;
assign micromat[89][85] = 9'b111111111;
assign micromat[89][86] = 9'b111111111;
assign micromat[89][87] = 9'b111111111;
assign micromat[89][88] = 9'b111111111;
assign micromat[89][89] = 9'b111111111;
assign micromat[89][90] = 9'b111111111;
assign micromat[89][91] = 9'b111111111;
assign micromat[89][92] = 9'b111111111;
assign micromat[89][93] = 9'b111111111;
assign micromat[89][94] = 9'b111111111;
assign micromat[89][95] = 9'b111111111;
assign micromat[89][96] = 9'b111111111;
assign micromat[89][97] = 9'b111111111;
assign micromat[89][98] = 9'b111111111;
assign micromat[89][99] = 9'b111111111;
assign micromat[90][0] = 9'b111111111;
assign micromat[90][1] = 9'b111111111;
assign micromat[90][2] = 9'b111111111;
assign micromat[90][3] = 9'b111111111;
assign micromat[90][4] = 9'b111111111;
assign micromat[90][5] = 9'b111111111;
assign micromat[90][6] = 9'b111111111;
assign micromat[90][7] = 9'b111111111;
assign micromat[90][8] = 9'b111111111;
assign micromat[90][9] = 9'b111111111;
assign micromat[90][10] = 9'b111111111;
assign micromat[90][11] = 9'b111111111;
assign micromat[90][12] = 9'b111111111;
assign micromat[90][13] = 9'b111111111;
assign micromat[90][14] = 9'b111111111;
assign micromat[90][15] = 9'b111111111;
assign micromat[90][16] = 9'b111111111;
assign micromat[90][17] = 9'b111111111;
assign micromat[90][18] = 9'b111111111;
assign micromat[90][19] = 9'b111111111;
assign micromat[90][20] = 9'b111111111;
assign micromat[90][21] = 9'b111111111;
assign micromat[90][22] = 9'b111111111;
assign micromat[90][23] = 9'b111111111;
assign micromat[90][24] = 9'b111111111;
assign micromat[90][25] = 9'b111111111;
assign micromat[90][26] = 9'b111111111;
assign micromat[90][27] = 9'b111111111;
assign micromat[90][28] = 9'b111111111;
assign micromat[90][29] = 9'b111111111;
assign micromat[90][30] = 9'b111111111;
assign micromat[90][31] = 9'b111111111;
assign micromat[90][32] = 9'b111111111;
assign micromat[90][33] = 9'b111111111;
assign micromat[90][34] = 9'b111111111;
assign micromat[90][35] = 9'b111111111;
assign micromat[90][36] = 9'b111111111;
assign micromat[90][37] = 9'b111111111;
assign micromat[90][38] = 9'b111111111;
assign micromat[90][39] = 9'b111111111;
assign micromat[90][40] = 9'b111111111;
assign micromat[90][41] = 9'b111111111;
assign micromat[90][42] = 9'b111111111;
assign micromat[90][43] = 9'b111111111;
assign micromat[90][44] = 9'b111111111;
assign micromat[90][45] = 9'b111111111;
assign micromat[90][46] = 9'b111111111;
assign micromat[90][47] = 9'b111111111;
assign micromat[90][48] = 9'b111111111;
assign micromat[90][49] = 9'b111111111;
assign micromat[90][50] = 9'b111111111;
assign micromat[90][51] = 9'b111111111;
assign micromat[90][52] = 9'b111111111;
assign micromat[90][53] = 9'b111111111;
assign micromat[90][54] = 9'b111111111;
assign micromat[90][55] = 9'b111111111;
assign micromat[90][56] = 9'b111111111;
assign micromat[90][57] = 9'b111111111;
assign micromat[90][58] = 9'b111111111;
assign micromat[90][59] = 9'b111111111;
assign micromat[90][60] = 9'b111111111;
assign micromat[90][61] = 9'b111111111;
assign micromat[90][62] = 9'b111111111;
assign micromat[90][63] = 9'b111111111;
assign micromat[90][64] = 9'b111111111;
assign micromat[90][65] = 9'b111111111;
assign micromat[90][66] = 9'b111111111;
assign micromat[90][67] = 9'b111111111;
assign micromat[90][68] = 9'b111111111;
assign micromat[90][69] = 9'b111111111;
assign micromat[90][70] = 9'b111111111;
assign micromat[90][71] = 9'b111111111;
assign micromat[90][72] = 9'b111111111;
assign micromat[90][73] = 9'b111111111;
assign micromat[90][74] = 9'b111111111;
assign micromat[90][75] = 9'b111111111;
assign micromat[90][76] = 9'b111111111;
assign micromat[90][77] = 9'b111111111;
assign micromat[90][78] = 9'b111111111;
assign micromat[90][79] = 9'b111111111;
assign micromat[90][80] = 9'b111111111;
assign micromat[90][81] = 9'b111111111;
assign micromat[90][82] = 9'b111111111;
assign micromat[90][83] = 9'b111111111;
assign micromat[90][84] = 9'b111111111;
assign micromat[90][85] = 9'b111111111;
assign micromat[90][86] = 9'b111111111;
assign micromat[90][87] = 9'b111111111;
assign micromat[90][88] = 9'b111111111;
assign micromat[90][89] = 9'b111111111;
assign micromat[90][90] = 9'b111111111;
assign micromat[90][91] = 9'b111111111;
assign micromat[90][92] = 9'b111111111;
assign micromat[90][93] = 9'b111111111;
assign micromat[90][94] = 9'b111111111;
assign micromat[90][95] = 9'b111111111;
assign micromat[90][96] = 9'b111111111;
assign micromat[90][97] = 9'b111111111;
assign micromat[90][98] = 9'b111111111;
assign micromat[90][99] = 9'b111111111;
assign micromat[91][0] = 9'b111111111;
assign micromat[91][1] = 9'b111111111;
assign micromat[91][2] = 9'b111111111;
assign micromat[91][3] = 9'b111111111;
assign micromat[91][4] = 9'b111111111;
assign micromat[91][5] = 9'b111111111;
assign micromat[91][6] = 9'b111111111;
assign micromat[91][7] = 9'b111111111;
assign micromat[91][8] = 9'b111111111;
assign micromat[91][9] = 9'b111111111;
assign micromat[91][10] = 9'b111111111;
assign micromat[91][11] = 9'b111111111;
assign micromat[91][12] = 9'b111111111;
assign micromat[91][13] = 9'b111111111;
assign micromat[91][14] = 9'b111111111;
assign micromat[91][15] = 9'b111111111;
assign micromat[91][16] = 9'b111111111;
assign micromat[91][17] = 9'b111111111;
assign micromat[91][18] = 9'b111111111;
assign micromat[91][19] = 9'b111111111;
assign micromat[91][20] = 9'b111111111;
assign micromat[91][21] = 9'b111111111;
assign micromat[91][22] = 9'b111111111;
assign micromat[91][23] = 9'b111111111;
assign micromat[91][24] = 9'b111111111;
assign micromat[91][25] = 9'b111111111;
assign micromat[91][26] = 9'b111111111;
assign micromat[91][27] = 9'b111111111;
assign micromat[91][28] = 9'b111111111;
assign micromat[91][29] = 9'b111111111;
assign micromat[91][30] = 9'b111111111;
assign micromat[91][31] = 9'b111111111;
assign micromat[91][32] = 9'b111111111;
assign micromat[91][33] = 9'b111111111;
assign micromat[91][34] = 9'b111111111;
assign micromat[91][35] = 9'b111111111;
assign micromat[91][36] = 9'b111111111;
assign micromat[91][37] = 9'b111111111;
assign micromat[91][38] = 9'b111111111;
assign micromat[91][39] = 9'b111111111;
assign micromat[91][40] = 9'b111111111;
assign micromat[91][41] = 9'b111111111;
assign micromat[91][42] = 9'b111111111;
assign micromat[91][43] = 9'b111111111;
assign micromat[91][44] = 9'b111111111;
assign micromat[91][45] = 9'b111111111;
assign micromat[91][46] = 9'b111111111;
assign micromat[91][47] = 9'b111111111;
assign micromat[91][48] = 9'b111111111;
assign micromat[91][49] = 9'b111111111;
assign micromat[91][50] = 9'b111111111;
assign micromat[91][51] = 9'b111111111;
assign micromat[91][52] = 9'b111111111;
assign micromat[91][53] = 9'b111111111;
assign micromat[91][54] = 9'b111111111;
assign micromat[91][55] = 9'b111111111;
assign micromat[91][56] = 9'b111111111;
assign micromat[91][57] = 9'b111111111;
assign micromat[91][58] = 9'b111111111;
assign micromat[91][59] = 9'b111111111;
assign micromat[91][60] = 9'b111111111;
assign micromat[91][61] = 9'b111111111;
assign micromat[91][62] = 9'b111111111;
assign micromat[91][63] = 9'b111111111;
assign micromat[91][64] = 9'b111111111;
assign micromat[91][65] = 9'b111111111;
assign micromat[91][66] = 9'b111111111;
assign micromat[91][67] = 9'b111111111;
assign micromat[91][68] = 9'b111111111;
assign micromat[91][69] = 9'b111111111;
assign micromat[91][70] = 9'b111111111;
assign micromat[91][71] = 9'b111111111;
assign micromat[91][72] = 9'b111111111;
assign micromat[91][73] = 9'b111111111;
assign micromat[91][74] = 9'b111111111;
assign micromat[91][75] = 9'b111111111;
assign micromat[91][76] = 9'b111111111;
assign micromat[91][77] = 9'b111111111;
assign micromat[91][78] = 9'b111111111;
assign micromat[91][79] = 9'b111111111;
assign micromat[91][80] = 9'b111111111;
assign micromat[91][81] = 9'b111111111;
assign micromat[91][82] = 9'b111111111;
assign micromat[91][83] = 9'b111111111;
assign micromat[91][84] = 9'b111111111;
assign micromat[91][85] = 9'b111111111;
assign micromat[91][86] = 9'b111111111;
assign micromat[91][87] = 9'b111111111;
assign micromat[91][88] = 9'b111111111;
assign micromat[91][89] = 9'b111111111;
assign micromat[91][90] = 9'b111111111;
assign micromat[91][91] = 9'b111111111;
assign micromat[91][92] = 9'b111111111;
assign micromat[91][93] = 9'b111111111;
assign micromat[91][94] = 9'b111111111;
assign micromat[91][95] = 9'b111111111;
assign micromat[91][96] = 9'b111111111;
assign micromat[91][97] = 9'b111111111;
assign micromat[91][98] = 9'b111111111;
assign micromat[91][99] = 9'b111111111;
assign micromat[92][0] = 9'b111111111;
assign micromat[92][1] = 9'b111111111;
assign micromat[92][2] = 9'b111111111;
assign micromat[92][3] = 9'b111111111;
assign micromat[92][4] = 9'b111111111;
assign micromat[92][5] = 9'b111111111;
assign micromat[92][6] = 9'b111111111;
assign micromat[92][7] = 9'b111111111;
assign micromat[92][8] = 9'b111111111;
assign micromat[92][9] = 9'b111111111;
assign micromat[92][10] = 9'b111111111;
assign micromat[92][11] = 9'b111111111;
assign micromat[92][12] = 9'b111111111;
assign micromat[92][13] = 9'b111111111;
assign micromat[92][14] = 9'b111111111;
assign micromat[92][15] = 9'b111111111;
assign micromat[92][16] = 9'b111111111;
assign micromat[92][17] = 9'b111111111;
assign micromat[92][18] = 9'b111111111;
assign micromat[92][19] = 9'b111111111;
assign micromat[92][20] = 9'b111111111;
assign micromat[92][21] = 9'b111111111;
assign micromat[92][22] = 9'b111111111;
assign micromat[92][23] = 9'b111111111;
assign micromat[92][24] = 9'b111111111;
assign micromat[92][25] = 9'b111111111;
assign micromat[92][26] = 9'b111111111;
assign micromat[92][27] = 9'b111111111;
assign micromat[92][28] = 9'b111111111;
assign micromat[92][29] = 9'b111111111;
assign micromat[92][30] = 9'b111111111;
assign micromat[92][31] = 9'b111111111;
assign micromat[92][32] = 9'b111111111;
assign micromat[92][33] = 9'b111111111;
assign micromat[92][34] = 9'b111111111;
assign micromat[92][35] = 9'b111111111;
assign micromat[92][36] = 9'b111111111;
assign micromat[92][37] = 9'b111111111;
assign micromat[92][38] = 9'b111111111;
assign micromat[92][39] = 9'b111111111;
assign micromat[92][40] = 9'b111111111;
assign micromat[92][41] = 9'b111111111;
assign micromat[92][42] = 9'b111111111;
assign micromat[92][43] = 9'b111111111;
assign micromat[92][44] = 9'b111111111;
assign micromat[92][45] = 9'b111111111;
assign micromat[92][46] = 9'b111111111;
assign micromat[92][47] = 9'b111111111;
assign micromat[92][48] = 9'b111111111;
assign micromat[92][49] = 9'b111111111;
assign micromat[92][50] = 9'b111111111;
assign micromat[92][51] = 9'b111111111;
assign micromat[92][52] = 9'b111111111;
assign micromat[92][53] = 9'b111111111;
assign micromat[92][54] = 9'b111111111;
assign micromat[92][55] = 9'b111111111;
assign micromat[92][56] = 9'b111111111;
assign micromat[92][57] = 9'b111111111;
assign micromat[92][58] = 9'b111111111;
assign micromat[92][59] = 9'b111111111;
assign micromat[92][60] = 9'b111111111;
assign micromat[92][61] = 9'b111111111;
assign micromat[92][62] = 9'b111111111;
assign micromat[92][63] = 9'b111111111;
assign micromat[92][64] = 9'b111111111;
assign micromat[92][65] = 9'b111111111;
assign micromat[92][66] = 9'b111111111;
assign micromat[92][67] = 9'b111111111;
assign micromat[92][68] = 9'b111111111;
assign micromat[92][69] = 9'b111111111;
assign micromat[92][70] = 9'b111111111;
assign micromat[92][71] = 9'b111111111;
assign micromat[92][72] = 9'b111111111;
assign micromat[92][73] = 9'b111111111;
assign micromat[92][74] = 9'b111111111;
assign micromat[92][75] = 9'b111111111;
assign micromat[92][76] = 9'b111111111;
assign micromat[92][77] = 9'b111111111;
assign micromat[92][78] = 9'b111111111;
assign micromat[92][79] = 9'b111111111;
assign micromat[92][80] = 9'b111111111;
assign micromat[92][81] = 9'b111111111;
assign micromat[92][82] = 9'b111111111;
assign micromat[92][83] = 9'b111111111;
assign micromat[92][84] = 9'b111111111;
assign micromat[92][85] = 9'b111111111;
assign micromat[92][86] = 9'b111111111;
assign micromat[92][87] = 9'b111111111;
assign micromat[92][88] = 9'b111111111;
assign micromat[92][89] = 9'b111111111;
assign micromat[92][90] = 9'b111111111;
assign micromat[92][91] = 9'b111111111;
assign micromat[92][92] = 9'b111111111;
assign micromat[92][93] = 9'b111111111;
assign micromat[92][94] = 9'b111111111;
assign micromat[92][95] = 9'b111111111;
assign micromat[92][96] = 9'b111111111;
assign micromat[92][97] = 9'b111111111;
assign micromat[92][98] = 9'b111111111;
assign micromat[92][99] = 9'b111111111;
assign micromat[93][0] = 9'b111111111;
assign micromat[93][1] = 9'b111111111;
assign micromat[93][2] = 9'b111111111;
assign micromat[93][3] = 9'b111111111;
assign micromat[93][4] = 9'b111111111;
assign micromat[93][5] = 9'b111111111;
assign micromat[93][6] = 9'b111111111;
assign micromat[93][7] = 9'b111111111;
assign micromat[93][8] = 9'b111111111;
assign micromat[93][9] = 9'b111111111;
assign micromat[93][10] = 9'b111111111;
assign micromat[93][11] = 9'b111111111;
assign micromat[93][12] = 9'b111111111;
assign micromat[93][13] = 9'b111111111;
assign micromat[93][14] = 9'b111111111;
assign micromat[93][15] = 9'b111111111;
assign micromat[93][16] = 9'b111111111;
assign micromat[93][17] = 9'b111111111;
assign micromat[93][18] = 9'b111111111;
assign micromat[93][19] = 9'b111111111;
assign micromat[93][20] = 9'b111111111;
assign micromat[93][21] = 9'b111111111;
assign micromat[93][22] = 9'b111111111;
assign micromat[93][23] = 9'b111111111;
assign micromat[93][24] = 9'b111111111;
assign micromat[93][25] = 9'b111111111;
assign micromat[93][26] = 9'b111111111;
assign micromat[93][27] = 9'b111111111;
assign micromat[93][28] = 9'b111111111;
assign micromat[93][29] = 9'b111111111;
assign micromat[93][30] = 9'b111111111;
assign micromat[93][31] = 9'b111111111;
assign micromat[93][32] = 9'b111111111;
assign micromat[93][33] = 9'b111111111;
assign micromat[93][34] = 9'b111111111;
assign micromat[93][35] = 9'b111111111;
assign micromat[93][36] = 9'b111111111;
assign micromat[93][37] = 9'b111111111;
assign micromat[93][38] = 9'b111111111;
assign micromat[93][39] = 9'b111111111;
assign micromat[93][40] = 9'b111111111;
assign micromat[93][41] = 9'b111111111;
assign micromat[93][42] = 9'b111111111;
assign micromat[93][43] = 9'b111111111;
assign micromat[93][44] = 9'b111111111;
assign micromat[93][45] = 9'b111111111;
assign micromat[93][46] = 9'b111111111;
assign micromat[93][47] = 9'b111111111;
assign micromat[93][48] = 9'b111111111;
assign micromat[93][49] = 9'b111111111;
assign micromat[93][50] = 9'b111111111;
assign micromat[93][51] = 9'b111111111;
assign micromat[93][52] = 9'b111111111;
assign micromat[93][53] = 9'b111111111;
assign micromat[93][54] = 9'b111111111;
assign micromat[93][55] = 9'b111111111;
assign micromat[93][56] = 9'b111111111;
assign micromat[93][57] = 9'b111111111;
assign micromat[93][58] = 9'b111111111;
assign micromat[93][59] = 9'b111111111;
assign micromat[93][60] = 9'b111111111;
assign micromat[93][61] = 9'b111111111;
assign micromat[93][62] = 9'b111111111;
assign micromat[93][63] = 9'b111111111;
assign micromat[93][64] = 9'b111111111;
assign micromat[93][65] = 9'b111111111;
assign micromat[93][66] = 9'b111111111;
assign micromat[93][67] = 9'b111111111;
assign micromat[93][68] = 9'b111111111;
assign micromat[93][69] = 9'b111111111;
assign micromat[93][70] = 9'b111111111;
assign micromat[93][71] = 9'b111111111;
assign micromat[93][72] = 9'b111111111;
assign micromat[93][73] = 9'b111111111;
assign micromat[93][74] = 9'b111111111;
assign micromat[93][75] = 9'b111111111;
assign micromat[93][76] = 9'b111111111;
assign micromat[93][77] = 9'b111111111;
assign micromat[93][78] = 9'b111111111;
assign micromat[93][79] = 9'b111111111;
assign micromat[93][80] = 9'b111111111;
assign micromat[93][81] = 9'b111111111;
assign micromat[93][82] = 9'b111111111;
assign micromat[93][83] = 9'b111111111;
assign micromat[93][84] = 9'b111111111;
assign micromat[93][85] = 9'b111111111;
assign micromat[93][86] = 9'b111111111;
assign micromat[93][87] = 9'b111111111;
assign micromat[93][88] = 9'b111111111;
assign micromat[93][89] = 9'b111111111;
assign micromat[93][90] = 9'b111111111;
assign micromat[93][91] = 9'b111111111;
assign micromat[93][92] = 9'b111111111;
assign micromat[93][93] = 9'b111111111;
assign micromat[93][94] = 9'b111111111;
assign micromat[93][95] = 9'b111111111;
assign micromat[93][96] = 9'b111111111;
assign micromat[93][97] = 9'b111111111;
assign micromat[93][98] = 9'b111111111;
assign micromat[93][99] = 9'b111111111;
assign micromat[94][0] = 9'b111111111;
assign micromat[94][1] = 9'b111111111;
assign micromat[94][2] = 9'b111111111;
assign micromat[94][3] = 9'b111111111;
assign micromat[94][4] = 9'b111111111;
assign micromat[94][5] = 9'b111111111;
assign micromat[94][6] = 9'b111111111;
assign micromat[94][7] = 9'b111111111;
assign micromat[94][8] = 9'b111111111;
assign micromat[94][9] = 9'b111111111;
assign micromat[94][10] = 9'b111111111;
assign micromat[94][11] = 9'b111111111;
assign micromat[94][12] = 9'b111111111;
assign micromat[94][13] = 9'b111111111;
assign micromat[94][14] = 9'b111111111;
assign micromat[94][15] = 9'b111111111;
assign micromat[94][16] = 9'b111111111;
assign micromat[94][17] = 9'b111111111;
assign micromat[94][18] = 9'b111111111;
assign micromat[94][19] = 9'b111111111;
assign micromat[94][20] = 9'b111111111;
assign micromat[94][21] = 9'b111111111;
assign micromat[94][22] = 9'b111111111;
assign micromat[94][23] = 9'b111111111;
assign micromat[94][24] = 9'b111111111;
assign micromat[94][25] = 9'b111111111;
assign micromat[94][26] = 9'b111111111;
assign micromat[94][27] = 9'b111111111;
assign micromat[94][28] = 9'b111111111;
assign micromat[94][29] = 9'b111111111;
assign micromat[94][30] = 9'b111111111;
assign micromat[94][31] = 9'b111111111;
assign micromat[94][32] = 9'b111111111;
assign micromat[94][33] = 9'b111111111;
assign micromat[94][34] = 9'b111111111;
assign micromat[94][35] = 9'b111111111;
assign micromat[94][36] = 9'b111111111;
assign micromat[94][37] = 9'b111111111;
assign micromat[94][38] = 9'b111111111;
assign micromat[94][39] = 9'b111111111;
assign micromat[94][40] = 9'b111111111;
assign micromat[94][41] = 9'b111111111;
assign micromat[94][42] = 9'b111111111;
assign micromat[94][43] = 9'b111111111;
assign micromat[94][44] = 9'b111111111;
assign micromat[94][45] = 9'b111111111;
assign micromat[94][46] = 9'b111111111;
assign micromat[94][47] = 9'b111111111;
assign micromat[94][48] = 9'b111111111;
assign micromat[94][49] = 9'b111111111;
assign micromat[94][50] = 9'b111111111;
assign micromat[94][51] = 9'b111111111;
assign micromat[94][52] = 9'b111111111;
assign micromat[94][53] = 9'b111111111;
assign micromat[94][54] = 9'b111111111;
assign micromat[94][55] = 9'b111111111;
assign micromat[94][56] = 9'b111111111;
assign micromat[94][57] = 9'b111111111;
assign micromat[94][58] = 9'b111111111;
assign micromat[94][59] = 9'b111111111;
assign micromat[94][60] = 9'b111111111;
assign micromat[94][61] = 9'b111111111;
assign micromat[94][62] = 9'b111111111;
assign micromat[94][63] = 9'b111111111;
assign micromat[94][64] = 9'b111111111;
assign micromat[94][65] = 9'b111111111;
assign micromat[94][66] = 9'b111111111;
assign micromat[94][67] = 9'b111111111;
assign micromat[94][68] = 9'b111111111;
assign micromat[94][69] = 9'b111111111;
assign micromat[94][70] = 9'b111111111;
assign micromat[94][71] = 9'b111111111;
assign micromat[94][72] = 9'b111111111;
assign micromat[94][73] = 9'b111111111;
assign micromat[94][74] = 9'b111111111;
assign micromat[94][75] = 9'b111111111;
assign micromat[94][76] = 9'b111111111;
assign micromat[94][77] = 9'b111111111;
assign micromat[94][78] = 9'b111111111;
assign micromat[94][79] = 9'b111111111;
assign micromat[94][80] = 9'b111111111;
assign micromat[94][81] = 9'b111111111;
assign micromat[94][82] = 9'b111111111;
assign micromat[94][83] = 9'b111111111;
assign micromat[94][84] = 9'b111111111;
assign micromat[94][85] = 9'b111111111;
assign micromat[94][86] = 9'b111111111;
assign micromat[94][87] = 9'b111111111;
assign micromat[94][88] = 9'b111111111;
assign micromat[94][89] = 9'b111111111;
assign micromat[94][90] = 9'b111111111;
assign micromat[94][91] = 9'b111111111;
assign micromat[94][92] = 9'b111111111;
assign micromat[94][93] = 9'b111111111;
assign micromat[94][94] = 9'b111111111;
assign micromat[94][95] = 9'b111111111;
assign micromat[94][96] = 9'b111111111;
assign micromat[94][97] = 9'b111111111;
assign micromat[94][98] = 9'b111111111;
assign micromat[94][99] = 9'b111111111;
assign micromat[95][0] = 9'b111111111;
assign micromat[95][1] = 9'b111111111;
assign micromat[95][2] = 9'b111111111;
assign micromat[95][3] = 9'b111111111;
assign micromat[95][4] = 9'b111111111;
assign micromat[95][5] = 9'b111111111;
assign micromat[95][6] = 9'b111111111;
assign micromat[95][7] = 9'b111111111;
assign micromat[95][8] = 9'b111111111;
assign micromat[95][9] = 9'b111111111;
assign micromat[95][10] = 9'b111111111;
assign micromat[95][11] = 9'b111111111;
assign micromat[95][12] = 9'b111111111;
assign micromat[95][13] = 9'b111111111;
assign micromat[95][14] = 9'b111111111;
assign micromat[95][15] = 9'b111111111;
assign micromat[95][16] = 9'b111111111;
assign micromat[95][17] = 9'b111111111;
assign micromat[95][18] = 9'b111111111;
assign micromat[95][19] = 9'b111111111;
assign micromat[95][20] = 9'b111111111;
assign micromat[95][21] = 9'b111111111;
assign micromat[95][22] = 9'b111111111;
assign micromat[95][23] = 9'b111111111;
assign micromat[95][24] = 9'b111111111;
assign micromat[95][25] = 9'b111111111;
assign micromat[95][26] = 9'b111111111;
assign micromat[95][27] = 9'b111111111;
assign micromat[95][28] = 9'b111111111;
assign micromat[95][29] = 9'b111111111;
assign micromat[95][30] = 9'b111111111;
assign micromat[95][31] = 9'b111111111;
assign micromat[95][32] = 9'b111111111;
assign micromat[95][33] = 9'b111111111;
assign micromat[95][34] = 9'b111111111;
assign micromat[95][35] = 9'b111111111;
assign micromat[95][36] = 9'b111111111;
assign micromat[95][37] = 9'b111111111;
assign micromat[95][38] = 9'b111111111;
assign micromat[95][39] = 9'b111111111;
assign micromat[95][40] = 9'b111111111;
assign micromat[95][41] = 9'b111111111;
assign micromat[95][42] = 9'b111111111;
assign micromat[95][43] = 9'b111111111;
assign micromat[95][44] = 9'b111111111;
assign micromat[95][45] = 9'b111111111;
assign micromat[95][46] = 9'b111111111;
assign micromat[95][47] = 9'b111111111;
assign micromat[95][48] = 9'b111111111;
assign micromat[95][49] = 9'b111111111;
assign micromat[95][50] = 9'b111111111;
assign micromat[95][51] = 9'b111111111;
assign micromat[95][52] = 9'b111111111;
assign micromat[95][53] = 9'b111111111;
assign micromat[95][54] = 9'b111111111;
assign micromat[95][55] = 9'b111111111;
assign micromat[95][56] = 9'b111111111;
assign micromat[95][57] = 9'b111111111;
assign micromat[95][58] = 9'b111111111;
assign micromat[95][59] = 9'b111111111;
assign micromat[95][60] = 9'b111111111;
assign micromat[95][61] = 9'b111111111;
assign micromat[95][62] = 9'b111111111;
assign micromat[95][63] = 9'b111111111;
assign micromat[95][64] = 9'b111111111;
assign micromat[95][65] = 9'b111111111;
assign micromat[95][66] = 9'b111111111;
assign micromat[95][67] = 9'b111111111;
assign micromat[95][68] = 9'b111111111;
assign micromat[95][69] = 9'b111111111;
assign micromat[95][70] = 9'b111111111;
assign micromat[95][71] = 9'b111111111;
assign micromat[95][72] = 9'b111111111;
assign micromat[95][73] = 9'b111111111;
assign micromat[95][74] = 9'b111111111;
assign micromat[95][75] = 9'b111111111;
assign micromat[95][76] = 9'b111111111;
assign micromat[95][77] = 9'b111111111;
assign micromat[95][78] = 9'b111111111;
assign micromat[95][79] = 9'b111111111;
assign micromat[95][80] = 9'b111111111;
assign micromat[95][81] = 9'b111111111;
assign micromat[95][82] = 9'b111111111;
assign micromat[95][83] = 9'b111111111;
assign micromat[95][84] = 9'b111111111;
assign micromat[95][85] = 9'b111111111;
assign micromat[95][86] = 9'b111111111;
assign micromat[95][87] = 9'b111111111;
assign micromat[95][88] = 9'b111111111;
assign micromat[95][89] = 9'b111111111;
assign micromat[95][90] = 9'b111111111;
assign micromat[95][91] = 9'b111111111;
assign micromat[95][92] = 9'b111111111;
assign micromat[95][93] = 9'b111111111;
assign micromat[95][94] = 9'b111111111;
assign micromat[95][95] = 9'b111111111;
assign micromat[95][96] = 9'b111111111;
assign micromat[95][97] = 9'b111111111;
assign micromat[95][98] = 9'b111111111;
assign micromat[95][99] = 9'b111111111;
assign micromat[96][0] = 9'b111111111;
assign micromat[96][1] = 9'b111111111;
assign micromat[96][2] = 9'b111111111;
assign micromat[96][3] = 9'b111111111;
assign micromat[96][4] = 9'b111111111;
assign micromat[96][5] = 9'b111111111;
assign micromat[96][6] = 9'b111111111;
assign micromat[96][7] = 9'b111111111;
assign micromat[96][8] = 9'b111111111;
assign micromat[96][9] = 9'b111111111;
assign micromat[96][10] = 9'b111111111;
assign micromat[96][11] = 9'b111111111;
assign micromat[96][12] = 9'b111111111;
assign micromat[96][13] = 9'b111111111;
assign micromat[96][14] = 9'b111111111;
assign micromat[96][15] = 9'b111111111;
assign micromat[96][16] = 9'b111111111;
assign micromat[96][17] = 9'b111111111;
assign micromat[96][18] = 9'b111111111;
assign micromat[96][19] = 9'b111111111;
assign micromat[96][20] = 9'b111111111;
assign micromat[96][21] = 9'b111111111;
assign micromat[96][22] = 9'b111111111;
assign micromat[96][23] = 9'b111111111;
assign micromat[96][24] = 9'b111111111;
assign micromat[96][25] = 9'b111111111;
assign micromat[96][26] = 9'b111111111;
assign micromat[96][27] = 9'b111111111;
assign micromat[96][28] = 9'b111111111;
assign micromat[96][29] = 9'b111111111;
assign micromat[96][30] = 9'b111111111;
assign micromat[96][31] = 9'b111111111;
assign micromat[96][32] = 9'b111111111;
assign micromat[96][33] = 9'b111111111;
assign micromat[96][34] = 9'b111111111;
assign micromat[96][35] = 9'b111111111;
assign micromat[96][36] = 9'b111111111;
assign micromat[96][37] = 9'b111111111;
assign micromat[96][38] = 9'b111111111;
assign micromat[96][39] = 9'b111111111;
assign micromat[96][40] = 9'b111111111;
assign micromat[96][41] = 9'b111111111;
assign micromat[96][42] = 9'b111111111;
assign micromat[96][43] = 9'b111111111;
assign micromat[96][44] = 9'b111111111;
assign micromat[96][45] = 9'b111111111;
assign micromat[96][46] = 9'b111111111;
assign micromat[96][47] = 9'b111111111;
assign micromat[96][48] = 9'b111111111;
assign micromat[96][49] = 9'b111111111;
assign micromat[96][50] = 9'b111111111;
assign micromat[96][51] = 9'b111111111;
assign micromat[96][52] = 9'b111111111;
assign micromat[96][53] = 9'b111111111;
assign micromat[96][54] = 9'b111111111;
assign micromat[96][55] = 9'b111111111;
assign micromat[96][56] = 9'b111111111;
assign micromat[96][57] = 9'b111111111;
assign micromat[96][58] = 9'b111111111;
assign micromat[96][59] = 9'b111111111;
assign micromat[96][60] = 9'b111111111;
assign micromat[96][61] = 9'b111111111;
assign micromat[96][62] = 9'b111111111;
assign micromat[96][63] = 9'b111111111;
assign micromat[96][64] = 9'b111111111;
assign micromat[96][65] = 9'b111111111;
assign micromat[96][66] = 9'b111111111;
assign micromat[96][67] = 9'b111111111;
assign micromat[96][68] = 9'b111111111;
assign micromat[96][69] = 9'b111111111;
assign micromat[96][70] = 9'b111111111;
assign micromat[96][71] = 9'b111111111;
assign micromat[96][72] = 9'b111111111;
assign micromat[96][73] = 9'b111111111;
assign micromat[96][74] = 9'b111111111;
assign micromat[96][75] = 9'b111111111;
assign micromat[96][76] = 9'b111111111;
assign micromat[96][77] = 9'b111111111;
assign micromat[96][78] = 9'b111111111;
assign micromat[96][79] = 9'b111111111;
assign micromat[96][80] = 9'b111111111;
assign micromat[96][81] = 9'b111111111;
assign micromat[96][82] = 9'b111111111;
assign micromat[96][83] = 9'b111111111;
assign micromat[96][84] = 9'b111111111;
assign micromat[96][85] = 9'b111111111;
assign micromat[96][86] = 9'b111111111;
assign micromat[96][87] = 9'b111111111;
assign micromat[96][88] = 9'b111111111;
assign micromat[96][89] = 9'b111111111;
assign micromat[96][90] = 9'b111111111;
assign micromat[96][91] = 9'b111111111;
assign micromat[96][92] = 9'b111111111;
assign micromat[96][93] = 9'b111111111;
assign micromat[96][94] = 9'b111111111;
assign micromat[96][95] = 9'b111111111;
assign micromat[96][96] = 9'b111111111;
assign micromat[96][97] = 9'b111111111;
assign micromat[96][98] = 9'b111111111;
assign micromat[96][99] = 9'b111111111;
assign micromat[97][0] = 9'b111111111;
assign micromat[97][1] = 9'b111111111;
assign micromat[97][2] = 9'b111111111;
assign micromat[97][3] = 9'b111111111;
assign micromat[97][4] = 9'b111111111;
assign micromat[97][5] = 9'b111111111;
assign micromat[97][6] = 9'b111111111;
assign micromat[97][7] = 9'b111111111;
assign micromat[97][8] = 9'b111111111;
assign micromat[97][9] = 9'b111111111;
assign micromat[97][10] = 9'b111111111;
assign micromat[97][11] = 9'b111111111;
assign micromat[97][12] = 9'b111111111;
assign micromat[97][13] = 9'b111111111;
assign micromat[97][14] = 9'b111111111;
assign micromat[97][15] = 9'b111111111;
assign micromat[97][16] = 9'b111111111;
assign micromat[97][17] = 9'b111111111;
assign micromat[97][18] = 9'b111111111;
assign micromat[97][19] = 9'b111111111;
assign micromat[97][20] = 9'b111111111;
assign micromat[97][21] = 9'b111111111;
assign micromat[97][22] = 9'b111111111;
assign micromat[97][23] = 9'b111111111;
assign micromat[97][24] = 9'b111111111;
assign micromat[97][25] = 9'b111111111;
assign micromat[97][26] = 9'b111111111;
assign micromat[97][27] = 9'b111111111;
assign micromat[97][28] = 9'b111111111;
assign micromat[97][29] = 9'b111111111;
assign micromat[97][30] = 9'b111111111;
assign micromat[97][31] = 9'b111111111;
assign micromat[97][32] = 9'b111111111;
assign micromat[97][33] = 9'b111111111;
assign micromat[97][34] = 9'b111111111;
assign micromat[97][35] = 9'b111111111;
assign micromat[97][36] = 9'b111111111;
assign micromat[97][37] = 9'b111111111;
assign micromat[97][38] = 9'b111111111;
assign micromat[97][39] = 9'b111111111;
assign micromat[97][40] = 9'b111111111;
assign micromat[97][41] = 9'b111111111;
assign micromat[97][42] = 9'b111111111;
assign micromat[97][43] = 9'b111111111;
assign micromat[97][44] = 9'b111111111;
assign micromat[97][45] = 9'b111111111;
assign micromat[97][46] = 9'b111111111;
assign micromat[97][47] = 9'b111111111;
assign micromat[97][48] = 9'b111111111;
assign micromat[97][49] = 9'b111111111;
assign micromat[97][50] = 9'b111111111;
assign micromat[97][51] = 9'b111111111;
assign micromat[97][52] = 9'b111111111;
assign micromat[97][53] = 9'b111111111;
assign micromat[97][54] = 9'b111111111;
assign micromat[97][55] = 9'b111111111;
assign micromat[97][56] = 9'b111111111;
assign micromat[97][57] = 9'b111111111;
assign micromat[97][58] = 9'b111111111;
assign micromat[97][59] = 9'b111111111;
assign micromat[97][60] = 9'b111111111;
assign micromat[97][61] = 9'b111111111;
assign micromat[97][62] = 9'b111111111;
assign micromat[97][63] = 9'b111111111;
assign micromat[97][64] = 9'b111111111;
assign micromat[97][65] = 9'b111111111;
assign micromat[97][66] = 9'b111111111;
assign micromat[97][67] = 9'b111111111;
assign micromat[97][68] = 9'b111111111;
assign micromat[97][69] = 9'b111111111;
assign micromat[97][70] = 9'b111111111;
assign micromat[97][71] = 9'b111111111;
assign micromat[97][72] = 9'b111111111;
assign micromat[97][73] = 9'b111111111;
assign micromat[97][74] = 9'b111111111;
assign micromat[97][75] = 9'b111111111;
assign micromat[97][76] = 9'b111111111;
assign micromat[97][77] = 9'b111111111;
assign micromat[97][78] = 9'b111111111;
assign micromat[97][79] = 9'b111111111;
assign micromat[97][80] = 9'b111111111;
assign micromat[97][81] = 9'b111111111;
assign micromat[97][82] = 9'b111111111;
assign micromat[97][83] = 9'b111111111;
assign micromat[97][84] = 9'b111111111;
assign micromat[97][85] = 9'b111111111;
assign micromat[97][86] = 9'b111111111;
assign micromat[97][87] = 9'b111111111;
assign micromat[97][88] = 9'b111111111;
assign micromat[97][89] = 9'b111111111;
assign micromat[97][90] = 9'b111111111;
assign micromat[97][91] = 9'b111111111;
assign micromat[97][92] = 9'b111111111;
assign micromat[97][93] = 9'b111111111;
assign micromat[97][94] = 9'b111111111;
assign micromat[97][95] = 9'b111111111;
assign micromat[97][96] = 9'b111111111;
assign micromat[97][97] = 9'b111111111;
assign micromat[97][98] = 9'b111111111;
assign micromat[97][99] = 9'b111111111;
assign micromat[98][0] = 9'b111111111;
assign micromat[98][1] = 9'b111111111;
assign micromat[98][2] = 9'b111111111;
assign micromat[98][3] = 9'b111111111;
assign micromat[98][4] = 9'b111111111;
assign micromat[98][5] = 9'b111111111;
assign micromat[98][6] = 9'b111111111;
assign micromat[98][7] = 9'b111111111;
assign micromat[98][8] = 9'b111111111;
assign micromat[98][9] = 9'b111111111;
assign micromat[98][10] = 9'b111111111;
assign micromat[98][11] = 9'b111111111;
assign micromat[98][12] = 9'b111111111;
assign micromat[98][13] = 9'b111111111;
assign micromat[98][14] = 9'b111111111;
assign micromat[98][15] = 9'b111111111;
assign micromat[98][16] = 9'b111111111;
assign micromat[98][17] = 9'b111111111;
assign micromat[98][18] = 9'b111111111;
assign micromat[98][19] = 9'b111111111;
assign micromat[98][20] = 9'b111111111;
assign micromat[98][21] = 9'b111111111;
assign micromat[98][22] = 9'b111111111;
assign micromat[98][23] = 9'b111111111;
assign micromat[98][24] = 9'b111111111;
assign micromat[98][25] = 9'b111111111;
assign micromat[98][26] = 9'b111111111;
assign micromat[98][27] = 9'b111111111;
assign micromat[98][28] = 9'b111111111;
assign micromat[98][29] = 9'b111111111;
assign micromat[98][30] = 9'b111111111;
assign micromat[98][31] = 9'b111111111;
assign micromat[98][32] = 9'b111111111;
assign micromat[98][33] = 9'b111111111;
assign micromat[98][34] = 9'b111111111;
assign micromat[98][35] = 9'b111111111;
assign micromat[98][36] = 9'b111111111;
assign micromat[98][37] = 9'b111111111;
assign micromat[98][38] = 9'b111111111;
assign micromat[98][39] = 9'b111111111;
assign micromat[98][40] = 9'b111111111;
assign micromat[98][41] = 9'b111111111;
assign micromat[98][42] = 9'b111111111;
assign micromat[98][43] = 9'b111111111;
assign micromat[98][44] = 9'b111111111;
assign micromat[98][45] = 9'b111111111;
assign micromat[98][46] = 9'b111111111;
assign micromat[98][47] = 9'b111111111;
assign micromat[98][48] = 9'b111111111;
assign micromat[98][49] = 9'b111111111;
assign micromat[98][50] = 9'b111111111;
assign micromat[98][51] = 9'b111111111;
assign micromat[98][52] = 9'b111111111;
assign micromat[98][53] = 9'b111111111;
assign micromat[98][54] = 9'b111111111;
assign micromat[98][55] = 9'b111111111;
assign micromat[98][56] = 9'b111111111;
assign micromat[98][57] = 9'b111111111;
assign micromat[98][58] = 9'b111111111;
assign micromat[98][59] = 9'b111111111;
assign micromat[98][60] = 9'b111111111;
assign micromat[98][61] = 9'b111111111;
assign micromat[98][62] = 9'b111111111;
assign micromat[98][63] = 9'b111111111;
assign micromat[98][64] = 9'b111111111;
assign micromat[98][65] = 9'b111111111;
assign micromat[98][66] = 9'b111111111;
assign micromat[98][67] = 9'b111111111;
assign micromat[98][68] = 9'b111111111;
assign micromat[98][69] = 9'b111111111;
assign micromat[98][70] = 9'b111111111;
assign micromat[98][71] = 9'b111111111;
assign micromat[98][72] = 9'b111111111;
assign micromat[98][73] = 9'b111111111;
assign micromat[98][74] = 9'b111111111;
assign micromat[98][75] = 9'b111111111;
assign micromat[98][76] = 9'b111111111;
assign micromat[98][77] = 9'b111111111;
assign micromat[98][78] = 9'b111111111;
assign micromat[98][79] = 9'b111111111;
assign micromat[98][80] = 9'b111111111;
assign micromat[98][81] = 9'b111111111;
assign micromat[98][82] = 9'b111111111;
assign micromat[98][83] = 9'b111111111;
assign micromat[98][84] = 9'b111111111;
assign micromat[98][85] = 9'b111111111;
assign micromat[98][86] = 9'b111111111;
assign micromat[98][87] = 9'b111111111;
assign micromat[98][88] = 9'b111111111;
assign micromat[98][89] = 9'b111111111;
assign micromat[98][90] = 9'b111111111;
assign micromat[98][91] = 9'b111111111;
assign micromat[98][92] = 9'b111111111;
assign micromat[98][93] = 9'b111111111;
assign micromat[98][94] = 9'b111111111;
assign micromat[98][95] = 9'b111111111;
assign micromat[98][96] = 9'b111111111;
assign micromat[98][97] = 9'b111111111;
assign micromat[98][98] = 9'b111111111;
assign micromat[98][99] = 9'b111111111;
assign micromat[99][0] = 9'b111111111;
assign micromat[99][1] = 9'b111111111;
assign micromat[99][2] = 9'b111111111;
assign micromat[99][3] = 9'b111111111;
assign micromat[99][4] = 9'b111111111;
assign micromat[99][5] = 9'b111111111;
assign micromat[99][6] = 9'b111111111;
assign micromat[99][7] = 9'b111111111;
assign micromat[99][8] = 9'b111111111;
assign micromat[99][9] = 9'b111111111;
assign micromat[99][10] = 9'b111111111;
assign micromat[99][11] = 9'b111111111;
assign micromat[99][12] = 9'b111111111;
assign micromat[99][13] = 9'b111111111;
assign micromat[99][14] = 9'b111111111;
assign micromat[99][15] = 9'b111111111;
assign micromat[99][16] = 9'b111111111;
assign micromat[99][17] = 9'b111111111;
assign micromat[99][18] = 9'b111111111;
assign micromat[99][19] = 9'b111111111;
assign micromat[99][20] = 9'b111111111;
assign micromat[99][21] = 9'b111111111;
assign micromat[99][22] = 9'b111111111;
assign micromat[99][23] = 9'b111111111;
assign micromat[99][24] = 9'b111111111;
assign micromat[99][25] = 9'b111111111;
assign micromat[99][26] = 9'b111111111;
assign micromat[99][27] = 9'b111111111;
assign micromat[99][28] = 9'b111111111;
assign micromat[99][29] = 9'b111111111;
assign micromat[99][30] = 9'b111111111;
assign micromat[99][31] = 9'b111111111;
assign micromat[99][32] = 9'b111111111;
assign micromat[99][33] = 9'b111111111;
assign micromat[99][34] = 9'b111111111;
assign micromat[99][35] = 9'b111111111;
assign micromat[99][36] = 9'b111111111;
assign micromat[99][37] = 9'b111111111;
assign micromat[99][38] = 9'b111111111;
assign micromat[99][39] = 9'b111111111;
assign micromat[99][40] = 9'b111111111;
assign micromat[99][41] = 9'b111111111;
assign micromat[99][42] = 9'b111111111;
assign micromat[99][43] = 9'b111111111;
assign micromat[99][44] = 9'b111111111;
assign micromat[99][45] = 9'b111111111;
assign micromat[99][46] = 9'b111111111;
assign micromat[99][47] = 9'b111111111;
assign micromat[99][48] = 9'b111111111;
assign micromat[99][49] = 9'b111111111;
assign micromat[99][50] = 9'b111111111;
assign micromat[99][51] = 9'b111111111;
assign micromat[99][52] = 9'b111111111;
assign micromat[99][53] = 9'b111111111;
assign micromat[99][54] = 9'b111111111;
assign micromat[99][55] = 9'b111111111;
assign micromat[99][56] = 9'b111111111;
assign micromat[99][57] = 9'b111111111;
assign micromat[99][58] = 9'b111111111;
assign micromat[99][59] = 9'b111111111;
assign micromat[99][60] = 9'b111111111;
assign micromat[99][61] = 9'b111111111;
assign micromat[99][62] = 9'b111111111;
assign micromat[99][63] = 9'b111111111;
assign micromat[99][64] = 9'b111111111;
assign micromat[99][65] = 9'b111111111;
assign micromat[99][66] = 9'b111111111;
assign micromat[99][67] = 9'b111111111;
assign micromat[99][68] = 9'b111111111;
assign micromat[99][69] = 9'b111111111;
assign micromat[99][70] = 9'b111111111;
assign micromat[99][71] = 9'b111111111;
assign micromat[99][72] = 9'b111111111;
assign micromat[99][73] = 9'b111111111;
assign micromat[99][74] = 9'b111111111;
assign micromat[99][75] = 9'b111111111;
assign micromat[99][76] = 9'b111111111;
assign micromat[99][77] = 9'b111111111;
assign micromat[99][78] = 9'b111111111;
assign micromat[99][79] = 9'b111111111;
assign micromat[99][80] = 9'b111111111;
assign micromat[99][81] = 9'b111111111;
assign micromat[99][82] = 9'b111111111;
assign micromat[99][83] = 9'b111111111;
assign micromat[99][84] = 9'b111111111;
assign micromat[99][85] = 9'b111111111;
assign micromat[99][86] = 9'b111111111;
assign micromat[99][87] = 9'b111111111;
assign micromat[99][88] = 9'b111111111;
assign micromat[99][89] = 9'b111111111;
assign micromat[99][90] = 9'b111111111;
assign micromat[99][91] = 9'b111111111;
assign micromat[99][92] = 9'b111111111;
assign micromat[99][93] = 9'b111111111;
assign micromat[99][94] = 9'b111111111;
assign micromat[99][95] = 9'b111111111;
assign micromat[99][96] = 9'b111111111;
assign micromat[99][97] = 9'b111111111;
assign micromat[99][98] = 9'b111111111;
assign micromat[99][99] = 9'b111111111;
//Total de Lineas = 10000
endmodule



