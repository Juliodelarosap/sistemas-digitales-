`timescale 1ns / 1ps
module gameover (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (f[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= f[vcount- posy][hcount- posx][7:5];
				green <= f[vcount- posy][hcount- posx][4:2];
            blue 	<= f[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 32;
parameter RESOLUCION_Y = 32;
wire [8:0] f[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign f[0][14] = 9'b101101101;
assign f[0][15] = 9'b101001001;
assign f[0][16] = 9'b101001000;
assign f[0][17] = 9'b100100100;
assign f[1][12] = 9'b101101101;
assign f[1][13] = 9'b101101101;
assign f[1][14] = 9'b101001001;
assign f[1][15] = 9'b101001000;
assign f[1][16] = 9'b100100100;
assign f[1][17] = 9'b100100100;
assign f[1][18] = 9'b100100100;
assign f[1][19] = 9'b100100100;
assign f[2][11] = 9'b110010001;
assign f[2][12] = 9'b101101101;
assign f[2][13] = 9'b101101101;
assign f[2][14] = 9'b101001001;
assign f[2][15] = 9'b101001000;
assign f[2][16] = 9'b100100100;
assign f[2][17] = 9'b100100100;
assign f[2][18] = 9'b100100100;
assign f[2][19] = 9'b100000000;
assign f[2][20] = 9'b100100100;
assign f[3][11] = 9'b110010001;
assign f[3][12] = 9'b101101101;
assign f[3][13] = 9'b101001001;
assign f[3][14] = 9'b101001001;
assign f[3][15] = 9'b100100100;
assign f[3][16] = 9'b100100100;
assign f[3][17] = 9'b100100100;
assign f[3][18] = 9'b100000000;
assign f[3][19] = 9'b100000000;
assign f[3][20] = 9'b100000000;
assign f[4][10] = 9'b110010001;
assign f[4][11] = 9'b110010001;
assign f[4][12] = 9'b111111101;
assign f[4][13] = 9'b101101101;
assign f[4][14] = 9'b110010001;
assign f[4][15] = 9'b101101100;
assign f[4][16] = 9'b101001000;
assign f[4][17] = 9'b101001000;
assign f[4][18] = 9'b101101100;
assign f[4][19] = 9'b110010000;
assign f[4][20] = 9'b101101100;
assign f[4][21] = 9'b100000000;
assign f[5][10] = 9'b110010001;
assign f[5][11] = 9'b110110101;
assign f[5][12] = 9'b110110101;
assign f[5][13] = 9'b101101101;
assign f[5][14] = 9'b111111101;
assign f[5][15] = 9'b110010000;
assign f[5][16] = 9'b110110100;
assign f[5][17] = 9'b110110100;
assign f[5][18] = 9'b111111100;
assign f[5][19] = 9'b101101100;
assign f[5][20] = 9'b100100100;
assign f[5][21] = 9'b100000000;
assign f[6][9] = 9'b110010010;
assign f[6][10] = 9'b110010010;
assign f[6][11] = 9'b111111101;
assign f[6][12] = 9'b101101101;
assign f[6][13] = 9'b110010001;
assign f[6][14] = 9'b101101101;
assign f[6][15] = 9'b110010000;
assign f[6][16] = 9'b111111100;
assign f[6][17] = 9'b111111100;
assign f[6][18] = 9'b111111100;
assign f[6][19] = 9'b101001000;
assign f[6][20] = 9'b100000000;
assign f[6][21] = 9'b100000000;
assign f[6][22] = 9'b100000000;
assign f[7][9] = 9'b110010010;
assign f[7][10] = 9'b110010001;
assign f[7][11] = 9'b110110101;
assign f[7][12] = 9'b110110101;
assign f[7][13] = 9'b111111101;
assign f[7][14] = 9'b110010001;
assign f[7][15] = 9'b110110100;
assign f[7][16] = 9'b111111100;
assign f[7][17] = 9'b111111100;
assign f[7][18] = 9'b111111100;
assign f[7][19] = 9'b111111100;
assign f[7][20] = 9'b100100100;
assign f[7][21] = 9'b100000000;
assign f[7][22] = 9'b100000000;
assign f[8][9] = 9'b110010001;
assign f[8][10] = 9'b110010001;
assign f[8][11] = 9'b110110101;
assign f[8][12] = 9'b110010001;
assign f[8][13] = 9'b111111101;
assign f[8][14] = 9'b111111101;
assign f[8][15] = 9'b111111100;
assign f[8][16] = 9'b110010000;
assign f[8][17] = 9'b101101100;
assign f[8][18] = 9'b111111100;
assign f[8][19] = 9'b100100100;
assign f[8][20] = 9'b100000000;
assign f[8][21] = 9'b100000000;
assign f[8][22] = 9'b100000000;
assign f[9][9] = 9'b110010001;
assign f[9][10] = 9'b101101101;
assign f[9][11] = 9'b110010001;
assign f[9][12] = 9'b111111101;
assign f[9][13] = 9'b111111101;
assign f[9][14] = 9'b101101101;
assign f[9][15] = 9'b110110100;
assign f[9][16] = 9'b110010000;
assign f[9][17] = 9'b101001000;
assign f[9][18] = 9'b111111100;
assign f[9][19] = 9'b110010000;
assign f[9][20] = 9'b101101000;
assign f[9][21] = 9'b100000000;
assign f[9][22] = 9'b100000000;
assign f[10][9] = 9'b110010001;
assign f[10][10] = 9'b101101101;
assign f[10][11] = 9'b110010001;
assign f[10][12] = 9'b111111101;
assign f[10][13] = 9'b110010001;
assign f[10][14] = 9'b101001000;
assign f[10][15] = 9'b101101100;
assign f[10][16] = 9'b101101100;
assign f[10][17] = 9'b101101000;
assign f[10][18] = 9'b101101100;
assign f[10][19] = 9'b110010000;
assign f[10][20] = 9'b101101000;
assign f[10][21] = 9'b100000000;
assign f[10][22] = 9'b100000000;
assign f[11][9] = 9'b110010001;
assign f[11][10] = 9'b101101101;
assign f[11][11] = 9'b110110101;
assign f[11][12] = 9'b111111101;
assign f[11][13] = 9'b110010001;
assign f[11][14] = 9'b101101100;
assign f[11][15] = 9'b110001100;
assign f[11][16] = 9'b111110000;
assign f[11][17] = 9'b110110000;
assign f[11][18] = 9'b110001100;
assign f[11][19] = 9'b111101100;
assign f[11][20] = 9'b101101000;
assign f[11][21] = 9'b100000000;
assign f[11][22] = 9'b100000000;
assign f[12][9] = 9'b110010001;
assign f[12][10] = 9'b110010001;
assign f[12][11] = 9'b110110001;
assign f[12][12] = 9'b110001101;
assign f[12][13] = 9'b111110001;
assign f[12][14] = 9'b101101000;
assign f[12][15] = 9'b110001100;
assign f[12][16] = 9'b110101100;
assign f[12][17] = 9'b100000000;
assign f[12][18] = 9'b101101000;
assign f[12][19] = 9'b101000100;
assign f[12][20] = 9'b110001000;
assign f[12][21] = 9'b100000000;
assign f[12][22] = 9'b100000000;
assign f[13][9] = 9'b110001101;
assign f[13][10] = 9'b101101101;
assign f[13][11] = 9'b110110001;
assign f[13][12] = 9'b101101101;
assign f[13][13] = 9'b111101101;
assign f[13][14] = 9'b110001000;
assign f[13][15] = 9'b110101000;
assign f[13][16] = 9'b111101000;
assign f[13][17] = 9'b101100100;
assign f[13][18] = 9'b101100100;
assign f[13][19] = 9'b101100100;
assign f[13][20] = 9'b110000100;
assign f[13][21] = 9'b100000000;
assign f[13][22] = 9'b100000000;
assign f[14][8] = 9'b111100000;
assign f[14][9] = 9'b110001001;
assign f[14][10] = 9'b101101101;
assign f[14][11] = 9'b110101101;
assign f[14][12] = 9'b101101001;
assign f[14][13] = 9'b111101000;
assign f[14][14] = 9'b111101000;
assign f[14][15] = 9'b111100100;
assign f[14][16] = 9'b111100100;
assign f[14][17] = 9'b101100100;
assign f[14][18] = 9'b101100000;
assign f[14][19] = 9'b111100000;
assign f[14][20] = 9'b101100000;
assign f[14][21] = 9'b100000000;
assign f[14][22] = 9'b100100000;
assign f[14][23] = 9'b101100000;
assign f[15][8] = 9'b111100000;
assign f[15][9] = 9'b101100100;
assign f[15][10] = 9'b101101101;
assign f[15][11] = 9'b110001001;
assign f[15][12] = 9'b101101001;
assign f[15][13] = 9'b110001000;
assign f[15][14] = 9'b111100100;
assign f[15][15] = 9'b110000100;
assign f[15][16] = 9'b110000100;
assign f[15][17] = 9'b100000100;
assign f[15][18] = 9'b101000000;
assign f[15][19] = 9'b111100000;
assign f[15][20] = 9'b101100000;
assign f[15][21] = 9'b100000000;
assign f[15][22] = 9'b100100000;
assign f[15][23] = 9'b101100000;
assign f[16][8] = 9'b111100000;
assign f[16][9] = 9'b101100000;
assign f[16][10] = 9'b101001101;
assign f[16][11] = 9'b111101001;
assign f[16][12] = 9'b111101001;
assign f[16][13] = 9'b101000100;
assign f[16][14] = 9'b110000100;
assign f[16][15] = 9'b101000100;
assign f[16][16] = 9'b111100100;
assign f[16][17] = 9'b110100100;
assign f[16][18] = 9'b110100000;
assign f[16][19] = 9'b110000000;
assign f[16][20] = 9'b111100000;
assign f[16][21] = 9'b100000000;
assign f[16][22] = 9'b101000000;
assign f[16][23] = 9'b101100000;
assign f[17][8] = 9'b111100000;
assign f[17][9] = 9'b101000000;
assign f[17][10] = 9'b100101000;
assign f[17][11] = 9'b101101001;
assign f[17][12] = 9'b101101000;
assign f[17][13] = 9'b100100100;
assign f[17][14] = 9'b100100100;
assign f[17][15] = 9'b100100100;
assign f[17][16] = 9'b101000100;
assign f[17][17] = 9'b101100000;
assign f[17][18] = 9'b101000000;
assign f[17][19] = 9'b100100000;
assign f[17][20] = 9'b101000000;
assign f[17][21] = 9'b100000000;
assign f[17][22] = 9'b101000000;
assign f[17][23] = 9'b101100000;
assign f[18][8] = 9'b111100000;
assign f[18][9] = 9'b101000000;
assign f[18][10] = 9'b100000000;
assign f[18][11] = 9'b101001001;
assign f[18][12] = 9'b100101000;
assign f[18][13] = 9'b100100100;
assign f[18][14] = 9'b100100100;
assign f[18][15] = 9'b100100100;
assign f[18][16] = 9'b100000100;
assign f[18][17] = 9'b100000000;
assign f[18][18] = 9'b100000000;
assign f[18][19] = 9'b100000000;
assign f[18][20] = 9'b100000000;
assign f[18][21] = 9'b100000000;
assign f[18][22] = 9'b101100000;
assign f[18][23] = 9'b101100000;
assign f[19][8] = 9'b111100100;
assign f[19][9] = 9'b101100000;
assign f[19][10] = 9'b100000000;
assign f[19][11] = 9'b100100100;
assign f[19][12] = 9'b101001000;
assign f[19][13] = 9'b100100100;
assign f[19][14] = 9'b100100100;
assign f[19][15] = 9'b100100100;
assign f[19][16] = 9'b100100100;
assign f[19][17] = 9'b100000000;
assign f[19][18] = 9'b100000000;
assign f[19][19] = 9'b100000000;
assign f[19][20] = 9'b100000000;
assign f[19][21] = 9'b100000000;
assign f[19][22] = 9'b101100000;
assign f[19][23] = 9'b101000000;
assign f[20][8] = 9'b111100100;
assign f[20][9] = 9'b110000000;
assign f[20][10] = 9'b100000000;
assign f[20][11] = 9'b100000000;
assign f[20][12] = 9'b100100100;
assign f[20][13] = 9'b100100100;
assign f[20][14] = 9'b100100100;
assign f[20][15] = 9'b100100100;
assign f[20][16] = 9'b100000000;
assign f[20][17] = 9'b100000000;
assign f[20][18] = 9'b100000000;
assign f[20][19] = 9'b100000000;
assign f[20][20] = 9'b100000000;
assign f[20][21] = 9'b100000000;
assign f[20][22] = 9'b101100000;
assign f[20][23] = 9'b101000000;
assign f[21][8] = 9'b111100100;
assign f[21][9] = 9'b110100000;
assign f[21][10] = 9'b100000000;
assign f[21][11] = 9'b100000000;
assign f[21][12] = 9'b100000000;
assign f[21][13] = 9'b101001001;
assign f[21][14] = 9'b100100100;
assign f[21][15] = 9'b100100100;
assign f[21][16] = 9'b100000000;
assign f[21][17] = 9'b100000000;
assign f[21][18] = 9'b100000000;
assign f[21][19] = 9'b100000000;
assign f[21][20] = 9'b100000000;
assign f[21][21] = 9'b100000000;
assign f[21][22] = 9'b101100000;
assign f[21][23] = 9'b100100000;
assign f[22][8] = 9'b111100100;
assign f[22][9] = 9'b111100000;
assign f[22][10] = 9'b100100000;
assign f[22][11] = 9'b100000000;
assign f[22][12] = 9'b100000000;
assign f[22][13] = 9'b101101101;
assign f[22][14] = 9'b110010001;
assign f[22][15] = 9'b101001001;
assign f[22][16] = 9'b100000000;
assign f[22][17] = 9'b100000000;
assign f[22][18] = 9'b100000000;
assign f[22][19] = 9'b100000000;
assign f[22][20] = 9'b100000000;
assign f[22][21] = 9'b100100000;
assign f[22][22] = 9'b101100000;
assign f[22][23] = 9'b100000000;
assign f[23][8] = 9'b111100100;
assign f[23][9] = 9'b111100100;
assign f[23][10] = 9'b101000000;
assign f[23][11] = 9'b100000000;
assign f[23][12] = 9'b100000000;
assign f[23][13] = 9'b101101101;
assign f[23][14] = 9'b110010001;
assign f[23][15] = 9'b101001001;
assign f[23][16] = 9'b100000000;
assign f[23][17] = 9'b100000000;
assign f[23][18] = 9'b100000000;
assign f[23][19] = 9'b100000000;
assign f[23][20] = 9'b100000000;
assign f[23][21] = 9'b101100000;
assign f[23][22] = 9'b101000000;
assign f[23][23] = 9'b100000000;
assign f[24][8] = 9'b111100000;
assign f[24][9] = 9'b111100100;
assign f[24][10] = 9'b110100000;
assign f[24][11] = 9'b100000000;
assign f[24][12] = 9'b100000000;
assign f[24][13] = 9'b101001001;
assign f[24][14] = 9'b110010001;
assign f[24][15] = 9'b101001001;
assign f[24][16] = 9'b100000000;
assign f[24][17] = 9'b100000000;
assign f[24][18] = 9'b100000000;
assign f[24][19] = 9'b100000000;
assign f[24][20] = 9'b100000000;
assign f[24][21] = 9'b101100000;
assign f[24][22] = 9'b100100000;
assign f[24][23] = 9'b100000000;
assign f[25][9] = 9'b111100100;
assign f[25][10] = 9'b111100000;
assign f[25][11] = 9'b101100000;
assign f[25][12] = 9'b100000000;
assign f[25][13] = 9'b101001001;
assign f[25][14] = 9'b110001101;
assign f[25][15] = 9'b101001001;
assign f[25][16] = 9'b100000000;
assign f[25][17] = 9'b100000000;
assign f[25][18] = 9'b100000000;
assign f[25][19] = 9'b100000000;
assign f[25][20] = 9'b101100000;
assign f[25][21] = 9'b101000000;
assign f[25][22] = 9'b100000000;
assign f[26][9] = 9'b111100000;
assign f[26][10] = 9'b111101000;
assign f[26][11] = 9'b111100000;
assign f[26][12] = 9'b101000000;
assign f[26][13] = 9'b101001001;
assign f[26][14] = 9'b101101101;
assign f[26][15] = 9'b101001000;
assign f[26][16] = 9'b100000000;
assign f[26][17] = 9'b100000000;
assign f[26][18] = 9'b100000000;
assign f[26][19] = 9'b101000000;
assign f[26][20] = 9'b101100000;
assign f[26][21] = 9'b100100000;
assign f[26][22] = 9'b100000000;
assign f[27][10] = 9'b111100100;
assign f[27][11] = 9'b111101001;
assign f[27][12] = 9'b111100000;
assign f[27][13] = 9'b101100000;
assign f[27][14] = 9'b101101001;
assign f[27][15] = 9'b101001000;
assign f[27][16] = 9'b100000000;
assign f[27][17] = 9'b100100000;
assign f[27][18] = 9'b101100000;
assign f[27][19] = 9'b101100000;
assign f[27][20] = 9'b101000000;
assign f[27][21] = 9'b100100000;
assign f[28][10] = 9'b111100000;
assign f[28][11] = 9'b111101000;
assign f[28][12] = 9'b111101000;
assign f[28][13] = 9'b110100000;
assign f[28][14] = 9'b110000000;
assign f[28][15] = 9'b110000000;
assign f[28][16] = 9'b101100000;
assign f[28][17] = 9'b110000000;
assign f[28][18] = 9'b101100000;
assign f[28][19] = 9'b101000000;
assign f[28][20] = 9'b101000000;
assign f[28][21] = 9'b100100000;
assign f[29][11] = 9'b111100000;
assign f[29][12] = 9'b111100100;
assign f[29][13] = 9'b111100100;
assign f[29][14] = 9'b110100000;
assign f[29][15] = 9'b110000000;
assign f[29][16] = 9'b101100000;
assign f[29][17] = 9'b101100000;
assign f[29][18] = 9'b101100000;
assign f[29][19] = 9'b101000000;
assign f[29][20] = 9'b100100000;
assign f[30][12] = 9'b111100000;
assign f[30][13] = 9'b111100000;
assign f[30][14] = 9'b110100000;
assign f[30][15] = 9'b110000000;
assign f[30][16] = 9'b110000000;
assign f[30][17] = 9'b101100000;
assign f[30][18] = 9'b101100000;
assign f[30][19] = 9'b101000000;
assign f[31][14] = 9'b110100000;
assign f[31][15] = 9'b110000000;
assign f[31][16] = 9'b110000000;
assign f[31][17] = 9'b101100000;
//Total de Lineas = 418
endmodule

