`timescale 1ns / 1ps
module logo (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (f[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= f[vcount- posy][hcount- posx][7:5];
				green <= f[vcount- posy][hcount- posx][4:2];
            blue 	<= f[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 200;
parameter RESOLUCION_Y = 100;
wire [8:0] f[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign f[31][20] = 9'b111111111;
assign f[31][21] = 9'b111111111;
assign f[31][22] = 9'b111111111;
assign f[31][23] = 9'b111111111;
assign f[31][24] = 9'b111111111;
assign f[31][25] = 9'b111111111;
assign f[31][26] = 9'b111111111;
assign f[31][27] = 9'b111111111;
assign f[31][28] = 9'b111111111;
assign f[31][29] = 9'b111111111;
assign f[31][30] = 9'b111111111;
assign f[31][32] = 9'b111111111;
assign f[31][33] = 9'b111111111;
assign f[31][34] = 9'b111111111;
assign f[31][35] = 9'b111111111;
assign f[31][38] = 9'b111111111;
assign f[31][39] = 9'b111111111;
assign f[31][42] = 9'b111111111;
assign f[31][43] = 9'b111111111;
assign f[31][44] = 9'b111111111;
assign f[31][45] = 9'b111111111;
assign f[31][46] = 9'b111111111;
assign f[31][47] = 9'b111111111;
assign f[31][56] = 9'b111111111;
assign f[31][57] = 9'b111111111;
assign f[31][58] = 9'b111111111;
assign f[31][59] = 9'b111111111;
assign f[31][60] = 9'b111111111;
assign f[31][61] = 9'b111111111;
assign f[31][62] = 9'b111111111;
assign f[31][66] = 9'b111111111;
assign f[31][67] = 9'b111111111;
assign f[31][68] = 9'b111111111;
assign f[31][69] = 9'b111111111;
assign f[31][70] = 9'b111111111;
assign f[31][71] = 9'b111111111;
assign f[31][72] = 9'b111111111;
assign f[31][73] = 9'b111111111;
assign f[31][74] = 9'b111111111;
assign f[31][75] = 9'b111111111;
assign f[31][76] = 9'b111111111;
assign f[31][77] = 9'b111111111;
assign f[31][78] = 9'b111111111;
assign f[31][79] = 9'b111111111;
assign f[31][80] = 9'b111111111;
assign f[31][81] = 9'b111111111;
assign f[31][94] = 9'b111111111;
assign f[31][95] = 9'b111111111;
assign f[31][96] = 9'b111111111;
assign f[31][97] = 9'b111111111;
assign f[31][98] = 9'b111111111;
assign f[31][99] = 9'b111111111;
assign f[31][100] = 9'b111111111;
assign f[31][101] = 9'b111111111;
assign f[31][102] = 9'b111111111;
assign f[31][103] = 9'b111111111;
assign f[31][104] = 9'b111111111;
assign f[31][105] = 9'b111111111;
assign f[31][106] = 9'b111111111;
assign f[31][107] = 9'b111111111;
assign f[31][117] = 9'b111111111;
assign f[31][118] = 9'b111111111;
assign f[31][119] = 9'b111111111;
assign f[31][120] = 9'b111111111;
assign f[31][121] = 9'b111111111;
assign f[31][122] = 9'b111111111;
assign f[31][123] = 9'b111111111;
assign f[31][146] = 9'b111111111;
assign f[31][147] = 9'b111111111;
assign f[31][148] = 9'b111111111;
assign f[31][149] = 9'b111111111;
assign f[31][150] = 9'b111111111;
assign f[31][151] = 9'b111111111;
assign f[31][152] = 9'b111111111;
assign f[31][153] = 9'b111111111;
assign f[31][164] = 9'b111111111;
assign f[31][165] = 9'b111111111;
assign f[31][166] = 9'b111111111;
assign f[31][167] = 9'b111111111;
assign f[31][168] = 9'b111111111;
assign f[31][169] = 9'b111111111;
assign f[31][170] = 9'b111111111;
assign f[31][171] = 9'b111111111;
assign f[31][172] = 9'b111111111;
assign f[31][180] = 9'b111111111;
assign f[31][181] = 9'b111111111;
assign f[31][182] = 9'b111111111;
assign f[31][183] = 9'b111111111;
assign f[31][184] = 9'b111111111;
assign f[31][185] = 9'b111111111;
assign f[32][19] = 9'b111111111;
assign f[32][20] = 9'b111111111;
assign f[32][21] = 9'b111111111;
assign f[32][22] = 9'b111111111;
assign f[32][23] = 9'b111111111;
assign f[32][24] = 9'b111111111;
assign f[32][25] = 9'b111111111;
assign f[32][26] = 9'b111111111;
assign f[32][27] = 9'b111111111;
assign f[32][28] = 9'b111111111;
assign f[32][29] = 9'b111111111;
assign f[32][30] = 9'b111111111;
assign f[32][31] = 9'b111111111;
assign f[32][32] = 9'b111111111;
assign f[32][33] = 9'b111111111;
assign f[32][34] = 9'b111111111;
assign f[32][35] = 9'b111111111;
assign f[32][36] = 9'b111111111;
assign f[32][37] = 9'b111111111;
assign f[32][38] = 9'b111111111;
assign f[32][39] = 9'b111111111;
assign f[32][40] = 9'b111111111;
assign f[32][42] = 9'b111111111;
assign f[32][43] = 9'b111111111;
assign f[32][44] = 9'b111111111;
assign f[32][45] = 9'b111111111;
assign f[32][46] = 9'b111111111;
assign f[32][47] = 9'b111111111;
assign f[32][48] = 9'b111111111;
assign f[32][56] = 9'b111111111;
assign f[32][57] = 9'b111111111;
assign f[32][58] = 9'b111111111;
assign f[32][59] = 9'b111111111;
assign f[32][60] = 9'b111111111;
assign f[32][61] = 9'b111111111;
assign f[32][62] = 9'b111111111;
assign f[32][65] = 9'b111111111;
assign f[32][66] = 9'b111111111;
assign f[32][67] = 9'b111111111;
assign f[32][68] = 9'b111111111;
assign f[32][69] = 9'b111111111;
assign f[32][70] = 9'b111111111;
assign f[32][71] = 9'b111111111;
assign f[32][72] = 9'b111111111;
assign f[32][73] = 9'b111111111;
assign f[32][74] = 9'b111111111;
assign f[32][75] = 9'b111111111;
assign f[32][76] = 9'b111111111;
assign f[32][77] = 9'b111111111;
assign f[32][78] = 9'b111111111;
assign f[32][79] = 9'b111111111;
assign f[32][80] = 9'b111111111;
assign f[32][81] = 9'b111111111;
assign f[32][94] = 9'b111111111;
assign f[32][95] = 9'b111111111;
assign f[32][96] = 9'b111111111;
assign f[32][97] = 9'b111111111;
assign f[32][98] = 9'b111111111;
assign f[32][99] = 9'b111111111;
assign f[32][100] = 9'b111111111;
assign f[32][101] = 9'b111111111;
assign f[32][102] = 9'b111111111;
assign f[32][103] = 9'b111111111;
assign f[32][104] = 9'b111111111;
assign f[32][105] = 9'b111111111;
assign f[32][106] = 9'b111111111;
assign f[32][107] = 9'b111111111;
assign f[32][108] = 9'b111111111;
assign f[32][109] = 9'b111111111;
assign f[32][110] = 9'b111111111;
assign f[32][117] = 9'b111111111;
assign f[32][118] = 9'b111111111;
assign f[32][119] = 9'b111111111;
assign f[32][120] = 9'b111111111;
assign f[32][121] = 9'b111111111;
assign f[32][122] = 9'b111111111;
assign f[32][123] = 9'b111111111;
assign f[32][145] = 9'b111111111;
assign f[32][146] = 9'b111111111;
assign f[32][147] = 9'b111111111;
assign f[32][148] = 9'b111111111;
assign f[32][149] = 9'b111111111;
assign f[32][150] = 9'b111111111;
assign f[32][151] = 9'b111111111;
assign f[32][152] = 9'b111111111;
assign f[32][153] = 9'b111111111;
assign f[32][154] = 9'b111111111;
assign f[32][164] = 9'b111111111;
assign f[32][165] = 9'b111111111;
assign f[32][166] = 9'b111111111;
assign f[32][167] = 9'b111111111;
assign f[32][168] = 9'b111111111;
assign f[32][169] = 9'b111111111;
assign f[32][170] = 9'b111111111;
assign f[32][171] = 9'b111111111;
assign f[32][172] = 9'b111111111;
assign f[32][179] = 9'b111111111;
assign f[32][180] = 9'b111111111;
assign f[32][181] = 9'b111111111;
assign f[32][182] = 9'b111111111;
assign f[32][183] = 9'b111111111;
assign f[32][184] = 9'b111111111;
assign f[32][185] = 9'b111111111;
assign f[33][19] = 9'b111111111;
assign f[33][20] = 9'b111111111;
assign f[33][21] = 9'b111111111;
assign f[33][22] = 9'b111111111;
assign f[33][23] = 9'b111111111;
assign f[33][24] = 9'b111111111;
assign f[33][25] = 9'b111111111;
assign f[33][26] = 9'b111111111;
assign f[33][27] = 9'b111111111;
assign f[33][28] = 9'b111111111;
assign f[33][29] = 9'b111111111;
assign f[33][30] = 9'b111111111;
assign f[33][31] = 9'b111111111;
assign f[33][32] = 9'b111111111;
assign f[33][33] = 9'b111111111;
assign f[33][34] = 9'b111111111;
assign f[33][35] = 9'b111111111;
assign f[33][36] = 9'b111111111;
assign f[33][37] = 9'b111111111;
assign f[33][38] = 9'b111111111;
assign f[33][39] = 9'b111111111;
assign f[33][40] = 9'b111111111;
assign f[33][42] = 9'b111111111;
assign f[33][43] = 9'b111111111;
assign f[33][44] = 9'b111111111;
assign f[33][45] = 9'b111111111;
assign f[33][46] = 9'b111111111;
assign f[33][47] = 9'b111111111;
assign f[33][48] = 9'b111111111;
assign f[33][56] = 9'b111111111;
assign f[33][57] = 9'b111111111;
assign f[33][58] = 9'b111111111;
assign f[33][59] = 9'b111111111;
assign f[33][60] = 9'b111111111;
assign f[33][61] = 9'b111111111;
assign f[33][62] = 9'b111111111;
assign f[33][66] = 9'b111111111;
assign f[33][67] = 9'b111111111;
assign f[33][68] = 9'b111111111;
assign f[33][69] = 9'b111111111;
assign f[33][70] = 9'b111111111;
assign f[33][71] = 9'b111111111;
assign f[33][72] = 9'b111111111;
assign f[33][73] = 9'b111111111;
assign f[33][74] = 9'b111111111;
assign f[33][75] = 9'b111111111;
assign f[33][76] = 9'b111111111;
assign f[33][77] = 9'b111111111;
assign f[33][78] = 9'b111111111;
assign f[33][79] = 9'b111111111;
assign f[33][80] = 9'b111111111;
assign f[33][81] = 9'b111111111;
assign f[33][94] = 9'b111111111;
assign f[33][95] = 9'b111111111;
assign f[33][96] = 9'b111111111;
assign f[33][97] = 9'b111111111;
assign f[33][98] = 9'b111111111;
assign f[33][99] = 9'b111111111;
assign f[33][100] = 9'b111111111;
assign f[33][101] = 9'b111111111;
assign f[33][102] = 9'b111111111;
assign f[33][103] = 9'b111111111;
assign f[33][104] = 9'b111111111;
assign f[33][105] = 9'b111111111;
assign f[33][106] = 9'b111111111;
assign f[33][107] = 9'b111111111;
assign f[33][108] = 9'b111111111;
assign f[33][109] = 9'b111111111;
assign f[33][110] = 9'b111111111;
assign f[33][111] = 9'b111111111;
assign f[33][117] = 9'b111111111;
assign f[33][118] = 9'b111111111;
assign f[33][119] = 9'b111111111;
assign f[33][120] = 9'b111111111;
assign f[33][121] = 9'b111111111;
assign f[33][122] = 9'b111111111;
assign f[33][123] = 9'b111111111;
assign f[33][145] = 9'b111111111;
assign f[33][146] = 9'b111111111;
assign f[33][147] = 9'b111111111;
assign f[33][148] = 9'b111111111;
assign f[33][149] = 9'b111111111;
assign f[33][150] = 9'b111111111;
assign f[33][151] = 9'b111111111;
assign f[33][152] = 9'b111111111;
assign f[33][153] = 9'b111111111;
assign f[33][154] = 9'b111111111;
assign f[33][164] = 9'b111111111;
assign f[33][165] = 9'b111111111;
assign f[33][166] = 9'b111111111;
assign f[33][167] = 9'b111111111;
assign f[33][168] = 9'b111111111;
assign f[33][169] = 9'b111111111;
assign f[33][170] = 9'b111111111;
assign f[33][171] = 9'b111111111;
assign f[33][172] = 9'b111111111;
assign f[33][173] = 9'b111111111;
assign f[33][179] = 9'b111111111;
assign f[33][180] = 9'b111111111;
assign f[33][181] = 9'b111111111;
assign f[33][182] = 9'b111111111;
assign f[33][183] = 9'b111111111;
assign f[33][184] = 9'b111111111;
assign f[33][185] = 9'b111111111;
assign f[34][19] = 9'b111111111;
assign f[34][20] = 9'b111111111;
assign f[34][21] = 9'b111111111;
assign f[34][22] = 9'b111111111;
assign f[34][23] = 9'b111111111;
assign f[34][24] = 9'b111111111;
assign f[34][25] = 9'b111111111;
assign f[34][26] = 9'b111111111;
assign f[34][27] = 9'b111111111;
assign f[34][28] = 9'b111111111;
assign f[34][29] = 9'b111111111;
assign f[34][30] = 9'b111111111;
assign f[34][31] = 9'b111111111;
assign f[34][32] = 9'b111111111;
assign f[34][33] = 9'b111111111;
assign f[34][34] = 9'b111111111;
assign f[34][35] = 9'b111111111;
assign f[34][36] = 9'b111111111;
assign f[34][37] = 9'b111111111;
assign f[34][38] = 9'b111111111;
assign f[34][39] = 9'b111111111;
assign f[34][40] = 9'b111111111;
assign f[34][42] = 9'b111111111;
assign f[34][43] = 9'b111111111;
assign f[34][44] = 9'b111111111;
assign f[34][45] = 9'b111111111;
assign f[34][46] = 9'b111111111;
assign f[34][47] = 9'b111111111;
assign f[34][48] = 9'b111111111;
assign f[34][56] = 9'b111111111;
assign f[34][57] = 9'b111111111;
assign f[34][58] = 9'b111111111;
assign f[34][59] = 9'b111111111;
assign f[34][60] = 9'b111111111;
assign f[34][61] = 9'b111111111;
assign f[34][62] = 9'b111111111;
assign f[34][65] = 9'b111111111;
assign f[34][66] = 9'b111111111;
assign f[34][67] = 9'b111111111;
assign f[34][68] = 9'b111111111;
assign f[34][69] = 9'b111111111;
assign f[34][70] = 9'b111111111;
assign f[34][71] = 9'b111111111;
assign f[34][72] = 9'b111111111;
assign f[34][73] = 9'b111111111;
assign f[34][74] = 9'b111111111;
assign f[34][75] = 9'b111111111;
assign f[34][76] = 9'b111111111;
assign f[34][77] = 9'b111111111;
assign f[34][78] = 9'b111111111;
assign f[34][79] = 9'b111111111;
assign f[34][80] = 9'b111111111;
assign f[34][81] = 9'b111111111;
assign f[34][94] = 9'b111111111;
assign f[34][95] = 9'b111111111;
assign f[34][96] = 9'b111111111;
assign f[34][97] = 9'b111111111;
assign f[34][98] = 9'b111111111;
assign f[34][99] = 9'b111111111;
assign f[34][100] = 9'b111111111;
assign f[34][101] = 9'b111111111;
assign f[34][102] = 9'b111111111;
assign f[34][103] = 9'b111111111;
assign f[34][104] = 9'b111111111;
assign f[34][105] = 9'b111111111;
assign f[34][106] = 9'b111111111;
assign f[34][107] = 9'b111111111;
assign f[34][108] = 9'b111111111;
assign f[34][109] = 9'b111111111;
assign f[34][110] = 9'b111111111;
assign f[34][111] = 9'b111111111;
assign f[34][112] = 9'b111111111;
assign f[34][117] = 9'b111111111;
assign f[34][118] = 9'b111111111;
assign f[34][119] = 9'b111111111;
assign f[34][120] = 9'b111111111;
assign f[34][121] = 9'b111111111;
assign f[34][122] = 9'b111111111;
assign f[34][123] = 9'b111111111;
assign f[34][146] = 9'b111111111;
assign f[34][147] = 9'b111111111;
assign f[34][148] = 9'b111111111;
assign f[34][149] = 9'b111111111;
assign f[34][150] = 9'b111111111;
assign f[34][151] = 9'b111111111;
assign f[34][152] = 9'b111111111;
assign f[34][153] = 9'b111111111;
assign f[34][154] = 9'b111111111;
assign f[34][164] = 9'b111111111;
assign f[34][165] = 9'b111111111;
assign f[34][166] = 9'b111111111;
assign f[34][167] = 9'b111111111;
assign f[34][168] = 9'b111111111;
assign f[34][169] = 9'b111111111;
assign f[34][170] = 9'b111111111;
assign f[34][171] = 9'b111111111;
assign f[34][172] = 9'b111111111;
assign f[34][173] = 9'b111111111;
assign f[34][179] = 9'b111111111;
assign f[34][180] = 9'b111111111;
assign f[34][181] = 9'b111111111;
assign f[34][182] = 9'b111111111;
assign f[34][183] = 9'b111111111;
assign f[34][184] = 9'b111111111;
assign f[34][185] = 9'b111111111;
assign f[35][19] = 9'b111111111;
assign f[35][20] = 9'b111111111;
assign f[35][21] = 9'b111111111;
assign f[35][22] = 9'b111111111;
assign f[35][23] = 9'b111111111;
assign f[35][24] = 9'b111111111;
assign f[35][25] = 9'b111111111;
assign f[35][26] = 9'b111111111;
assign f[35][27] = 9'b111111111;
assign f[35][28] = 9'b111111111;
assign f[35][29] = 9'b111111111;
assign f[35][30] = 9'b111111111;
assign f[35][31] = 9'b111111111;
assign f[35][32] = 9'b111111111;
assign f[35][33] = 9'b111111111;
assign f[35][34] = 9'b111111111;
assign f[35][35] = 9'b111111111;
assign f[35][36] = 9'b111111111;
assign f[35][37] = 9'b111111111;
assign f[35][38] = 9'b111111111;
assign f[35][39] = 9'b111111111;
assign f[35][42] = 9'b111111111;
assign f[35][43] = 9'b111111111;
assign f[35][44] = 9'b111111111;
assign f[35][45] = 9'b111111111;
assign f[35][46] = 9'b111111111;
assign f[35][47] = 9'b111111111;
assign f[35][48] = 9'b111111111;
assign f[35][56] = 9'b111111111;
assign f[35][57] = 9'b111111111;
assign f[35][58] = 9'b111111111;
assign f[35][59] = 9'b111111111;
assign f[35][60] = 9'b111111111;
assign f[35][61] = 9'b111111111;
assign f[35][62] = 9'b111111111;
assign f[35][65] = 9'b111111111;
assign f[35][66] = 9'b111111111;
assign f[35][67] = 9'b111111111;
assign f[35][68] = 9'b111111111;
assign f[35][69] = 9'b111111111;
assign f[35][70] = 9'b111111111;
assign f[35][71] = 9'b111111111;
assign f[35][72] = 9'b111111111;
assign f[35][73] = 9'b111111111;
assign f[35][74] = 9'b111111111;
assign f[35][75] = 9'b111111111;
assign f[35][76] = 9'b111111111;
assign f[35][77] = 9'b111111111;
assign f[35][78] = 9'b111111111;
assign f[35][79] = 9'b111111111;
assign f[35][80] = 9'b111111111;
assign f[35][81] = 9'b111111111;
assign f[35][94] = 9'b111111111;
assign f[35][95] = 9'b111111111;
assign f[35][96] = 9'b111111111;
assign f[35][97] = 9'b111111111;
assign f[35][98] = 9'b111111111;
assign f[35][99] = 9'b111111111;
assign f[35][100] = 9'b111111111;
assign f[35][101] = 9'b111111111;
assign f[35][102] = 9'b111111111;
assign f[35][103] = 9'b111111111;
assign f[35][104] = 9'b111111111;
assign f[35][105] = 9'b111111111;
assign f[35][106] = 9'b111111111;
assign f[35][107] = 9'b111111111;
assign f[35][108] = 9'b111111111;
assign f[35][109] = 9'b111111111;
assign f[35][110] = 9'b111111111;
assign f[35][111] = 9'b111111111;
assign f[35][112] = 9'b111111111;
assign f[35][117] = 9'b111111111;
assign f[35][118] = 9'b111111111;
assign f[35][119] = 9'b111111111;
assign f[35][120] = 9'b111111111;
assign f[35][121] = 9'b111111111;
assign f[35][122] = 9'b111111111;
assign f[35][123] = 9'b111111111;
assign f[35][144] = 9'b111111111;
assign f[35][145] = 9'b111111111;
assign f[35][146] = 9'b111111111;
assign f[35][147] = 9'b111111111;
assign f[35][148] = 9'b111111111;
assign f[35][149] = 9'b111111111;
assign f[35][150] = 9'b111111111;
assign f[35][151] = 9'b111111111;
assign f[35][152] = 9'b111111111;
assign f[35][153] = 9'b111111111;
assign f[35][154] = 9'b111111111;
assign f[35][163] = 9'b111111111;
assign f[35][164] = 9'b111111111;
assign f[35][165] = 9'b111111111;
assign f[35][166] = 9'b111111111;
assign f[35][167] = 9'b111111111;
assign f[35][168] = 9'b111111111;
assign f[35][169] = 9'b111111111;
assign f[35][170] = 9'b111111111;
assign f[35][171] = 9'b111111111;
assign f[35][172] = 9'b111111111;
assign f[35][173] = 9'b111111111;
assign f[35][179] = 9'b111111111;
assign f[35][180] = 9'b111111111;
assign f[35][181] = 9'b111111111;
assign f[35][182] = 9'b111111111;
assign f[35][183] = 9'b111111111;
assign f[35][184] = 9'b111111111;
assign f[35][185] = 9'b111111111;
assign f[36][19] = 9'b111111111;
assign f[36][20] = 9'b111111111;
assign f[36][21] = 9'b111111111;
assign f[36][22] = 9'b111111111;
assign f[36][23] = 9'b111111111;
assign f[36][24] = 9'b111111111;
assign f[36][25] = 9'b111111111;
assign f[36][26] = 9'b111111111;
assign f[36][27] = 9'b111111111;
assign f[36][28] = 9'b111111111;
assign f[36][29] = 9'b111111111;
assign f[36][30] = 9'b111111111;
assign f[36][31] = 9'b111111111;
assign f[36][32] = 9'b111111111;
assign f[36][33] = 9'b111111111;
assign f[36][34] = 9'b111111111;
assign f[36][35] = 9'b111111111;
assign f[36][36] = 9'b111111111;
assign f[36][37] = 9'b111111111;
assign f[36][38] = 9'b111111111;
assign f[36][39] = 9'b111111111;
assign f[36][42] = 9'b111111111;
assign f[36][43] = 9'b111111111;
assign f[36][44] = 9'b111111111;
assign f[36][45] = 9'b111111111;
assign f[36][46] = 9'b111111111;
assign f[36][47] = 9'b111111111;
assign f[36][48] = 9'b111111111;
assign f[36][56] = 9'b111111111;
assign f[36][57] = 9'b111111111;
assign f[36][58] = 9'b111111111;
assign f[36][59] = 9'b111111111;
assign f[36][60] = 9'b111111111;
assign f[36][61] = 9'b111111111;
assign f[36][62] = 9'b111111111;
assign f[36][65] = 9'b111111111;
assign f[36][66] = 9'b111111111;
assign f[36][67] = 9'b111111111;
assign f[36][68] = 9'b111111111;
assign f[36][69] = 9'b111111111;
assign f[36][70] = 9'b111111111;
assign f[36][71] = 9'b111111111;
assign f[36][72] = 9'b111111111;
assign f[36][73] = 9'b111111111;
assign f[36][74] = 9'b111111111;
assign f[36][75] = 9'b111111111;
assign f[36][76] = 9'b111111111;
assign f[36][77] = 9'b111111111;
assign f[36][78] = 9'b111111111;
assign f[36][79] = 9'b111111111;
assign f[36][80] = 9'b111111111;
assign f[36][94] = 9'b111111111;
assign f[36][95] = 9'b111111111;
assign f[36][96] = 9'b111111111;
assign f[36][97] = 9'b111111111;
assign f[36][98] = 9'b111111111;
assign f[36][99] = 9'b111111111;
assign f[36][100] = 9'b111111111;
assign f[36][101] = 9'b111111111;
assign f[36][102] = 9'b111111111;
assign f[36][103] = 9'b111111111;
assign f[36][104] = 9'b111111111;
assign f[36][105] = 9'b111111111;
assign f[36][106] = 9'b111111111;
assign f[36][107] = 9'b111111111;
assign f[36][108] = 9'b111111111;
assign f[36][109] = 9'b111111111;
assign f[36][110] = 9'b111111111;
assign f[36][111] = 9'b111111111;
assign f[36][112] = 9'b111111111;
assign f[36][113] = 9'b111111111;
assign f[36][117] = 9'b111111111;
assign f[36][118] = 9'b111111111;
assign f[36][119] = 9'b111111111;
assign f[36][120] = 9'b111111111;
assign f[36][121] = 9'b111111111;
assign f[36][122] = 9'b111111111;
assign f[36][123] = 9'b111111111;
assign f[36][144] = 9'b111111111;
assign f[36][145] = 9'b111111111;
assign f[36][146] = 9'b111111111;
assign f[36][147] = 9'b111111111;
assign f[36][148] = 9'b111111111;
assign f[36][149] = 9'b111111111;
assign f[36][150] = 9'b111111111;
assign f[36][151] = 9'b111111111;
assign f[36][152] = 9'b111111111;
assign f[36][153] = 9'b111111111;
assign f[36][154] = 9'b111111111;
assign f[36][163] = 9'b111111111;
assign f[36][164] = 9'b111111111;
assign f[36][165] = 9'b111111111;
assign f[36][166] = 9'b111111111;
assign f[36][167] = 9'b111111111;
assign f[36][168] = 9'b111111111;
assign f[36][169] = 9'b111111111;
assign f[36][170] = 9'b111111111;
assign f[36][171] = 9'b111111111;
assign f[36][172] = 9'b111111111;
assign f[36][173] = 9'b111111111;
assign f[36][180] = 9'b111111111;
assign f[36][181] = 9'b111111111;
assign f[36][182] = 9'b111111111;
assign f[36][183] = 9'b111111111;
assign f[36][184] = 9'b111111111;
assign f[36][185] = 9'b111111111;
assign f[37][26] = 9'b111111111;
assign f[37][27] = 9'b111111111;
assign f[37][28] = 9'b111111111;
assign f[37][29] = 9'b111111111;
assign f[37][30] = 9'b111111111;
assign f[37][31] = 9'b111111111;
assign f[37][32] = 9'b111111111;
assign f[37][42] = 9'b111111111;
assign f[37][43] = 9'b111111111;
assign f[37][44] = 9'b111111111;
assign f[37][45] = 9'b111111111;
assign f[37][46] = 9'b111111111;
assign f[37][47] = 9'b111111111;
assign f[37][48] = 9'b111111111;
assign f[37][56] = 9'b111111111;
assign f[37][57] = 9'b111111111;
assign f[37][58] = 9'b111111111;
assign f[37][59] = 9'b111111111;
assign f[37][60] = 9'b111111111;
assign f[37][61] = 9'b111111111;
assign f[37][62] = 9'b111111111;
assign f[37][65] = 9'b111111111;
assign f[37][66] = 9'b111111111;
assign f[37][67] = 9'b111111111;
assign f[37][68] = 9'b111111111;
assign f[37][69] = 9'b111111111;
assign f[37][70] = 9'b111111111;
assign f[37][71] = 9'b111111111;
assign f[37][94] = 9'b111111111;
assign f[37][95] = 9'b111111111;
assign f[37][96] = 9'b111111111;
assign f[37][97] = 9'b111111111;
assign f[37][98] = 9'b111111111;
assign f[37][99] = 9'b111111111;
assign f[37][100] = 9'b111111111;
assign f[37][106] = 9'b111111111;
assign f[37][107] = 9'b111111111;
assign f[37][108] = 9'b111111111;
assign f[37][109] = 9'b111111111;
assign f[37][110] = 9'b111111111;
assign f[37][111] = 9'b111111111;
assign f[37][112] = 9'b111111111;
assign f[37][113] = 9'b111111111;
assign f[37][117] = 9'b111111111;
assign f[37][118] = 9'b111111111;
assign f[37][119] = 9'b111111111;
assign f[37][120] = 9'b111111111;
assign f[37][121] = 9'b111111111;
assign f[37][122] = 9'b111111111;
assign f[37][123] = 9'b111111111;
assign f[37][144] = 9'b111111111;
assign f[37][145] = 9'b111111111;
assign f[37][146] = 9'b111111111;
assign f[37][147] = 9'b111111111;
assign f[37][148] = 9'b111111111;
assign f[37][149] = 9'b111111111;
assign f[37][150] = 9'b111111111;
assign f[37][151] = 9'b111111111;
assign f[37][152] = 9'b111111111;
assign f[37][153] = 9'b111111111;
assign f[37][154] = 9'b111111111;
assign f[37][155] = 9'b111111111;
assign f[37][163] = 9'b111111111;
assign f[37][164] = 9'b111111111;
assign f[37][165] = 9'b111111111;
assign f[37][166] = 9'b111111111;
assign f[37][167] = 9'b111111111;
assign f[37][168] = 9'b111111111;
assign f[37][169] = 9'b111111111;
assign f[37][170] = 9'b111111111;
assign f[37][171] = 9'b111111111;
assign f[37][172] = 9'b111111111;
assign f[37][173] = 9'b111111111;
assign f[37][174] = 9'b111111111;
assign f[37][180] = 9'b111111111;
assign f[37][181] = 9'b111111111;
assign f[37][182] = 9'b111111111;
assign f[37][183] = 9'b111111111;
assign f[37][184] = 9'b111111111;
assign f[37][185] = 9'b111111111;
assign f[38][26] = 9'b111111111;
assign f[38][27] = 9'b111111111;
assign f[38][28] = 9'b111111111;
assign f[38][29] = 9'b111111111;
assign f[38][30] = 9'b111111111;
assign f[38][31] = 9'b111111111;
assign f[38][32] = 9'b111111111;
assign f[38][42] = 9'b111111111;
assign f[38][43] = 9'b111111111;
assign f[38][44] = 9'b111111111;
assign f[38][45] = 9'b111111111;
assign f[38][46] = 9'b111111111;
assign f[38][47] = 9'b111111111;
assign f[38][48] = 9'b111111111;
assign f[38][56] = 9'b111111111;
assign f[38][57] = 9'b111111111;
assign f[38][58] = 9'b111111111;
assign f[38][59] = 9'b111111111;
assign f[38][60] = 9'b111111111;
assign f[38][61] = 9'b111111111;
assign f[38][62] = 9'b111111111;
assign f[38][65] = 9'b111111111;
assign f[38][66] = 9'b111111111;
assign f[38][67] = 9'b111111111;
assign f[38][68] = 9'b111111111;
assign f[38][69] = 9'b111111111;
assign f[38][70] = 9'b111111111;
assign f[38][71] = 9'b111111111;
assign f[38][94] = 9'b111111111;
assign f[38][95] = 9'b111111111;
assign f[38][96] = 9'b111111111;
assign f[38][97] = 9'b111111111;
assign f[38][98] = 9'b111111111;
assign f[38][99] = 9'b111111111;
assign f[38][100] = 9'b111111111;
assign f[38][107] = 9'b111111111;
assign f[38][108] = 9'b111111111;
assign f[38][109] = 9'b111111111;
assign f[38][110] = 9'b111111111;
assign f[38][111] = 9'b111111111;
assign f[38][112] = 9'b111111111;
assign f[38][113] = 9'b111111111;
assign f[38][117] = 9'b111111111;
assign f[38][118] = 9'b111111111;
assign f[38][119] = 9'b111111111;
assign f[38][120] = 9'b111111111;
assign f[38][121] = 9'b111111111;
assign f[38][122] = 9'b111111111;
assign f[38][123] = 9'b111111111;
assign f[38][143] = 9'b111111111;
assign f[38][144] = 9'b111111111;
assign f[38][145] = 9'b111111111;
assign f[38][146] = 9'b111111111;
assign f[38][147] = 9'b111111111;
assign f[38][148] = 9'b111111111;
assign f[38][150] = 9'b111111111;
assign f[38][151] = 9'b111111111;
assign f[38][152] = 9'b111111111;
assign f[38][153] = 9'b111111111;
assign f[38][154] = 9'b111111111;
assign f[38][155] = 9'b111111111;
assign f[38][163] = 9'b111111111;
assign f[38][164] = 9'b111111111;
assign f[38][165] = 9'b111111111;
assign f[38][166] = 9'b111111111;
assign f[38][167] = 9'b111111111;
assign f[38][168] = 9'b111111111;
assign f[38][169] = 9'b111111111;
assign f[38][170] = 9'b111111111;
assign f[38][171] = 9'b111111111;
assign f[38][172] = 9'b111111111;
assign f[38][173] = 9'b111111111;
assign f[38][174] = 9'b111111111;
assign f[38][180] = 9'b111111111;
assign f[38][181] = 9'b111111111;
assign f[38][182] = 9'b111111111;
assign f[38][183] = 9'b111111111;
assign f[38][184] = 9'b111111111;
assign f[38][185] = 9'b111111111;
assign f[39][26] = 9'b111111111;
assign f[39][27] = 9'b111111111;
assign f[39][28] = 9'b111111111;
assign f[39][29] = 9'b111111111;
assign f[39][30] = 9'b111111111;
assign f[39][31] = 9'b111111111;
assign f[39][32] = 9'b111111111;
assign f[39][42] = 9'b111111111;
assign f[39][43] = 9'b111111111;
assign f[39][44] = 9'b111111111;
assign f[39][45] = 9'b111111111;
assign f[39][46] = 9'b111111111;
assign f[39][47] = 9'b111111111;
assign f[39][48] = 9'b111111111;
assign f[39][56] = 9'b111111111;
assign f[39][57] = 9'b111111111;
assign f[39][58] = 9'b111111111;
assign f[39][59] = 9'b111111111;
assign f[39][60] = 9'b111111111;
assign f[39][61] = 9'b111111111;
assign f[39][62] = 9'b111111111;
assign f[39][65] = 9'b111111111;
assign f[39][66] = 9'b111111111;
assign f[39][67] = 9'b111111111;
assign f[39][68] = 9'b111111111;
assign f[39][69] = 9'b111111111;
assign f[39][70] = 9'b111111111;
assign f[39][71] = 9'b111111111;
assign f[39][94] = 9'b111111111;
assign f[39][95] = 9'b111111111;
assign f[39][96] = 9'b111111111;
assign f[39][97] = 9'b111111111;
assign f[39][98] = 9'b111111111;
assign f[39][99] = 9'b111111111;
assign f[39][100] = 9'b111111111;
assign f[39][107] = 9'b111111111;
assign f[39][108] = 9'b111111111;
assign f[39][109] = 9'b111111111;
assign f[39][110] = 9'b111111111;
assign f[39][111] = 9'b111111111;
assign f[39][112] = 9'b111111111;
assign f[39][113] = 9'b111111111;
assign f[39][117] = 9'b111111111;
assign f[39][118] = 9'b111111111;
assign f[39][119] = 9'b111111111;
assign f[39][120] = 9'b111111111;
assign f[39][121] = 9'b111111111;
assign f[39][122] = 9'b111111111;
assign f[39][123] = 9'b111111111;
assign f[39][143] = 9'b111111111;
assign f[39][144] = 9'b111111111;
assign f[39][147] = 9'b111111111;
assign f[39][148] = 9'b111111111;
assign f[39][150] = 9'b111111111;
assign f[39][151] = 9'b111111111;
assign f[39][152] = 9'b111111111;
assign f[39][153] = 9'b111111111;
assign f[39][154] = 9'b111111111;
assign f[39][155] = 9'b111111111;
assign f[39][163] = 9'b111111111;
assign f[39][164] = 9'b111111111;
assign f[39][165] = 9'b111111111;
assign f[39][166] = 9'b111111111;
assign f[39][167] = 9'b111111111;
assign f[39][168] = 9'b111111111;
assign f[39][169] = 9'b111111111;
assign f[39][170] = 9'b111111111;
assign f[39][171] = 9'b111111111;
assign f[39][172] = 9'b111111111;
assign f[39][173] = 9'b111111111;
assign f[39][174] = 9'b111111111;
assign f[39][180] = 9'b111111111;
assign f[39][181] = 9'b111111111;
assign f[39][183] = 9'b111111111;
assign f[39][184] = 9'b111111111;
assign f[39][185] = 9'b111111111;
assign f[40][26] = 9'b111111111;
assign f[40][27] = 9'b111111111;
assign f[40][28] = 9'b111111111;
assign f[40][29] = 9'b111111111;
assign f[40][30] = 9'b111111111;
assign f[40][31] = 9'b111111111;
assign f[40][32] = 9'b111111111;
assign f[40][33] = 9'b111111111;
assign f[40][42] = 9'b111111111;
assign f[40][43] = 9'b111111111;
assign f[40][44] = 9'b111111111;
assign f[40][45] = 9'b111111111;
assign f[40][46] = 9'b111111111;
assign f[40][47] = 9'b111111111;
assign f[40][48] = 9'b111111111;
assign f[40][56] = 9'b111111111;
assign f[40][57] = 9'b111111111;
assign f[40][58] = 9'b111111111;
assign f[40][59] = 9'b111111111;
assign f[40][60] = 9'b111111111;
assign f[40][61] = 9'b111111111;
assign f[40][62] = 9'b111111111;
assign f[40][65] = 9'b111111111;
assign f[40][66] = 9'b111111111;
assign f[40][67] = 9'b111111111;
assign f[40][68] = 9'b111111111;
assign f[40][69] = 9'b111111111;
assign f[40][70] = 9'b111111111;
assign f[40][71] = 9'b111111111;
assign f[40][94] = 9'b111111111;
assign f[40][95] = 9'b111111111;
assign f[40][96] = 9'b111111111;
assign f[40][97] = 9'b111111111;
assign f[40][98] = 9'b111111111;
assign f[40][99] = 9'b111111111;
assign f[40][100] = 9'b111111111;
assign f[40][107] = 9'b111111111;
assign f[40][108] = 9'b111111111;
assign f[40][109] = 9'b111111111;
assign f[40][110] = 9'b111111111;
assign f[40][111] = 9'b111111111;
assign f[40][112] = 9'b111111111;
assign f[40][113] = 9'b111111111;
assign f[40][117] = 9'b111111111;
assign f[40][118] = 9'b111111111;
assign f[40][119] = 9'b111111111;
assign f[40][120] = 9'b111111111;
assign f[40][121] = 9'b111111111;
assign f[40][122] = 9'b111111111;
assign f[40][123] = 9'b111111111;
assign f[40][143] = 9'b111111111;
assign f[40][144] = 9'b111111111;
assign f[40][145] = 9'b111111111;
assign f[40][146] = 9'b111111111;
assign f[40][147] = 9'b111111111;
assign f[40][148] = 9'b111111111;
assign f[40][150] = 9'b111111111;
assign f[40][151] = 9'b111111111;
assign f[40][152] = 9'b111111111;
assign f[40][153] = 9'b111111111;
assign f[40][154] = 9'b111111111;
assign f[40][155] = 9'b111111111;
assign f[40][163] = 9'b111111111;
assign f[40][164] = 9'b111111111;
assign f[40][165] = 9'b111111111;
assign f[40][166] = 9'b111111111;
assign f[40][167] = 9'b111111111;
assign f[40][168] = 9'b111111111;
assign f[40][169] = 9'b111111111;
assign f[40][170] = 9'b111111111;
assign f[40][171] = 9'b111111111;
assign f[40][172] = 9'b111111111;
assign f[40][173] = 9'b111111111;
assign f[40][174] = 9'b111111111;
assign f[40][175] = 9'b111111111;
assign f[40][180] = 9'b111111111;
assign f[40][181] = 9'b111111111;
assign f[40][182] = 9'b111111111;
assign f[40][183] = 9'b111111111;
assign f[40][184] = 9'b111111111;
assign f[40][185] = 9'b111111111;
assign f[41][26] = 9'b111111111;
assign f[41][27] = 9'b111111111;
assign f[41][28] = 9'b111111111;
assign f[41][29] = 9'b111111111;
assign f[41][30] = 9'b111111111;
assign f[41][31] = 9'b111111111;
assign f[41][32] = 9'b111111111;
assign f[41][42] = 9'b111111111;
assign f[41][43] = 9'b111111111;
assign f[41][44] = 9'b111111111;
assign f[41][45] = 9'b111111111;
assign f[41][47] = 9'b111111111;
assign f[41][48] = 9'b111111111;
assign f[41][56] = 9'b111111111;
assign f[41][57] = 9'b111111111;
assign f[41][58] = 9'b111111111;
assign f[41][59] = 9'b111111111;
assign f[41][60] = 9'b111111111;
assign f[41][61] = 9'b111111111;
assign f[41][62] = 9'b111111111;
assign f[41][65] = 9'b111111111;
assign f[41][66] = 9'b111111111;
assign f[41][67] = 9'b111111111;
assign f[41][68] = 9'b111111111;
assign f[41][69] = 9'b111111111;
assign f[41][70] = 9'b111111111;
assign f[41][71] = 9'b111111111;
assign f[41][94] = 9'b111111111;
assign f[41][95] = 9'b111111111;
assign f[41][96] = 9'b111111111;
assign f[41][97] = 9'b111111111;
assign f[41][98] = 9'b111111111;
assign f[41][99] = 9'b111111111;
assign f[41][100] = 9'b111111111;
assign f[41][107] = 9'b111111111;
assign f[41][108] = 9'b111111111;
assign f[41][109] = 9'b111111111;
assign f[41][110] = 9'b111111111;
assign f[41][111] = 9'b111111111;
assign f[41][112] = 9'b111111111;
assign f[41][113] = 9'b111111111;
assign f[41][117] = 9'b111111111;
assign f[41][118] = 9'b111111111;
assign f[41][119] = 9'b111111111;
assign f[41][120] = 9'b111111111;
assign f[41][121] = 9'b111111111;
assign f[41][122] = 9'b111111111;
assign f[41][123] = 9'b111111111;
assign f[41][142] = 9'b111111111;
assign f[41][143] = 9'b111111111;
assign f[41][146] = 9'b111111111;
assign f[41][147] = 9'b111111111;
assign f[41][148] = 9'b111111111;
assign f[41][150] = 9'b111111111;
assign f[41][151] = 9'b111111111;
assign f[41][152] = 9'b111111111;
assign f[41][153] = 9'b111111111;
assign f[41][154] = 9'b111111111;
assign f[41][155] = 9'b111111111;
assign f[41][156] = 9'b111111111;
assign f[41][163] = 9'b111111111;
assign f[41][164] = 9'b111111111;
assign f[41][165] = 9'b111111111;
assign f[41][166] = 9'b111111111;
assign f[41][167] = 9'b111111111;
assign f[41][168] = 9'b111111111;
assign f[41][169] = 9'b111111111;
assign f[41][170] = 9'b111111111;
assign f[41][171] = 9'b111111111;
assign f[41][172] = 9'b111111111;
assign f[41][173] = 9'b111111111;
assign f[41][174] = 9'b111111111;
assign f[41][175] = 9'b111111111;
assign f[41][180] = 9'b111111111;
assign f[41][181] = 9'b111111111;
assign f[41][182] = 9'b111111111;
assign f[41][183] = 9'b111111111;
assign f[41][184] = 9'b111111111;
assign f[41][185] = 9'b111111111;
assign f[42][26] = 9'b111111111;
assign f[42][27] = 9'b111111111;
assign f[42][28] = 9'b111111111;
assign f[42][29] = 9'b111111111;
assign f[42][30] = 9'b111111111;
assign f[42][31] = 9'b111111111;
assign f[42][32] = 9'b111111111;
assign f[42][42] = 9'b111111111;
assign f[42][43] = 9'b111111111;
assign f[42][44] = 9'b111111111;
assign f[42][45] = 9'b111111111;
assign f[42][46] = 9'b111111111;
assign f[42][47] = 9'b111111111;
assign f[42][48] = 9'b111111111;
assign f[42][56] = 9'b111111111;
assign f[42][57] = 9'b111111111;
assign f[42][58] = 9'b111111111;
assign f[42][59] = 9'b111111111;
assign f[42][60] = 9'b111111111;
assign f[42][61] = 9'b111111111;
assign f[42][62] = 9'b111111111;
assign f[42][65] = 9'b111111111;
assign f[42][66] = 9'b111111111;
assign f[42][67] = 9'b111111111;
assign f[42][68] = 9'b111111111;
assign f[42][69] = 9'b111111111;
assign f[42][70] = 9'b111111111;
assign f[42][71] = 9'b111111111;
assign f[42][94] = 9'b111111111;
assign f[42][95] = 9'b111111111;
assign f[42][96] = 9'b111111111;
assign f[42][97] = 9'b111111111;
assign f[42][98] = 9'b111111111;
assign f[42][99] = 9'b111111111;
assign f[42][100] = 9'b111111111;
assign f[42][107] = 9'b111111111;
assign f[42][108] = 9'b111111111;
assign f[42][109] = 9'b111111111;
assign f[42][110] = 9'b111111111;
assign f[42][111] = 9'b111111111;
assign f[42][112] = 9'b111111111;
assign f[42][113] = 9'b111111111;
assign f[42][117] = 9'b111111111;
assign f[42][118] = 9'b111111111;
assign f[42][119] = 9'b111111111;
assign f[42][120] = 9'b111111111;
assign f[42][121] = 9'b111111111;
assign f[42][122] = 9'b111111111;
assign f[42][123] = 9'b111111111;
assign f[42][142] = 9'b111111111;
assign f[42][143] = 9'b111111111;
assign f[42][146] = 9'b111111111;
assign f[42][147] = 9'b111111111;
assign f[42][151] = 9'b111111111;
assign f[42][152] = 9'b111111111;
assign f[42][153] = 9'b111111111;
assign f[42][154] = 9'b111111111;
assign f[42][155] = 9'b111111111;
assign f[42][156] = 9'b111111111;
assign f[42][163] = 9'b111111111;
assign f[42][164] = 9'b111111111;
assign f[42][165] = 9'b111111111;
assign f[42][166] = 9'b111111111;
assign f[42][167] = 9'b111111111;
assign f[42][168] = 9'b111111111;
assign f[42][169] = 9'b111111111;
assign f[42][170] = 9'b111111111;
assign f[42][171] = 9'b111111111;
assign f[42][172] = 9'b111111111;
assign f[42][173] = 9'b111111111;
assign f[42][174] = 9'b111111111;
assign f[42][175] = 9'b111111111;
assign f[42][180] = 9'b111111111;
assign f[42][181] = 9'b111111111;
assign f[42][182] = 9'b111111111;
assign f[42][183] = 9'b111111111;
assign f[42][184] = 9'b111111111;
assign f[42][185] = 9'b111111111;
assign f[43][26] = 9'b111111111;
assign f[43][27] = 9'b111111111;
assign f[43][28] = 9'b111111111;
assign f[43][29] = 9'b111111111;
assign f[43][30] = 9'b111111111;
assign f[43][31] = 9'b111111111;
assign f[43][32] = 9'b111111111;
assign f[43][42] = 9'b111111111;
assign f[43][43] = 9'b111111111;
assign f[43][44] = 9'b111111111;
assign f[43][45] = 9'b111111111;
assign f[43][46] = 9'b111111111;
assign f[43][47] = 9'b111111111;
assign f[43][48] = 9'b111111111;
assign f[43][56] = 9'b111111111;
assign f[43][57] = 9'b111111111;
assign f[43][58] = 9'b111111111;
assign f[43][59] = 9'b111111111;
assign f[43][60] = 9'b111111111;
assign f[43][61] = 9'b111111111;
assign f[43][62] = 9'b111111111;
assign f[43][65] = 9'b111111111;
assign f[43][66] = 9'b111111111;
assign f[43][67] = 9'b111111111;
assign f[43][68] = 9'b111111111;
assign f[43][69] = 9'b111111111;
assign f[43][70] = 9'b111111111;
assign f[43][71] = 9'b111111111;
assign f[43][94] = 9'b111111111;
assign f[43][95] = 9'b111111111;
assign f[43][96] = 9'b111111111;
assign f[43][97] = 9'b111111111;
assign f[43][98] = 9'b111111111;
assign f[43][99] = 9'b111111111;
assign f[43][100] = 9'b111111111;
assign f[43][107] = 9'b111111111;
assign f[43][108] = 9'b111111111;
assign f[43][109] = 9'b111111111;
assign f[43][110] = 9'b111111111;
assign f[43][111] = 9'b111111111;
assign f[43][112] = 9'b111111111;
assign f[43][113] = 9'b111111111;
assign f[43][117] = 9'b111111111;
assign f[43][118] = 9'b111111111;
assign f[43][119] = 9'b111111111;
assign f[43][120] = 9'b111111111;
assign f[43][121] = 9'b111111111;
assign f[43][122] = 9'b111111111;
assign f[43][123] = 9'b111111111;
assign f[43][143] = 9'b111111111;
assign f[43][144] = 9'b111111111;
assign f[43][150] = 9'b111111111;
assign f[43][151] = 9'b111111111;
assign f[43][152] = 9'b111111111;
assign f[43][153] = 9'b111111111;
assign f[43][154] = 9'b111111111;
assign f[43][155] = 9'b111111111;
assign f[43][156] = 9'b111111111;
assign f[43][163] = 9'b111111111;
assign f[43][164] = 9'b111111111;
assign f[43][165] = 9'b111111111;
assign f[43][166] = 9'b111111111;
assign f[43][167] = 9'b111111111;
assign f[43][168] = 9'b111111111;
assign f[43][170] = 9'b111111111;
assign f[43][171] = 9'b111111111;
assign f[43][172] = 9'b111111111;
assign f[43][173] = 9'b111111111;
assign f[43][174] = 9'b111111111;
assign f[43][175] = 9'b111111111;
assign f[43][180] = 9'b111111111;
assign f[43][181] = 9'b111111111;
assign f[43][182] = 9'b111111111;
assign f[43][183] = 9'b111111111;
assign f[43][184] = 9'b111111111;
assign f[43][185] = 9'b111111111;
assign f[44][26] = 9'b111111111;
assign f[44][27] = 9'b111111111;
assign f[44][28] = 9'b111111111;
assign f[44][29] = 9'b111111111;
assign f[44][30] = 9'b111111111;
assign f[44][31] = 9'b111111111;
assign f[44][32] = 9'b111111111;
assign f[44][42] = 9'b111111111;
assign f[44][43] = 9'b111111111;
assign f[44][44] = 9'b111111111;
assign f[44][45] = 9'b111111111;
assign f[44][46] = 9'b111111111;
assign f[44][47] = 9'b111111111;
assign f[44][48] = 9'b111111111;
assign f[44][55] = 9'b111111111;
assign f[44][56] = 9'b111111111;
assign f[44][57] = 9'b111111111;
assign f[44][58] = 9'b111111111;
assign f[44][59] = 9'b111111111;
assign f[44][60] = 9'b111111111;
assign f[44][61] = 9'b111111111;
assign f[44][62] = 9'b111111111;
assign f[44][65] = 9'b111111111;
assign f[44][66] = 9'b111111111;
assign f[44][67] = 9'b111111111;
assign f[44][68] = 9'b111111111;
assign f[44][69] = 9'b111111111;
assign f[44][70] = 9'b111111111;
assign f[44][71] = 9'b111111111;
assign f[44][94] = 9'b111111111;
assign f[44][95] = 9'b111111111;
assign f[44][96] = 9'b111111111;
assign f[44][97] = 9'b111111111;
assign f[44][98] = 9'b111111111;
assign f[44][99] = 9'b111111111;
assign f[44][100] = 9'b111111111;
assign f[44][107] = 9'b111111111;
assign f[44][108] = 9'b111111111;
assign f[44][109] = 9'b111111111;
assign f[44][110] = 9'b111111111;
assign f[44][111] = 9'b111111111;
assign f[44][112] = 9'b111111111;
assign f[44][113] = 9'b111111111;
assign f[44][117] = 9'b111111111;
assign f[44][118] = 9'b111111111;
assign f[44][119] = 9'b111111111;
assign f[44][120] = 9'b111111111;
assign f[44][121] = 9'b111111111;
assign f[44][122] = 9'b111111111;
assign f[44][123] = 9'b111111111;
assign f[44][142] = 9'b111111111;
assign f[44][143] = 9'b111111111;
assign f[44][144] = 9'b111111111;
assign f[44][145] = 9'b111111111;
assign f[44][146] = 9'b111111111;
assign f[44][151] = 9'b111111111;
assign f[44][152] = 9'b111111111;
assign f[44][153] = 9'b111111111;
assign f[44][154] = 9'b111111111;
assign f[44][155] = 9'b111111111;
assign f[44][156] = 9'b111111111;
assign f[44][164] = 9'b111111111;
assign f[44][165] = 9'b111111111;
assign f[44][166] = 9'b111111111;
assign f[44][167] = 9'b111111111;
assign f[44][168] = 9'b111111111;
assign f[44][170] = 9'b111111111;
assign f[44][171] = 9'b111111111;
assign f[44][172] = 9'b111111111;
assign f[44][173] = 9'b111111111;
assign f[44][174] = 9'b111111111;
assign f[44][175] = 9'b111111111;
assign f[44][176] = 9'b111111111;
assign f[44][180] = 9'b111111111;
assign f[44][181] = 9'b111111111;
assign f[44][182] = 9'b111111111;
assign f[44][183] = 9'b111111111;
assign f[44][184] = 9'b111111111;
assign f[44][185] = 9'b111111111;
assign f[45][26] = 9'b111111111;
assign f[45][27] = 9'b111111111;
assign f[45][28] = 9'b111111111;
assign f[45][29] = 9'b111111111;
assign f[45][30] = 9'b111111111;
assign f[45][31] = 9'b111111111;
assign f[45][32] = 9'b111111111;
assign f[45][42] = 9'b111111111;
assign f[45][43] = 9'b111111111;
assign f[45][44] = 9'b111111111;
assign f[45][45] = 9'b111111111;
assign f[45][46] = 9'b111111111;
assign f[45][47] = 9'b111111111;
assign f[45][48] = 9'b111111111;
assign f[45][49] = 9'b111111111;
assign f[45][50] = 9'b111111111;
assign f[45][51] = 9'b111111111;
assign f[45][52] = 9'b111111111;
assign f[45][54] = 9'b111111111;
assign f[45][55] = 9'b111111111;
assign f[45][56] = 9'b111111111;
assign f[45][57] = 9'b111111111;
assign f[45][58] = 9'b111111111;
assign f[45][59] = 9'b111111111;
assign f[45][60] = 9'b111111111;
assign f[45][61] = 9'b111111111;
assign f[45][62] = 9'b111111111;
assign f[45][65] = 9'b111111111;
assign f[45][66] = 9'b111111111;
assign f[45][67] = 9'b111111111;
assign f[45][68] = 9'b111111111;
assign f[45][69] = 9'b111111111;
assign f[45][70] = 9'b111111111;
assign f[45][71] = 9'b111111111;
assign f[45][72] = 9'b111111111;
assign f[45][73] = 9'b111111111;
assign f[45][74] = 9'b111111111;
assign f[45][75] = 9'b111111111;
assign f[45][76] = 9'b111111111;
assign f[45][77] = 9'b111111111;
assign f[45][78] = 9'b111111111;
assign f[45][79] = 9'b111111111;
assign f[45][80] = 9'b111111111;
assign f[45][94] = 9'b111111111;
assign f[45][95] = 9'b111111111;
assign f[45][96] = 9'b111111111;
assign f[45][97] = 9'b111111111;
assign f[45][98] = 9'b111111111;
assign f[45][99] = 9'b111111111;
assign f[45][100] = 9'b111111111;
assign f[45][107] = 9'b111111111;
assign f[45][108] = 9'b111111111;
assign f[45][109] = 9'b111111111;
assign f[45][110] = 9'b111111111;
assign f[45][111] = 9'b111111111;
assign f[45][112] = 9'b111111111;
assign f[45][113] = 9'b111111111;
assign f[45][117] = 9'b111111111;
assign f[45][118] = 9'b111111111;
assign f[45][120] = 9'b111111111;
assign f[45][121] = 9'b111111111;
assign f[45][122] = 9'b111111111;
assign f[45][123] = 9'b111111111;
assign f[45][142] = 9'b111111111;
assign f[45][143] = 9'b111111111;
assign f[45][144] = 9'b111111111;
assign f[45][145] = 9'b111111111;
assign f[45][146] = 9'b111111111;
assign f[45][151] = 9'b111111111;
assign f[45][152] = 9'b111111111;
assign f[45][153] = 9'b111111111;
assign f[45][154] = 9'b111111111;
assign f[45][155] = 9'b111111111;
assign f[45][156] = 9'b111111111;
assign f[45][157] = 9'b111111111;
assign f[45][163] = 9'b111111111;
assign f[45][164] = 9'b111111111;
assign f[45][165] = 9'b111111111;
assign f[45][166] = 9'b111111111;
assign f[45][167] = 9'b111111111;
assign f[45][168] = 9'b111111111;
assign f[45][171] = 9'b111111111;
assign f[45][172] = 9'b111111111;
assign f[45][173] = 9'b111111111;
assign f[45][174] = 9'b111111111;
assign f[45][175] = 9'b111111111;
assign f[45][176] = 9'b111111111;
assign f[45][180] = 9'b111111111;
assign f[45][181] = 9'b111111111;
assign f[45][182] = 9'b111111111;
assign f[45][183] = 9'b111111111;
assign f[45][184] = 9'b111111111;
assign f[45][185] = 9'b111111111;
assign f[46][26] = 9'b111111111;
assign f[46][27] = 9'b111111111;
assign f[46][28] = 9'b111111111;
assign f[46][29] = 9'b111111111;
assign f[46][30] = 9'b111111111;
assign f[46][31] = 9'b111111111;
assign f[46][32] = 9'b111111111;
assign f[46][42] = 9'b111111111;
assign f[46][43] = 9'b111111111;
assign f[46][44] = 9'b111111111;
assign f[46][45] = 9'b111111111;
assign f[46][46] = 9'b111111111;
assign f[46][47] = 9'b111111111;
assign f[46][48] = 9'b111111111;
assign f[46][49] = 9'b111111111;
assign f[46][50] = 9'b111111111;
assign f[46][51] = 9'b111111111;
assign f[46][52] = 9'b111111111;
assign f[46][53] = 9'b111111111;
assign f[46][54] = 9'b111111111;
assign f[46][55] = 9'b111111111;
assign f[46][56] = 9'b111111111;
assign f[46][57] = 9'b111111111;
assign f[46][58] = 9'b111111111;
assign f[46][59] = 9'b111111111;
assign f[46][60] = 9'b111111111;
assign f[46][61] = 9'b111111111;
assign f[46][62] = 9'b111111111;
assign f[46][65] = 9'b111111111;
assign f[46][66] = 9'b111111111;
assign f[46][67] = 9'b111111111;
assign f[46][68] = 9'b111111111;
assign f[46][69] = 9'b111111111;
assign f[46][70] = 9'b111111111;
assign f[46][71] = 9'b111111111;
assign f[46][72] = 9'b111111111;
assign f[46][73] = 9'b111111111;
assign f[46][74] = 9'b111111111;
assign f[46][75] = 9'b111111111;
assign f[46][76] = 9'b111111111;
assign f[46][77] = 9'b111111111;
assign f[46][78] = 9'b111111111;
assign f[46][79] = 9'b111111111;
assign f[46][80] = 9'b111111111;
assign f[46][81] = 9'b111111111;
assign f[46][94] = 9'b111111111;
assign f[46][95] = 9'b111111111;
assign f[46][96] = 9'b111111111;
assign f[46][97] = 9'b111111111;
assign f[46][98] = 9'b111111111;
assign f[46][99] = 9'b111111111;
assign f[46][100] = 9'b111111111;
assign f[46][101] = 9'b111111111;
assign f[46][102] = 9'b111111111;
assign f[46][103] = 9'b111111111;
assign f[46][104] = 9'b111111111;
assign f[46][105] = 9'b111111111;
assign f[46][106] = 9'b111111111;
assign f[46][107] = 9'b111111111;
assign f[46][108] = 9'b111111111;
assign f[46][109] = 9'b111111111;
assign f[46][110] = 9'b111111111;
assign f[46][111] = 9'b111111111;
assign f[46][112] = 9'b111111111;
assign f[46][113] = 9'b111111111;
assign f[46][118] = 9'b111111111;
assign f[46][119] = 9'b111111111;
assign f[46][120] = 9'b111111111;
assign f[46][121] = 9'b111111111;
assign f[46][122] = 9'b111111111;
assign f[46][123] = 9'b111111111;
assign f[46][142] = 9'b111111111;
assign f[46][144] = 9'b111111111;
assign f[46][145] = 9'b111111111;
assign f[46][146] = 9'b111111111;
assign f[46][151] = 9'b111111111;
assign f[46][152] = 9'b111111111;
assign f[46][153] = 9'b111111111;
assign f[46][154] = 9'b111111111;
assign f[46][155] = 9'b111111111;
assign f[46][156] = 9'b111111111;
assign f[46][157] = 9'b111111111;
assign f[46][163] = 9'b111111111;
assign f[46][164] = 9'b111111111;
assign f[46][165] = 9'b111111111;
assign f[46][166] = 9'b111111111;
assign f[46][167] = 9'b111111111;
assign f[46][168] = 9'b111111111;
assign f[46][171] = 9'b111111111;
assign f[46][172] = 9'b111111111;
assign f[46][173] = 9'b111111111;
assign f[46][174] = 9'b111111111;
assign f[46][175] = 9'b111111111;
assign f[46][176] = 9'b111111111;
assign f[46][180] = 9'b111111111;
assign f[46][181] = 9'b111111111;
assign f[46][182] = 9'b111111111;
assign f[46][183] = 9'b111111111;
assign f[46][184] = 9'b111111111;
assign f[46][185] = 9'b111111111;
assign f[47][26] = 9'b111111111;
assign f[47][27] = 9'b111111111;
assign f[47][28] = 9'b111111111;
assign f[47][29] = 9'b111111111;
assign f[47][30] = 9'b111111111;
assign f[47][31] = 9'b111111111;
assign f[47][32] = 9'b111111111;
assign f[47][42] = 9'b111111111;
assign f[47][43] = 9'b111111111;
assign f[47][44] = 9'b111111111;
assign f[47][45] = 9'b111111111;
assign f[47][46] = 9'b111111111;
assign f[47][47] = 9'b111111111;
assign f[47][48] = 9'b111111111;
assign f[47][49] = 9'b111111111;
assign f[47][50] = 9'b111111111;
assign f[47][51] = 9'b111111111;
assign f[47][52] = 9'b111111111;
assign f[47][53] = 9'b111111111;
assign f[47][54] = 9'b111111111;
assign f[47][55] = 9'b111111111;
assign f[47][56] = 9'b111111111;
assign f[47][57] = 9'b111111111;
assign f[47][58] = 9'b111111111;
assign f[47][59] = 9'b111111111;
assign f[47][60] = 9'b111111111;
assign f[47][61] = 9'b111111111;
assign f[47][62] = 9'b111111111;
assign f[47][65] = 9'b111111111;
assign f[47][66] = 9'b111111111;
assign f[47][67] = 9'b111111111;
assign f[47][68] = 9'b111111111;
assign f[47][69] = 9'b111111111;
assign f[47][70] = 9'b111111111;
assign f[47][71] = 9'b111111111;
assign f[47][72] = 9'b111111111;
assign f[47][73] = 9'b111111111;
assign f[47][74] = 9'b111111111;
assign f[47][75] = 9'b111111111;
assign f[47][76] = 9'b111111111;
assign f[47][77] = 9'b111111111;
assign f[47][78] = 9'b111111111;
assign f[47][79] = 9'b111111111;
assign f[47][80] = 9'b111111111;
assign f[47][81] = 9'b111111111;
assign f[47][94] = 9'b111111111;
assign f[47][95] = 9'b111111111;
assign f[47][96] = 9'b111111111;
assign f[47][97] = 9'b111111111;
assign f[47][98] = 9'b111111111;
assign f[47][99] = 9'b111111111;
assign f[47][100] = 9'b111111111;
assign f[47][101] = 9'b111111111;
assign f[47][102] = 9'b111111111;
assign f[47][103] = 9'b111111111;
assign f[47][104] = 9'b111111111;
assign f[47][105] = 9'b111111111;
assign f[47][106] = 9'b111111111;
assign f[47][107] = 9'b111111111;
assign f[47][108] = 9'b111111111;
assign f[47][109] = 9'b111111111;
assign f[47][110] = 9'b111111111;
assign f[47][111] = 9'b111111111;
assign f[47][112] = 9'b111111111;
assign f[47][113] = 9'b111111111;
assign f[47][118] = 9'b111111111;
assign f[47][119] = 9'b111111111;
assign f[47][120] = 9'b111111111;
assign f[47][121] = 9'b111111111;
assign f[47][122] = 9'b111111111;
assign f[47][123] = 9'b111111111;
assign f[47][143] = 9'b111111111;
assign f[47][145] = 9'b111111111;
assign f[47][146] = 9'b111111111;
assign f[47][151] = 9'b111111111;
assign f[47][152] = 9'b111111111;
assign f[47][153] = 9'b111111111;
assign f[47][154] = 9'b111111111;
assign f[47][155] = 9'b111111111;
assign f[47][156] = 9'b111111111;
assign f[47][157] = 9'b111111111;
assign f[47][163] = 9'b111111111;
assign f[47][164] = 9'b111111111;
assign f[47][165] = 9'b111111111;
assign f[47][166] = 9'b111111111;
assign f[47][167] = 9'b111111111;
assign f[47][168] = 9'b111111111;
assign f[47][172] = 9'b111111111;
assign f[47][173] = 9'b111111111;
assign f[47][174] = 9'b111111111;
assign f[47][175] = 9'b111111111;
assign f[47][176] = 9'b111111111;
assign f[47][177] = 9'b111111111;
assign f[47][180] = 9'b111111111;
assign f[47][181] = 9'b111111111;
assign f[47][182] = 9'b111111111;
assign f[47][183] = 9'b111111111;
assign f[47][184] = 9'b111111111;
assign f[47][185] = 9'b111111111;
assign f[48][26] = 9'b111111111;
assign f[48][27] = 9'b111111111;
assign f[48][28] = 9'b111111111;
assign f[48][29] = 9'b111111111;
assign f[48][30] = 9'b111111111;
assign f[48][31] = 9'b111111111;
assign f[48][32] = 9'b111111111;
assign f[48][42] = 9'b111111111;
assign f[48][43] = 9'b111111111;
assign f[48][44] = 9'b111111111;
assign f[48][45] = 9'b111111111;
assign f[48][46] = 9'b111111111;
assign f[48][47] = 9'b111111111;
assign f[48][48] = 9'b111111111;
assign f[48][49] = 9'b111111111;
assign f[48][50] = 9'b111111111;
assign f[48][51] = 9'b111111111;
assign f[48][52] = 9'b111111111;
assign f[48][53] = 9'b111111111;
assign f[48][54] = 9'b111111111;
assign f[48][55] = 9'b111111111;
assign f[48][56] = 9'b111111111;
assign f[48][57] = 9'b111111111;
assign f[48][58] = 9'b111111111;
assign f[48][59] = 9'b111111111;
assign f[48][60] = 9'b111111111;
assign f[48][61] = 9'b111111111;
assign f[48][62] = 9'b111111111;
assign f[48][65] = 9'b111111111;
assign f[48][66] = 9'b111111111;
assign f[48][67] = 9'b111111111;
assign f[48][68] = 9'b111111111;
assign f[48][69] = 9'b111111111;
assign f[48][70] = 9'b111111111;
assign f[48][71] = 9'b111111111;
assign f[48][72] = 9'b111111111;
assign f[48][73] = 9'b111111111;
assign f[48][74] = 9'b111111111;
assign f[48][75] = 9'b111111111;
assign f[48][76] = 9'b111111111;
assign f[48][77] = 9'b111111111;
assign f[48][78] = 9'b111111111;
assign f[48][79] = 9'b111111111;
assign f[48][80] = 9'b111111111;
assign f[48][81] = 9'b111111111;
assign f[48][94] = 9'b111111111;
assign f[48][96] = 9'b111111111;
assign f[48][97] = 9'b111111111;
assign f[48][98] = 9'b111111111;
assign f[48][99] = 9'b111111111;
assign f[48][100] = 9'b111111111;
assign f[48][101] = 9'b111111111;
assign f[48][102] = 9'b111111111;
assign f[48][103] = 9'b111111111;
assign f[48][104] = 9'b111111111;
assign f[48][105] = 9'b111111111;
assign f[48][106] = 9'b111111111;
assign f[48][107] = 9'b111111111;
assign f[48][108] = 9'b111111111;
assign f[48][109] = 9'b111111111;
assign f[48][110] = 9'b111111111;
assign f[48][111] = 9'b111111111;
assign f[48][112] = 9'b111111111;
assign f[48][118] = 9'b111111111;
assign f[48][119] = 9'b111111111;
assign f[48][120] = 9'b111111111;
assign f[48][121] = 9'b111111111;
assign f[48][122] = 9'b111111111;
assign f[48][123] = 9'b111111111;
assign f[48][142] = 9'b111111111;
assign f[48][143] = 9'b111111111;
assign f[48][144] = 9'b111111111;
assign f[48][145] = 9'b111111111;
assign f[48][146] = 9'b111111111;
assign f[48][152] = 9'b111111111;
assign f[48][153] = 9'b111111111;
assign f[48][154] = 9'b111111111;
assign f[48][155] = 9'b111111111;
assign f[48][156] = 9'b111111111;
assign f[48][157] = 9'b111111111;
assign f[48][163] = 9'b111111111;
assign f[48][164] = 9'b111111111;
assign f[48][165] = 9'b111111111;
assign f[48][166] = 9'b111111111;
assign f[48][167] = 9'b111111111;
assign f[48][168] = 9'b111111111;
assign f[48][172] = 9'b111111111;
assign f[48][173] = 9'b111111111;
assign f[48][174] = 9'b111111111;
assign f[48][175] = 9'b111111111;
assign f[48][176] = 9'b111111111;
assign f[48][177] = 9'b111111111;
assign f[48][180] = 9'b111111111;
assign f[48][181] = 9'b111111111;
assign f[48][184] = 9'b111111111;
assign f[48][185] = 9'b111111111;
assign f[49][26] = 9'b111111111;
assign f[49][27] = 9'b111111111;
assign f[49][28] = 9'b111111111;
assign f[49][29] = 9'b111111111;
assign f[49][30] = 9'b111111111;
assign f[49][31] = 9'b111111111;
assign f[49][32] = 9'b111111111;
assign f[49][42] = 9'b111111111;
assign f[49][43] = 9'b111111111;
assign f[49][44] = 9'b111111111;
assign f[49][45] = 9'b111111111;
assign f[49][46] = 9'b111111111;
assign f[49][47] = 9'b111111111;
assign f[49][50] = 9'b111111111;
assign f[49][51] = 9'b111111111;
assign f[49][52] = 9'b111111111;
assign f[49][53] = 9'b111111111;
assign f[49][54] = 9'b111111111;
assign f[49][55] = 9'b111111111;
assign f[49][56] = 9'b111111111;
assign f[49][57] = 9'b111111111;
assign f[49][58] = 9'b111111111;
assign f[49][59] = 9'b111111111;
assign f[49][60] = 9'b111111111;
assign f[49][61] = 9'b111111111;
assign f[49][62] = 9'b111111111;
assign f[49][65] = 9'b111111111;
assign f[49][66] = 9'b111111111;
assign f[49][67] = 9'b111111111;
assign f[49][68] = 9'b111111111;
assign f[49][69] = 9'b111111111;
assign f[49][70] = 9'b111111111;
assign f[49][71] = 9'b111111111;
assign f[49][72] = 9'b111111111;
assign f[49][73] = 9'b111111111;
assign f[49][74] = 9'b111111111;
assign f[49][75] = 9'b111111111;
assign f[49][76] = 9'b111111111;
assign f[49][77] = 9'b111111111;
assign f[49][78] = 9'b111111111;
assign f[49][79] = 9'b111111111;
assign f[49][80] = 9'b111111111;
assign f[49][81] = 9'b111111111;
assign f[49][94] = 9'b111111111;
assign f[49][95] = 9'b111111111;
assign f[49][96] = 9'b111111111;
assign f[49][97] = 9'b111111111;
assign f[49][98] = 9'b111111111;
assign f[49][99] = 9'b111111111;
assign f[49][100] = 9'b111111111;
assign f[49][101] = 9'b111111111;
assign f[49][102] = 9'b111111111;
assign f[49][103] = 9'b111111111;
assign f[49][104] = 9'b111111111;
assign f[49][105] = 9'b111111111;
assign f[49][106] = 9'b111111111;
assign f[49][107] = 9'b111111111;
assign f[49][108] = 9'b111111111;
assign f[49][109] = 9'b111111111;
assign f[49][110] = 9'b111111111;
assign f[49][111] = 9'b111111111;
assign f[49][117] = 9'b111111111;
assign f[49][118] = 9'b111111111;
assign f[49][119] = 9'b111111111;
assign f[49][120] = 9'b111111111;
assign f[49][121] = 9'b111111111;
assign f[49][122] = 9'b111111111;
assign f[49][123] = 9'b111111111;
assign f[49][141] = 9'b111111111;
assign f[49][142] = 9'b111111111;
assign f[49][143] = 9'b111111111;
assign f[49][144] = 9'b111111111;
assign f[49][145] = 9'b111111111;
assign f[49][146] = 9'b111111111;
assign f[49][152] = 9'b111111111;
assign f[49][153] = 9'b111111111;
assign f[49][154] = 9'b111111111;
assign f[49][155] = 9'b111111111;
assign f[49][156] = 9'b111111111;
assign f[49][157] = 9'b111111111;
assign f[49][158] = 9'b111111111;
assign f[49][163] = 9'b111111111;
assign f[49][164] = 9'b111111111;
assign f[49][165] = 9'b111111111;
assign f[49][166] = 9'b111111111;
assign f[49][167] = 9'b111111111;
assign f[49][168] = 9'b111111111;
assign f[49][169] = 9'b111111111;
assign f[49][172] = 9'b111111111;
assign f[49][173] = 9'b111111111;
assign f[49][174] = 9'b111111111;
assign f[49][175] = 9'b111111111;
assign f[49][176] = 9'b111111111;
assign f[49][177] = 9'b111111111;
assign f[49][180] = 9'b111111111;
assign f[49][181] = 9'b111111111;
assign f[49][182] = 9'b111111111;
assign f[49][183] = 9'b111111111;
assign f[49][184] = 9'b111111111;
assign f[49][185] = 9'b111111111;
assign f[50][26] = 9'b111111111;
assign f[50][27] = 9'b111111111;
assign f[50][28] = 9'b111111111;
assign f[50][29] = 9'b111111111;
assign f[50][30] = 9'b111111111;
assign f[50][31] = 9'b111111111;
assign f[50][32] = 9'b111111111;
assign f[50][42] = 9'b111111111;
assign f[50][43] = 9'b111111111;
assign f[50][44] = 9'b111111111;
assign f[50][45] = 9'b111111111;
assign f[50][46] = 9'b111111111;
assign f[50][47] = 9'b111111111;
assign f[50][48] = 9'b111111111;
assign f[50][55] = 9'b111111111;
assign f[50][56] = 9'b111111111;
assign f[50][57] = 9'b111111111;
assign f[50][58] = 9'b111111111;
assign f[50][59] = 9'b111111111;
assign f[50][60] = 9'b111111111;
assign f[50][61] = 9'b111111111;
assign f[50][62] = 9'b111111111;
assign f[50][65] = 9'b111111111;
assign f[50][66] = 9'b111111111;
assign f[50][67] = 9'b111111111;
assign f[50][68] = 9'b111111111;
assign f[50][69] = 9'b111111111;
assign f[50][70] = 9'b111111111;
assign f[50][71] = 9'b111111111;
assign f[50][72] = 9'b111111111;
assign f[50][73] = 9'b111111111;
assign f[50][74] = 9'b111111111;
assign f[50][75] = 9'b111111111;
assign f[50][76] = 9'b111111111;
assign f[50][77] = 9'b111111111;
assign f[50][78] = 9'b111111111;
assign f[50][79] = 9'b111111111;
assign f[50][80] = 9'b111111111;
assign f[50][94] = 9'b111111111;
assign f[50][95] = 9'b111111111;
assign f[50][96] = 9'b111111111;
assign f[50][97] = 9'b111111111;
assign f[50][98] = 9'b111111111;
assign f[50][99] = 9'b111111111;
assign f[50][100] = 9'b111111111;
assign f[50][101] = 9'b111111111;
assign f[50][102] = 9'b111111111;
assign f[50][103] = 9'b111111111;
assign f[50][104] = 9'b111111111;
assign f[50][105] = 9'b111111111;
assign f[50][106] = 9'b111111111;
assign f[50][107] = 9'b111111111;
assign f[50][108] = 9'b111111111;
assign f[50][109] = 9'b111111111;
assign f[50][110] = 9'b111111111;
assign f[50][117] = 9'b111111111;
assign f[50][118] = 9'b111111111;
assign f[50][119] = 9'b111111111;
assign f[50][120] = 9'b111111111;
assign f[50][121] = 9'b111111111;
assign f[50][122] = 9'b111111111;
assign f[50][123] = 9'b111111111;
assign f[50][141] = 9'b111111111;
assign f[50][142] = 9'b111111111;
assign f[50][143] = 9'b111111111;
assign f[50][144] = 9'b111111111;
assign f[50][145] = 9'b111111111;
assign f[50][152] = 9'b111111111;
assign f[50][153] = 9'b111111111;
assign f[50][154] = 9'b111111111;
assign f[50][155] = 9'b111111111;
assign f[50][156] = 9'b111111111;
assign f[50][157] = 9'b111111111;
assign f[50][158] = 9'b111111111;
assign f[50][164] = 9'b111111111;
assign f[50][165] = 9'b111111111;
assign f[50][166] = 9'b111111111;
assign f[50][167] = 9'b111111111;
assign f[50][168] = 9'b111111111;
assign f[50][169] = 9'b111111111;
assign f[50][172] = 9'b111111111;
assign f[50][173] = 9'b111111111;
assign f[50][174] = 9'b111111111;
assign f[50][176] = 9'b111111111;
assign f[50][177] = 9'b111111111;
assign f[50][180] = 9'b111111111;
assign f[50][181] = 9'b111111111;
assign f[50][182] = 9'b111111111;
assign f[50][183] = 9'b111111111;
assign f[50][184] = 9'b111111111;
assign f[50][185] = 9'b111111111;
assign f[51][26] = 9'b111111111;
assign f[51][27] = 9'b111111111;
assign f[51][28] = 9'b111111111;
assign f[51][29] = 9'b111111111;
assign f[51][30] = 9'b111111111;
assign f[51][31] = 9'b111111111;
assign f[51][32] = 9'b111111111;
assign f[51][42] = 9'b111111111;
assign f[51][43] = 9'b111111111;
assign f[51][44] = 9'b111111111;
assign f[51][45] = 9'b111111111;
assign f[51][46] = 9'b111111111;
assign f[51][47] = 9'b111111111;
assign f[51][48] = 9'b111111111;
assign f[51][56] = 9'b111111111;
assign f[51][57] = 9'b111111111;
assign f[51][58] = 9'b111111111;
assign f[51][59] = 9'b111111111;
assign f[51][60] = 9'b111111111;
assign f[51][61] = 9'b111111111;
assign f[51][62] = 9'b111111111;
assign f[51][65] = 9'b111111111;
assign f[51][66] = 9'b111111111;
assign f[51][67] = 9'b111111111;
assign f[51][68] = 9'b111111111;
assign f[51][69] = 9'b111111111;
assign f[51][70] = 9'b111111111;
assign f[51][71] = 9'b111111111;
assign f[51][94] = 9'b111111111;
assign f[51][95] = 9'b111111111;
assign f[51][96] = 9'b111111111;
assign f[51][97] = 9'b111111111;
assign f[51][98] = 9'b111111111;
assign f[51][99] = 9'b111111111;
assign f[51][100] = 9'b111111111;
assign f[51][101] = 9'b111111111;
assign f[51][102] = 9'b111111111;
assign f[51][103] = 9'b111111111;
assign f[51][104] = 9'b111111111;
assign f[51][105] = 9'b111111111;
assign f[51][106] = 9'b111111111;
assign f[51][107] = 9'b111111111;
assign f[51][108] = 9'b111111111;
assign f[51][109] = 9'b111111111;
assign f[51][117] = 9'b111111111;
assign f[51][118] = 9'b111111111;
assign f[51][119] = 9'b111111111;
assign f[51][120] = 9'b111111111;
assign f[51][121] = 9'b111111111;
assign f[51][122] = 9'b111111111;
assign f[51][123] = 9'b111111111;
assign f[51][142] = 9'b111111111;
assign f[51][143] = 9'b111111111;
assign f[51][144] = 9'b111111111;
assign f[51][145] = 9'b111111111;
assign f[51][152] = 9'b111111111;
assign f[51][153] = 9'b111111111;
assign f[51][154] = 9'b111111111;
assign f[51][155] = 9'b111111111;
assign f[51][156] = 9'b111111111;
assign f[51][157] = 9'b111111111;
assign f[51][158] = 9'b111111111;
assign f[51][163] = 9'b111111111;
assign f[51][164] = 9'b111111111;
assign f[51][165] = 9'b111111111;
assign f[51][166] = 9'b111111111;
assign f[51][167] = 9'b111111111;
assign f[51][168] = 9'b111111111;
assign f[51][173] = 9'b111111111;
assign f[51][176] = 9'b111111111;
assign f[51][177] = 9'b111111111;
assign f[51][180] = 9'b111111111;
assign f[51][181] = 9'b111111111;
assign f[51][182] = 9'b111111111;
assign f[51][183] = 9'b111111111;
assign f[51][184] = 9'b111111111;
assign f[51][185] = 9'b111111111;
assign f[52][26] = 9'b111111111;
assign f[52][27] = 9'b111111111;
assign f[52][28] = 9'b111111111;
assign f[52][29] = 9'b111111111;
assign f[52][30] = 9'b111111111;
assign f[52][31] = 9'b111111111;
assign f[52][32] = 9'b111111111;
assign f[52][42] = 9'b111111111;
assign f[52][43] = 9'b111111111;
assign f[52][44] = 9'b111111111;
assign f[52][45] = 9'b111111111;
assign f[52][46] = 9'b111111111;
assign f[52][47] = 9'b111111111;
assign f[52][48] = 9'b111111111;
assign f[52][56] = 9'b111111111;
assign f[52][57] = 9'b111111111;
assign f[52][58] = 9'b111111111;
assign f[52][59] = 9'b111111111;
assign f[52][60] = 9'b111111111;
assign f[52][61] = 9'b111111111;
assign f[52][62] = 9'b111111111;
assign f[52][65] = 9'b111111111;
assign f[52][66] = 9'b111111111;
assign f[52][67] = 9'b111111111;
assign f[52][68] = 9'b111111111;
assign f[52][69] = 9'b111111111;
assign f[52][70] = 9'b111111111;
assign f[52][71] = 9'b111111111;
assign f[52][95] = 9'b111111111;
assign f[52][96] = 9'b111111111;
assign f[52][97] = 9'b111111111;
assign f[52][98] = 9'b111111111;
assign f[52][99] = 9'b111111111;
assign f[52][100] = 9'b111111111;
assign f[52][117] = 9'b111111111;
assign f[52][118] = 9'b111111111;
assign f[52][120] = 9'b111111111;
assign f[52][121] = 9'b111111111;
assign f[52][122] = 9'b111111111;
assign f[52][123] = 9'b111111111;
assign f[52][140] = 9'b111111111;
assign f[52][141] = 9'b111111111;
assign f[52][142] = 9'b111111111;
assign f[52][143] = 9'b111111111;
assign f[52][144] = 9'b111111111;
assign f[52][145] = 9'b111111111;
assign f[52][149] = 9'b111111111;
assign f[52][151] = 9'b111111111;
assign f[52][152] = 9'b111111111;
assign f[52][153] = 9'b111111111;
assign f[52][154] = 9'b111111111;
assign f[52][155] = 9'b111111111;
assign f[52][156] = 9'b111111111;
assign f[52][157] = 9'b111111111;
assign f[52][158] = 9'b111111111;
assign f[52][163] = 9'b111111111;
assign f[52][164] = 9'b111111111;
assign f[52][165] = 9'b111111111;
assign f[52][166] = 9'b111111111;
assign f[52][167] = 9'b111111111;
assign f[52][168] = 9'b111111111;
assign f[52][172] = 9'b111111111;
assign f[52][173] = 9'b111111111;
assign f[52][176] = 9'b111111111;
assign f[52][177] = 9'b111111111;
assign f[52][178] = 9'b111111111;
assign f[52][180] = 9'b111111111;
assign f[52][181] = 9'b111111111;
assign f[52][182] = 9'b111111111;
assign f[52][183] = 9'b111111111;
assign f[52][184] = 9'b111111111;
assign f[52][185] = 9'b111111111;
assign f[53][26] = 9'b111111111;
assign f[53][27] = 9'b111111111;
assign f[53][28] = 9'b111111111;
assign f[53][29] = 9'b111111111;
assign f[53][30] = 9'b111111111;
assign f[53][31] = 9'b111111111;
assign f[53][32] = 9'b111111111;
assign f[53][33] = 9'b111111111;
assign f[53][42] = 9'b111111111;
assign f[53][43] = 9'b111111111;
assign f[53][44] = 9'b111111111;
assign f[53][45] = 9'b111111111;
assign f[53][46] = 9'b111111111;
assign f[53][47] = 9'b111111111;
assign f[53][48] = 9'b111111111;
assign f[53][56] = 9'b111111111;
assign f[53][57] = 9'b111111111;
assign f[53][58] = 9'b111111111;
assign f[53][59] = 9'b111111111;
assign f[53][60] = 9'b111111111;
assign f[53][61] = 9'b111111111;
assign f[53][62] = 9'b111111111;
assign f[53][65] = 9'b111111111;
assign f[53][66] = 9'b111111111;
assign f[53][67] = 9'b111111111;
assign f[53][68] = 9'b111111111;
assign f[53][69] = 9'b111111111;
assign f[53][70] = 9'b111111111;
assign f[53][71] = 9'b111111111;
assign f[53][94] = 9'b111111111;
assign f[53][95] = 9'b111111111;
assign f[53][96] = 9'b111111111;
assign f[53][97] = 9'b111111111;
assign f[53][98] = 9'b111111111;
assign f[53][99] = 9'b111111111;
assign f[53][100] = 9'b111111111;
assign f[53][117] = 9'b111111111;
assign f[53][118] = 9'b111111111;
assign f[53][121] = 9'b111111111;
assign f[53][122] = 9'b111111111;
assign f[53][123] = 9'b111111111;
assign f[53][140] = 9'b111111111;
assign f[53][141] = 9'b111111111;
assign f[53][142] = 9'b111111111;
assign f[53][143] = 9'b111111111;
assign f[53][144] = 9'b111111111;
assign f[53][145] = 9'b111111111;
assign f[53][146] = 9'b111111111;
assign f[53][147] = 9'b111111111;
assign f[53][148] = 9'b111111111;
assign f[53][149] = 9'b111111111;
assign f[53][150] = 9'b111111111;
assign f[53][151] = 9'b111111111;
assign f[53][152] = 9'b111111111;
assign f[53][153] = 9'b111111111;
assign f[53][154] = 9'b111111111;
assign f[53][155] = 9'b111111111;
assign f[53][156] = 9'b111111111;
assign f[53][157] = 9'b111111111;
assign f[53][158] = 9'b111111111;
assign f[53][163] = 9'b111111111;
assign f[53][164] = 9'b111111111;
assign f[53][165] = 9'b111111111;
assign f[53][166] = 9'b111111111;
assign f[53][167] = 9'b111111111;
assign f[53][168] = 9'b111111111;
assign f[53][173] = 9'b111111111;
assign f[53][174] = 9'b111111111;
assign f[53][175] = 9'b111111111;
assign f[53][176] = 9'b111111111;
assign f[53][177] = 9'b111111111;
assign f[53][178] = 9'b111111111;
assign f[53][180] = 9'b111111111;
assign f[53][181] = 9'b111111111;
assign f[53][182] = 9'b111111111;
assign f[53][183] = 9'b111111111;
assign f[53][184] = 9'b111111111;
assign f[53][185] = 9'b111111111;
assign f[54][26] = 9'b111111111;
assign f[54][27] = 9'b111111111;
assign f[54][28] = 9'b111111111;
assign f[54][29] = 9'b111111111;
assign f[54][30] = 9'b111111111;
assign f[54][31] = 9'b111111111;
assign f[54][32] = 9'b111111111;
assign f[54][42] = 9'b111111111;
assign f[54][43] = 9'b111111111;
assign f[54][44] = 9'b111111111;
assign f[54][45] = 9'b111111111;
assign f[54][46] = 9'b111111111;
assign f[54][47] = 9'b111111111;
assign f[54][48] = 9'b111111111;
assign f[54][56] = 9'b111111111;
assign f[54][57] = 9'b111111111;
assign f[54][58] = 9'b111111111;
assign f[54][59] = 9'b111111111;
assign f[54][60] = 9'b111111111;
assign f[54][61] = 9'b111111111;
assign f[54][62] = 9'b111111111;
assign f[54][65] = 9'b111111111;
assign f[54][66] = 9'b111111111;
assign f[54][67] = 9'b111111111;
assign f[54][68] = 9'b111111111;
assign f[54][69] = 9'b111111111;
assign f[54][70] = 9'b111111111;
assign f[54][71] = 9'b111111111;
assign f[54][72] = 9'b111111111;
assign f[54][94] = 9'b111111111;
assign f[54][95] = 9'b111111111;
assign f[54][96] = 9'b111111111;
assign f[54][97] = 9'b111111111;
assign f[54][98] = 9'b111111111;
assign f[54][99] = 9'b111111111;
assign f[54][100] = 9'b111111111;
assign f[54][117] = 9'b111111111;
assign f[54][118] = 9'b111111111;
assign f[54][119] = 9'b111111111;
assign f[54][120] = 9'b111111111;
assign f[54][121] = 9'b111111111;
assign f[54][122] = 9'b111111111;
assign f[54][123] = 9'b111111111;
assign f[54][139] = 9'b111111111;
assign f[54][140] = 9'b111111111;
assign f[54][141] = 9'b111111111;
assign f[54][142] = 9'b111111111;
assign f[54][143] = 9'b111111111;
assign f[54][144] = 9'b111111111;
assign f[54][145] = 9'b111111111;
assign f[54][146] = 9'b111111111;
assign f[54][147] = 9'b111111111;
assign f[54][148] = 9'b111111111;
assign f[54][149] = 9'b111111111;
assign f[54][150] = 9'b111111111;
assign f[54][151] = 9'b111111111;
assign f[54][152] = 9'b111111111;
assign f[54][153] = 9'b111111111;
assign f[54][154] = 9'b111111111;
assign f[54][155] = 9'b111111111;
assign f[54][156] = 9'b111111111;
assign f[54][157] = 9'b111111111;
assign f[54][158] = 9'b111111111;
assign f[54][159] = 9'b111111111;
assign f[54][163] = 9'b111111111;
assign f[54][164] = 9'b111111111;
assign f[54][165] = 9'b111111111;
assign f[54][166] = 9'b111111111;
assign f[54][167] = 9'b111111111;
assign f[54][168] = 9'b111111111;
assign f[54][169] = 9'b111111111;
assign f[54][173] = 9'b111111111;
assign f[54][174] = 9'b111111111;
assign f[54][175] = 9'b111111111;
assign f[54][176] = 9'b111111111;
assign f[54][177] = 9'b111111111;
assign f[54][178] = 9'b111111111;
assign f[54][180] = 9'b111111111;
assign f[54][181] = 9'b111111111;
assign f[54][182] = 9'b111111111;
assign f[54][183] = 9'b111111111;
assign f[54][184] = 9'b111111111;
assign f[54][185] = 9'b111111111;
assign f[55][26] = 9'b111111111;
assign f[55][27] = 9'b111111111;
assign f[55][28] = 9'b111111111;
assign f[55][29] = 9'b111111111;
assign f[55][30] = 9'b111111111;
assign f[55][31] = 9'b111111111;
assign f[55][32] = 9'b111111111;
assign f[55][42] = 9'b111111111;
assign f[55][43] = 9'b111111111;
assign f[55][44] = 9'b111111111;
assign f[55][45] = 9'b111111111;
assign f[55][46] = 9'b111111111;
assign f[55][47] = 9'b111111111;
assign f[55][48] = 9'b111111111;
assign f[55][56] = 9'b111111111;
assign f[55][57] = 9'b111111111;
assign f[55][58] = 9'b111111111;
assign f[55][59] = 9'b111111111;
assign f[55][60] = 9'b111111111;
assign f[55][61] = 9'b111111111;
assign f[55][62] = 9'b111111111;
assign f[55][65] = 9'b111111111;
assign f[55][66] = 9'b111111111;
assign f[55][67] = 9'b111111111;
assign f[55][68] = 9'b111111111;
assign f[55][69] = 9'b111111111;
assign f[55][70] = 9'b111111111;
assign f[55][71] = 9'b111111111;
assign f[55][94] = 9'b111111111;
assign f[55][95] = 9'b111111111;
assign f[55][96] = 9'b111111111;
assign f[55][97] = 9'b111111111;
assign f[55][98] = 9'b111111111;
assign f[55][99] = 9'b111111111;
assign f[55][100] = 9'b111111111;
assign f[55][117] = 9'b111111111;
assign f[55][118] = 9'b111111111;
assign f[55][120] = 9'b111111111;
assign f[55][121] = 9'b111111111;
assign f[55][122] = 9'b111111111;
assign f[55][123] = 9'b111111111;
assign f[55][139] = 9'b111111111;
assign f[55][140] = 9'b111111111;
assign f[55][141] = 9'b111111111;
assign f[55][142] = 9'b111111111;
assign f[55][143] = 9'b111111111;
assign f[55][144] = 9'b111111111;
assign f[55][145] = 9'b111111111;
assign f[55][146] = 9'b111111111;
assign f[55][147] = 9'b111111111;
assign f[55][148] = 9'b111111111;
assign f[55][149] = 9'b111111111;
assign f[55][150] = 9'b111111111;
assign f[55][151] = 9'b111111111;
assign f[55][152] = 9'b111111111;
assign f[55][153] = 9'b111111111;
assign f[55][154] = 9'b111111111;
assign f[55][155] = 9'b111111111;
assign f[55][156] = 9'b111111111;
assign f[55][157] = 9'b111111111;
assign f[55][158] = 9'b111111111;
assign f[55][159] = 9'b111111111;
assign f[55][163] = 9'b111111111;
assign f[55][164] = 9'b111111111;
assign f[55][165] = 9'b111111111;
assign f[55][166] = 9'b111111111;
assign f[55][167] = 9'b111111111;
assign f[55][168] = 9'b111111111;
assign f[55][169] = 9'b111111111;
assign f[55][173] = 9'b111111111;
assign f[55][174] = 9'b111111111;
assign f[55][175] = 9'b111111111;
assign f[55][176] = 9'b111111111;
assign f[55][177] = 9'b111111111;
assign f[55][178] = 9'b111111111;
assign f[55][179] = 9'b111111111;
assign f[55][180] = 9'b111111111;
assign f[55][181] = 9'b111111111;
assign f[55][182] = 9'b111111111;
assign f[55][183] = 9'b111111111;
assign f[55][184] = 9'b111111111;
assign f[55][185] = 9'b111111111;
assign f[56][26] = 9'b111111111;
assign f[56][27] = 9'b111111111;
assign f[56][28] = 9'b111111111;
assign f[56][29] = 9'b111111111;
assign f[56][30] = 9'b111111111;
assign f[56][31] = 9'b111111111;
assign f[56][32] = 9'b111111111;
assign f[56][42] = 9'b111111111;
assign f[56][43] = 9'b111111111;
assign f[56][44] = 9'b111111111;
assign f[56][45] = 9'b111111111;
assign f[56][46] = 9'b111111111;
assign f[56][47] = 9'b111111111;
assign f[56][48] = 9'b111111111;
assign f[56][56] = 9'b111111111;
assign f[56][57] = 9'b111111111;
assign f[56][58] = 9'b111111111;
assign f[56][59] = 9'b111111111;
assign f[56][60] = 9'b111111111;
assign f[56][61] = 9'b111111111;
assign f[56][62] = 9'b111111111;
assign f[56][65] = 9'b111111111;
assign f[56][66] = 9'b111111111;
assign f[56][67] = 9'b111111111;
assign f[56][68] = 9'b111111111;
assign f[56][69] = 9'b111111111;
assign f[56][70] = 9'b111111111;
assign f[56][71] = 9'b111111111;
assign f[56][94] = 9'b111111111;
assign f[56][95] = 9'b111111111;
assign f[56][96] = 9'b111111111;
assign f[56][97] = 9'b111111111;
assign f[56][98] = 9'b111111111;
assign f[56][99] = 9'b111111111;
assign f[56][100] = 9'b111111111;
assign f[56][117] = 9'b111111111;
assign f[56][118] = 9'b111111111;
assign f[56][119] = 9'b111111111;
assign f[56][120] = 9'b111111111;
assign f[56][121] = 9'b111111111;
assign f[56][122] = 9'b111111111;
assign f[56][123] = 9'b111111111;
assign f[56][139] = 9'b111111111;
assign f[56][140] = 9'b111111111;
assign f[56][141] = 9'b111111111;
assign f[56][142] = 9'b111111111;
assign f[56][143] = 9'b111111111;
assign f[56][144] = 9'b111111111;
assign f[56][145] = 9'b111111111;
assign f[56][146] = 9'b111111111;
assign f[56][147] = 9'b111111111;
assign f[56][148] = 9'b111111111;
assign f[56][149] = 9'b111111111;
assign f[56][150] = 9'b111111111;
assign f[56][151] = 9'b111111111;
assign f[56][152] = 9'b111111111;
assign f[56][153] = 9'b111111111;
assign f[56][154] = 9'b111111111;
assign f[56][155] = 9'b111111111;
assign f[56][156] = 9'b111111111;
assign f[56][157] = 9'b111111111;
assign f[56][158] = 9'b111111111;
assign f[56][159] = 9'b111111111;
assign f[56][163] = 9'b111111111;
assign f[56][164] = 9'b111111111;
assign f[56][165] = 9'b111111111;
assign f[56][166] = 9'b111111111;
assign f[56][167] = 9'b111111111;
assign f[56][168] = 9'b111111111;
assign f[56][169] = 9'b111111111;
assign f[56][174] = 9'b111111111;
assign f[56][175] = 9'b111111111;
assign f[56][176] = 9'b111111111;
assign f[56][177] = 9'b111111111;
assign f[56][178] = 9'b111111111;
assign f[56][179] = 9'b111111111;
assign f[56][180] = 9'b111111111;
assign f[56][181] = 9'b111111111;
assign f[56][183] = 9'b111111111;
assign f[56][184] = 9'b111111111;
assign f[56][185] = 9'b111111111;
assign f[57][26] = 9'b111111111;
assign f[57][27] = 9'b111111111;
assign f[57][28] = 9'b111111111;
assign f[57][29] = 9'b111111111;
assign f[57][30] = 9'b111111111;
assign f[57][31] = 9'b111111111;
assign f[57][32] = 9'b111111111;
assign f[57][33] = 9'b111111111;
assign f[57][42] = 9'b111111111;
assign f[57][43] = 9'b111111111;
assign f[57][44] = 9'b111111111;
assign f[57][45] = 9'b111111111;
assign f[57][46] = 9'b111111111;
assign f[57][47] = 9'b111111111;
assign f[57][48] = 9'b111111111;
assign f[57][56] = 9'b111111111;
assign f[57][57] = 9'b111111111;
assign f[57][58] = 9'b111111111;
assign f[57][59] = 9'b111111111;
assign f[57][60] = 9'b111111111;
assign f[57][61] = 9'b111111111;
assign f[57][62] = 9'b111111111;
assign f[57][65] = 9'b111111111;
assign f[57][66] = 9'b111111111;
assign f[57][67] = 9'b111111111;
assign f[57][68] = 9'b111111111;
assign f[57][69] = 9'b111111111;
assign f[57][70] = 9'b111111111;
assign f[57][71] = 9'b111111111;
assign f[57][94] = 9'b111111111;
assign f[57][95] = 9'b111111111;
assign f[57][96] = 9'b111111111;
assign f[57][97] = 9'b111111111;
assign f[57][98] = 9'b111111111;
assign f[57][99] = 9'b111111111;
assign f[57][100] = 9'b111111111;
assign f[57][117] = 9'b111111111;
assign f[57][118] = 9'b111111111;
assign f[57][119] = 9'b111111111;
assign f[57][120] = 9'b111111111;
assign f[57][121] = 9'b111111111;
assign f[57][122] = 9'b111111111;
assign f[57][123] = 9'b111111111;
assign f[57][138] = 9'b111111111;
assign f[57][139] = 9'b111111111;
assign f[57][140] = 9'b111111111;
assign f[57][141] = 9'b111111111;
assign f[57][142] = 9'b111111111;
assign f[57][143] = 9'b111111111;
assign f[57][144] = 9'b111111111;
assign f[57][145] = 9'b111111111;
assign f[57][146] = 9'b111111111;
assign f[57][147] = 9'b111111111;
assign f[57][148] = 9'b111111111;
assign f[57][149] = 9'b111111111;
assign f[57][150] = 9'b111111111;
assign f[57][151] = 9'b111111111;
assign f[57][152] = 9'b111111111;
assign f[57][153] = 9'b111111111;
assign f[57][154] = 9'b111111111;
assign f[57][155] = 9'b111111111;
assign f[57][156] = 9'b111111111;
assign f[57][157] = 9'b111111111;
assign f[57][158] = 9'b111111111;
assign f[57][159] = 9'b111111111;
assign f[57][163] = 9'b111111111;
assign f[57][164] = 9'b111111111;
assign f[57][165] = 9'b111111111;
assign f[57][166] = 9'b111111111;
assign f[57][167] = 9'b111111111;
assign f[57][168] = 9'b111111111;
assign f[57][169] = 9'b111111111;
assign f[57][174] = 9'b111111111;
assign f[57][175] = 9'b111111111;
assign f[57][176] = 9'b111111111;
assign f[57][177] = 9'b111111111;
assign f[57][178] = 9'b111111111;
assign f[57][179] = 9'b111111111;
assign f[57][180] = 9'b111111111;
assign f[57][181] = 9'b111111111;
assign f[57][182] = 9'b111111111;
assign f[57][183] = 9'b111111111;
assign f[57][184] = 9'b111111111;
assign f[57][185] = 9'b111111111;
assign f[58][26] = 9'b111111111;
assign f[58][27] = 9'b111111111;
assign f[58][28] = 9'b111111111;
assign f[58][29] = 9'b111111111;
assign f[58][30] = 9'b111111111;
assign f[58][31] = 9'b111111111;
assign f[58][32] = 9'b111111111;
assign f[58][33] = 9'b111111111;
assign f[58][42] = 9'b111111111;
assign f[58][43] = 9'b111111111;
assign f[58][44] = 9'b111111111;
assign f[58][45] = 9'b111111111;
assign f[58][46] = 9'b111111111;
assign f[58][47] = 9'b111111111;
assign f[58][48] = 9'b111111111;
assign f[58][56] = 9'b111111111;
assign f[58][57] = 9'b111111111;
assign f[58][58] = 9'b111111111;
assign f[58][59] = 9'b111111111;
assign f[58][60] = 9'b111111111;
assign f[58][61] = 9'b111111111;
assign f[58][62] = 9'b111111111;
assign f[58][65] = 9'b111111111;
assign f[58][66] = 9'b111111111;
assign f[58][67] = 9'b111111111;
assign f[58][68] = 9'b111111111;
assign f[58][69] = 9'b111111111;
assign f[58][70] = 9'b111111111;
assign f[58][71] = 9'b111111111;
assign f[58][94] = 9'b111111111;
assign f[58][95] = 9'b111111111;
assign f[58][96] = 9'b111111111;
assign f[58][97] = 9'b111111111;
assign f[58][98] = 9'b111111111;
assign f[58][99] = 9'b111111111;
assign f[58][100] = 9'b111111111;
assign f[58][117] = 9'b111111111;
assign f[58][118] = 9'b111111111;
assign f[58][119] = 9'b111111111;
assign f[58][120] = 9'b111111111;
assign f[58][121] = 9'b111111111;
assign f[58][122] = 9'b111111111;
assign f[58][123] = 9'b111111111;
assign f[58][138] = 9'b111111111;
assign f[58][139] = 9'b111111111;
assign f[58][140] = 9'b111111111;
assign f[58][141] = 9'b111111111;
assign f[58][142] = 9'b111111111;
assign f[58][143] = 9'b111111111;
assign f[58][153] = 9'b111111111;
assign f[58][154] = 9'b111111111;
assign f[58][155] = 9'b111111111;
assign f[58][156] = 9'b111111111;
assign f[58][157] = 9'b111111111;
assign f[58][158] = 9'b111111111;
assign f[58][159] = 9'b111111111;
assign f[58][160] = 9'b111111111;
assign f[58][163] = 9'b111111111;
assign f[58][164] = 9'b111111111;
assign f[58][165] = 9'b111111111;
assign f[58][166] = 9'b111111111;
assign f[58][167] = 9'b111111111;
assign f[58][168] = 9'b111111111;
assign f[58][169] = 9'b111111111;
assign f[58][174] = 9'b111111111;
assign f[58][175] = 9'b111111111;
assign f[58][176] = 9'b111111111;
assign f[58][177] = 9'b111111111;
assign f[58][178] = 9'b111111111;
assign f[58][179] = 9'b111111111;
assign f[58][180] = 9'b111111111;
assign f[58][181] = 9'b111111111;
assign f[58][182] = 9'b111111111;
assign f[58][183] = 9'b111111111;
assign f[58][184] = 9'b111111111;
assign f[58][185] = 9'b111111111;
assign f[59][26] = 9'b111111111;
assign f[59][27] = 9'b111111111;
assign f[59][28] = 9'b111111111;
assign f[59][29] = 9'b111111111;
assign f[59][30] = 9'b111111111;
assign f[59][31] = 9'b111111111;
assign f[59][32] = 9'b111111111;
assign f[59][42] = 9'b111111111;
assign f[59][43] = 9'b111111111;
assign f[59][44] = 9'b111111111;
assign f[59][45] = 9'b111111111;
assign f[59][46] = 9'b111111111;
assign f[59][47] = 9'b111111111;
assign f[59][48] = 9'b111111111;
assign f[59][56] = 9'b111111111;
assign f[59][57] = 9'b111111111;
assign f[59][58] = 9'b111111111;
assign f[59][59] = 9'b111111111;
assign f[59][60] = 9'b111111111;
assign f[59][61] = 9'b111111111;
assign f[59][62] = 9'b111111111;
assign f[59][65] = 9'b111111111;
assign f[59][66] = 9'b111111111;
assign f[59][67] = 9'b111111111;
assign f[59][68] = 9'b111111111;
assign f[59][69] = 9'b111111111;
assign f[59][70] = 9'b111111111;
assign f[59][71] = 9'b111111111;
assign f[59][72] = 9'b111111111;
assign f[59][94] = 9'b111111111;
assign f[59][95] = 9'b111111111;
assign f[59][96] = 9'b111111111;
assign f[59][97] = 9'b111111111;
assign f[59][98] = 9'b111111111;
assign f[59][99] = 9'b111111111;
assign f[59][100] = 9'b111111111;
assign f[59][117] = 9'b111111111;
assign f[59][118] = 9'b111111111;
assign f[59][119] = 9'b111111111;
assign f[59][120] = 9'b111111111;
assign f[59][121] = 9'b111111111;
assign f[59][122] = 9'b111111111;
assign f[59][123] = 9'b111111111;
assign f[59][124] = 9'b111111111;
assign f[59][138] = 9'b111111111;
assign f[59][139] = 9'b111111111;
assign f[59][140] = 9'b111111111;
assign f[59][141] = 9'b111111111;
assign f[59][142] = 9'b111111111;
assign f[59][143] = 9'b111111111;
assign f[59][153] = 9'b111111111;
assign f[59][154] = 9'b111111111;
assign f[59][155] = 9'b111111111;
assign f[59][156] = 9'b111111111;
assign f[59][157] = 9'b111111111;
assign f[59][158] = 9'b111111111;
assign f[59][159] = 9'b111111111;
assign f[59][160] = 9'b111111111;
assign f[59][163] = 9'b111111111;
assign f[59][164] = 9'b111111111;
assign f[59][165] = 9'b111111111;
assign f[59][166] = 9'b111111111;
assign f[59][167] = 9'b111111111;
assign f[59][168] = 9'b111111111;
assign f[59][169] = 9'b111111111;
assign f[59][174] = 9'b111111111;
assign f[59][175] = 9'b111111111;
assign f[59][176] = 9'b111111111;
assign f[59][177] = 9'b111111111;
assign f[59][178] = 9'b111111111;
assign f[59][179] = 9'b111111111;
assign f[59][180] = 9'b111111111;
assign f[59][181] = 9'b111111111;
assign f[59][182] = 9'b111111111;
assign f[59][183] = 9'b111111111;
assign f[59][184] = 9'b111111111;
assign f[59][185] = 9'b111111111;
assign f[60][26] = 9'b111111111;
assign f[60][27] = 9'b111111111;
assign f[60][28] = 9'b111111111;
assign f[60][29] = 9'b111111111;
assign f[60][30] = 9'b111111111;
assign f[60][31] = 9'b111111111;
assign f[60][32] = 9'b111111111;
assign f[60][33] = 9'b111111111;
assign f[60][41] = 9'b111111111;
assign f[60][42] = 9'b111111111;
assign f[60][43] = 9'b111111111;
assign f[60][44] = 9'b111111111;
assign f[60][45] = 9'b111111111;
assign f[60][46] = 9'b111111111;
assign f[60][47] = 9'b111111111;
assign f[60][48] = 9'b111111111;
assign f[60][56] = 9'b111111111;
assign f[60][57] = 9'b111111111;
assign f[60][58] = 9'b111111111;
assign f[60][59] = 9'b111111111;
assign f[60][60] = 9'b111111111;
assign f[60][61] = 9'b111111111;
assign f[60][62] = 9'b111111111;
assign f[60][65] = 9'b111111111;
assign f[60][66] = 9'b111111111;
assign f[60][67] = 9'b111111111;
assign f[60][68] = 9'b111111111;
assign f[60][69] = 9'b111111111;
assign f[60][70] = 9'b111111111;
assign f[60][71] = 9'b111111111;
assign f[60][72] = 9'b111111111;
assign f[60][73] = 9'b111111111;
assign f[60][74] = 9'b111111111;
assign f[60][75] = 9'b111111111;
assign f[60][76] = 9'b111111111;
assign f[60][77] = 9'b111111111;
assign f[60][78] = 9'b111111111;
assign f[60][79] = 9'b111111111;
assign f[60][80] = 9'b111111111;
assign f[60][81] = 9'b111111111;
assign f[60][94] = 9'b111111111;
assign f[60][95] = 9'b111111111;
assign f[60][96] = 9'b111111111;
assign f[60][97] = 9'b111111111;
assign f[60][98] = 9'b111111111;
assign f[60][99] = 9'b111111111;
assign f[60][100] = 9'b111111111;
assign f[60][117] = 9'b111111111;
assign f[60][118] = 9'b111111111;
assign f[60][119] = 9'b111111111;
assign f[60][120] = 9'b111111111;
assign f[60][121] = 9'b111111111;
assign f[60][122] = 9'b111111111;
assign f[60][123] = 9'b111111111;
assign f[60][124] = 9'b111111111;
assign f[60][125] = 9'b111111111;
assign f[60][126] = 9'b111111111;
assign f[60][127] = 9'b111111111;
assign f[60][129] = 9'b111111111;
assign f[60][130] = 9'b111111111;
assign f[60][131] = 9'b111111111;
assign f[60][138] = 9'b111111111;
assign f[60][139] = 9'b111111111;
assign f[60][140] = 9'b111111111;
assign f[60][141] = 9'b111111111;
assign f[60][142] = 9'b111111111;
assign f[60][143] = 9'b111111111;
assign f[60][154] = 9'b111111111;
assign f[60][155] = 9'b111111111;
assign f[60][156] = 9'b111111111;
assign f[60][157] = 9'b111111111;
assign f[60][158] = 9'b111111111;
assign f[60][159] = 9'b111111111;
assign f[60][160] = 9'b111111111;
assign f[60][163] = 9'b111111111;
assign f[60][164] = 9'b111111111;
assign f[60][165] = 9'b111111111;
assign f[60][166] = 9'b111111111;
assign f[60][167] = 9'b111111111;
assign f[60][168] = 9'b111111111;
assign f[60][169] = 9'b111111111;
assign f[60][175] = 9'b111111111;
assign f[60][176] = 9'b111111111;
assign f[60][177] = 9'b111111111;
assign f[60][178] = 9'b111111111;
assign f[60][179] = 9'b111111111;
assign f[60][180] = 9'b111111111;
assign f[60][181] = 9'b111111111;
assign f[60][182] = 9'b111111111;
assign f[60][183] = 9'b111111111;
assign f[60][184] = 9'b111111111;
assign f[60][185] = 9'b111111111;
assign f[61][26] = 9'b111111111;
assign f[61][27] = 9'b111111111;
assign f[61][28] = 9'b111111111;
assign f[61][29] = 9'b111111111;
assign f[61][30] = 9'b111111111;
assign f[61][31] = 9'b111111111;
assign f[61][32] = 9'b111111111;
assign f[61][33] = 9'b111111111;
assign f[61][41] = 9'b111111111;
assign f[61][42] = 9'b111111111;
assign f[61][43] = 9'b111111111;
assign f[61][44] = 9'b111111111;
assign f[61][45] = 9'b111111111;
assign f[61][46] = 9'b111111111;
assign f[61][47] = 9'b111111111;
assign f[61][48] = 9'b111111111;
assign f[61][56] = 9'b111111111;
assign f[61][57] = 9'b111111111;
assign f[61][58] = 9'b111111111;
assign f[61][59] = 9'b111111111;
assign f[61][60] = 9'b111111111;
assign f[61][61] = 9'b111111111;
assign f[61][62] = 9'b111111111;
assign f[61][65] = 9'b111111111;
assign f[61][66] = 9'b111111111;
assign f[61][67] = 9'b111111111;
assign f[61][68] = 9'b111111111;
assign f[61][69] = 9'b111111111;
assign f[61][70] = 9'b111111111;
assign f[61][71] = 9'b111111111;
assign f[61][72] = 9'b111111111;
assign f[61][73] = 9'b111111111;
assign f[61][74] = 9'b111111111;
assign f[61][75] = 9'b111111111;
assign f[61][76] = 9'b111111111;
assign f[61][77] = 9'b111111111;
assign f[61][78] = 9'b111111111;
assign f[61][79] = 9'b111111111;
assign f[61][80] = 9'b111111111;
assign f[61][81] = 9'b111111111;
assign f[61][94] = 9'b111111111;
assign f[61][95] = 9'b111111111;
assign f[61][96] = 9'b111111111;
assign f[61][97] = 9'b111111111;
assign f[61][98] = 9'b111111111;
assign f[61][99] = 9'b111111111;
assign f[61][100] = 9'b111111111;
assign f[61][117] = 9'b111111111;
assign f[61][118] = 9'b111111111;
assign f[61][119] = 9'b111111111;
assign f[61][120] = 9'b111111111;
assign f[61][121] = 9'b111111111;
assign f[61][122] = 9'b111111111;
assign f[61][123] = 9'b111111111;
assign f[61][124] = 9'b111111111;
assign f[61][125] = 9'b111111111;
assign f[61][126] = 9'b111111111;
assign f[61][127] = 9'b111111111;
assign f[61][128] = 9'b111111111;
assign f[61][129] = 9'b111111111;
assign f[61][130] = 9'b111111111;
assign f[61][131] = 9'b111111111;
assign f[61][132] = 9'b111111111;
assign f[61][137] = 9'b111111111;
assign f[61][138] = 9'b111111111;
assign f[61][139] = 9'b111111111;
assign f[61][140] = 9'b111111111;
assign f[61][141] = 9'b111111111;
assign f[61][142] = 9'b111111111;
assign f[61][143] = 9'b111111111;
assign f[61][154] = 9'b111111111;
assign f[61][155] = 9'b111111111;
assign f[61][156] = 9'b111111111;
assign f[61][157] = 9'b111111111;
assign f[61][158] = 9'b111111111;
assign f[61][159] = 9'b111111111;
assign f[61][160] = 9'b111111111;
assign f[61][163] = 9'b111111111;
assign f[61][164] = 9'b111111111;
assign f[61][165] = 9'b111111111;
assign f[61][166] = 9'b111111111;
assign f[61][167] = 9'b111111111;
assign f[61][168] = 9'b111111111;
assign f[61][169] = 9'b111111111;
assign f[61][175] = 9'b111111111;
assign f[61][176] = 9'b111111111;
assign f[61][177] = 9'b111111111;
assign f[61][178] = 9'b111111111;
assign f[61][179] = 9'b111111111;
assign f[61][180] = 9'b111111111;
assign f[61][181] = 9'b111111111;
assign f[61][182] = 9'b111111111;
assign f[61][183] = 9'b111111111;
assign f[61][184] = 9'b111111111;
assign f[61][185] = 9'b111111111;
assign f[62][26] = 9'b111111111;
assign f[62][27] = 9'b111111111;
assign f[62][28] = 9'b111111111;
assign f[62][29] = 9'b111111111;
assign f[62][30] = 9'b111111111;
assign f[62][31] = 9'b111111111;
assign f[62][32] = 9'b111111111;
assign f[62][33] = 9'b111111111;
assign f[62][41] = 9'b111111111;
assign f[62][42] = 9'b111111111;
assign f[62][43] = 9'b111111111;
assign f[62][44] = 9'b111111111;
assign f[62][45] = 9'b111111111;
assign f[62][46] = 9'b111111111;
assign f[62][47] = 9'b111111111;
assign f[62][48] = 9'b111111111;
assign f[62][56] = 9'b111111111;
assign f[62][57] = 9'b111111111;
assign f[62][58] = 9'b111111111;
assign f[62][59] = 9'b111111111;
assign f[62][60] = 9'b111111111;
assign f[62][61] = 9'b111111111;
assign f[62][62] = 9'b111111111;
assign f[62][65] = 9'b111111111;
assign f[62][66] = 9'b111111111;
assign f[62][67] = 9'b111111111;
assign f[62][68] = 9'b111111111;
assign f[62][69] = 9'b111111111;
assign f[62][70] = 9'b111111111;
assign f[62][71] = 9'b111111111;
assign f[62][72] = 9'b111111111;
assign f[62][73] = 9'b111111111;
assign f[62][74] = 9'b111111111;
assign f[62][75] = 9'b111111111;
assign f[62][76] = 9'b111111111;
assign f[62][77] = 9'b111111111;
assign f[62][78] = 9'b111111111;
assign f[62][79] = 9'b111111111;
assign f[62][80] = 9'b111111111;
assign f[62][81] = 9'b111111111;
assign f[62][94] = 9'b111111111;
assign f[62][95] = 9'b111111111;
assign f[62][96] = 9'b111111111;
assign f[62][97] = 9'b111111111;
assign f[62][98] = 9'b111111111;
assign f[62][99] = 9'b111111111;
assign f[62][100] = 9'b111111111;
assign f[62][117] = 9'b111111111;
assign f[62][118] = 9'b111111111;
assign f[62][119] = 9'b111111111;
assign f[62][120] = 9'b111111111;
assign f[62][121] = 9'b111111111;
assign f[62][122] = 9'b111111111;
assign f[62][123] = 9'b111111111;
assign f[62][124] = 9'b111111111;
assign f[62][125] = 9'b111111111;
assign f[62][126] = 9'b111111111;
assign f[62][127] = 9'b111111111;
assign f[62][128] = 9'b111111111;
assign f[62][129] = 9'b111111111;
assign f[62][130] = 9'b111111111;
assign f[62][131] = 9'b111111111;
assign f[62][132] = 9'b111111111;
assign f[62][137] = 9'b111111111;
assign f[62][138] = 9'b111111111;
assign f[62][139] = 9'b111111111;
assign f[62][140] = 9'b111111111;
assign f[62][141] = 9'b111111111;
assign f[62][142] = 9'b111111111;
assign f[62][143] = 9'b111111111;
assign f[62][154] = 9'b111111111;
assign f[62][155] = 9'b111111111;
assign f[62][156] = 9'b111111111;
assign f[62][157] = 9'b111111111;
assign f[62][158] = 9'b111111111;
assign f[62][159] = 9'b111111111;
assign f[62][160] = 9'b111111111;
assign f[62][163] = 9'b111111111;
assign f[62][164] = 9'b111111111;
assign f[62][165] = 9'b111111111;
assign f[62][166] = 9'b111111111;
assign f[62][167] = 9'b111111111;
assign f[62][168] = 9'b111111111;
assign f[62][169] = 9'b111111111;
assign f[62][175] = 9'b111111111;
assign f[62][176] = 9'b111111111;
assign f[62][177] = 9'b111111111;
assign f[62][178] = 9'b111111111;
assign f[62][179] = 9'b111111111;
assign f[62][180] = 9'b111111111;
assign f[62][181] = 9'b111111111;
assign f[62][182] = 9'b111111111;
assign f[62][183] = 9'b111111111;
assign f[62][184] = 9'b111111111;
assign f[62][185] = 9'b111111111;
assign f[63][26] = 9'b111111111;
assign f[63][27] = 9'b111111111;
assign f[63][28] = 9'b111111111;
assign f[63][29] = 9'b111111111;
assign f[63][30] = 9'b111111111;
assign f[63][31] = 9'b111111111;
assign f[63][32] = 9'b111111111;
assign f[63][33] = 9'b111111111;
assign f[63][42] = 9'b111111111;
assign f[63][43] = 9'b111111111;
assign f[63][44] = 9'b111111111;
assign f[63][45] = 9'b111111111;
assign f[63][46] = 9'b111111111;
assign f[63][47] = 9'b111111111;
assign f[63][48] = 9'b111111111;
assign f[63][56] = 9'b111111111;
assign f[63][57] = 9'b111111111;
assign f[63][58] = 9'b111111111;
assign f[63][59] = 9'b111111111;
assign f[63][60] = 9'b111111111;
assign f[63][61] = 9'b111111111;
assign f[63][62] = 9'b111111111;
assign f[63][65] = 9'b111111111;
assign f[63][66] = 9'b111111111;
assign f[63][67] = 9'b111111111;
assign f[63][68] = 9'b111111111;
assign f[63][69] = 9'b111111111;
assign f[63][70] = 9'b111111111;
assign f[63][71] = 9'b111111111;
assign f[63][72] = 9'b111111111;
assign f[63][73] = 9'b111111111;
assign f[63][74] = 9'b111111111;
assign f[63][75] = 9'b111111111;
assign f[63][76] = 9'b111111111;
assign f[63][77] = 9'b111111111;
assign f[63][78] = 9'b111111111;
assign f[63][79] = 9'b111111111;
assign f[63][80] = 9'b111111111;
assign f[63][81] = 9'b111111111;
assign f[63][94] = 9'b111111111;
assign f[63][95] = 9'b111111111;
assign f[63][96] = 9'b111111111;
assign f[63][97] = 9'b111111111;
assign f[63][98] = 9'b111111111;
assign f[63][99] = 9'b111111111;
assign f[63][100] = 9'b111111111;
assign f[63][117] = 9'b111111111;
assign f[63][118] = 9'b111111111;
assign f[63][119] = 9'b111111111;
assign f[63][120] = 9'b111111111;
assign f[63][121] = 9'b111111111;
assign f[63][122] = 9'b111111111;
assign f[63][123] = 9'b111111111;
assign f[63][124] = 9'b111111111;
assign f[63][125] = 9'b111111111;
assign f[63][126] = 9'b111111111;
assign f[63][127] = 9'b111111111;
assign f[63][128] = 9'b111111111;
assign f[63][129] = 9'b111111111;
assign f[63][130] = 9'b111111111;
assign f[63][131] = 9'b111111111;
assign f[63][137] = 9'b111111111;
assign f[63][138] = 9'b111111111;
assign f[63][139] = 9'b111111111;
assign f[63][140] = 9'b111111111;
assign f[63][141] = 9'b111111111;
assign f[63][142] = 9'b111111111;
assign f[63][154] = 9'b111111111;
assign f[63][155] = 9'b111111111;
assign f[63][156] = 9'b111111111;
assign f[63][157] = 9'b111111111;
assign f[63][158] = 9'b111111111;
assign f[63][159] = 9'b111111111;
assign f[63][160] = 9'b111111111;
assign f[63][161] = 9'b111111111;
assign f[63][163] = 9'b111111111;
assign f[63][164] = 9'b111111111;
assign f[63][165] = 9'b111111111;
assign f[63][166] = 9'b111111111;
assign f[63][167] = 9'b111111111;
assign f[63][168] = 9'b111111111;
assign f[63][169] = 9'b111111111;
assign f[63][175] = 9'b111111111;
assign f[63][176] = 9'b111111111;
assign f[63][177] = 9'b111111111;
assign f[63][178] = 9'b111111111;
assign f[63][179] = 9'b111111111;
assign f[63][180] = 9'b111111111;
assign f[63][181] = 9'b111111111;
assign f[63][182] = 9'b111111111;
assign f[63][183] = 9'b111111111;
assign f[63][184] = 9'b111111111;
assign f[63][185] = 9'b111111111;
assign f[64][26] = 9'b111111111;
assign f[64][27] = 9'b111111111;
assign f[64][28] = 9'b111111111;
assign f[64][29] = 9'b111111111;
assign f[64][30] = 9'b111111111;
assign f[64][31] = 9'b111111111;
assign f[64][32] = 9'b111111111;
assign f[64][33] = 9'b111111111;
assign f[64][42] = 9'b111111111;
assign f[64][43] = 9'b111111111;
assign f[64][44] = 9'b111111111;
assign f[64][45] = 9'b111111111;
assign f[64][46] = 9'b111111111;
assign f[64][47] = 9'b111111111;
assign f[64][48] = 9'b111111111;
assign f[64][55] = 9'b111111111;
assign f[64][56] = 9'b111111111;
assign f[64][57] = 9'b111111111;
assign f[64][58] = 9'b111111111;
assign f[64][59] = 9'b111111111;
assign f[64][60] = 9'b111111111;
assign f[64][61] = 9'b111111111;
assign f[64][62] = 9'b111111111;
assign f[64][65] = 9'b111111111;
assign f[64][66] = 9'b111111111;
assign f[64][67] = 9'b111111111;
assign f[64][68] = 9'b111111111;
assign f[64][69] = 9'b111111111;
assign f[64][70] = 9'b111111111;
assign f[64][71] = 9'b111111111;
assign f[64][72] = 9'b111111111;
assign f[64][73] = 9'b111111111;
assign f[64][74] = 9'b111111111;
assign f[64][75] = 9'b111111111;
assign f[64][76] = 9'b111111111;
assign f[64][77] = 9'b111111111;
assign f[64][78] = 9'b111111111;
assign f[64][79] = 9'b111111111;
assign f[64][80] = 9'b111111111;
assign f[64][81] = 9'b111111111;
assign f[64][82] = 9'b111111111;
assign f[64][94] = 9'b111111111;
assign f[64][95] = 9'b111111111;
assign f[64][96] = 9'b111111111;
assign f[64][97] = 9'b111111111;
assign f[64][98] = 9'b111111111;
assign f[64][99] = 9'b111111111;
assign f[64][100] = 9'b111111111;
assign f[64][117] = 9'b111111111;
assign f[64][118] = 9'b111111111;
assign f[64][119] = 9'b111111111;
assign f[64][120] = 9'b111111111;
assign f[64][121] = 9'b111111111;
assign f[64][122] = 9'b111111111;
assign f[64][123] = 9'b111111111;
assign f[64][124] = 9'b111111111;
assign f[64][125] = 9'b111111111;
assign f[64][126] = 9'b111111111;
assign f[64][127] = 9'b111111111;
assign f[64][128] = 9'b111111111;
assign f[64][129] = 9'b111111111;
assign f[64][130] = 9'b111111111;
assign f[64][131] = 9'b111111111;
assign f[64][132] = 9'b111111111;
assign f[64][137] = 9'b111111111;
assign f[64][138] = 9'b111111111;
assign f[64][139] = 9'b111111111;
assign f[64][140] = 9'b111111111;
assign f[64][141] = 9'b111111111;
assign f[64][142] = 9'b111111111;
assign f[64][155] = 9'b111111111;
assign f[64][156] = 9'b111111111;
assign f[64][157] = 9'b111111111;
assign f[64][158] = 9'b111111111;
assign f[64][159] = 9'b111111111;
assign f[64][160] = 9'b111111111;
assign f[64][161] = 9'b111111111;
assign f[64][163] = 9'b111111111;
assign f[64][164] = 9'b111111111;
assign f[64][165] = 9'b111111111;
assign f[64][166] = 9'b111111111;
assign f[64][167] = 9'b111111111;
assign f[64][168] = 9'b111111111;
assign f[64][169] = 9'b111111111;
assign f[64][176] = 9'b111111111;
assign f[64][177] = 9'b111111111;
assign f[64][178] = 9'b111111111;
assign f[64][179] = 9'b111111111;
assign f[64][180] = 9'b111111111;
assign f[64][181] = 9'b111111111;
assign f[64][182] = 9'b111111111;
assign f[64][183] = 9'b111111111;
assign f[64][184] = 9'b111111111;
assign f[64][185] = 9'b111111111;
assign f[65][27] = 9'b111111111;
assign f[65][28] = 9'b111111111;
assign f[65][29] = 9'b111111111;
assign f[65][30] = 9'b111111111;
assign f[65][31] = 9'b111111111;
assign f[65][32] = 9'b111111111;
assign f[65][42] = 9'b111111111;
assign f[65][43] = 9'b111111111;
assign f[65][44] = 9'b111111111;
assign f[65][45] = 9'b111111111;
assign f[65][46] = 9'b111111111;
assign f[65][47] = 9'b111111111;
assign f[65][56] = 9'b111111111;
assign f[65][57] = 9'b111111111;
assign f[65][58] = 9'b111111111;
assign f[65][59] = 9'b111111111;
assign f[65][60] = 9'b111111111;
assign f[65][61] = 9'b111111111;
assign f[65][65] = 9'b111111111;
assign f[65][66] = 9'b111111111;
assign f[65][67] = 9'b111111111;
assign f[65][68] = 9'b111111111;
assign f[65][69] = 9'b111111111;
assign f[65][70] = 9'b111111111;
assign f[65][71] = 9'b111111111;
assign f[65][72] = 9'b111111111;
assign f[65][74] = 9'b111111111;
assign f[65][75] = 9'b111111111;
assign f[65][76] = 9'b111111111;
assign f[65][77] = 9'b111111111;
assign f[65][78] = 9'b111111111;
assign f[65][79] = 9'b111111111;
assign f[65][80] = 9'b111111111;
assign f[65][81] = 9'b111111111;
assign f[65][95] = 9'b111111111;
assign f[65][96] = 9'b111111111;
assign f[65][97] = 9'b111111111;
assign f[65][98] = 9'b111111111;
assign f[65][99] = 9'b111111111;
assign f[65][100] = 9'b111111111;
assign f[65][117] = 9'b111111111;
assign f[65][118] = 9'b111111111;
assign f[65][119] = 9'b111111111;
assign f[65][120] = 9'b111111111;
assign f[65][121] = 9'b111111111;
assign f[65][122] = 9'b111111111;
assign f[65][123] = 9'b111111111;
assign f[65][124] = 9'b111111111;
assign f[65][125] = 9'b111111111;
assign f[65][126] = 9'b111111111;
assign f[65][127] = 9'b111111111;
assign f[65][129] = 9'b111111111;
assign f[65][130] = 9'b111111111;
assign f[65][137] = 9'b111111111;
assign f[65][138] = 9'b111111111;
assign f[65][139] = 9'b111111111;
assign f[65][140] = 9'b111111111;
assign f[65][141] = 9'b111111111;
assign f[65][155] = 9'b111111111;
assign f[65][156] = 9'b111111111;
assign f[65][157] = 9'b111111111;
assign f[65][158] = 9'b111111111;
assign f[65][159] = 9'b111111111;
assign f[65][160] = 9'b111111111;
assign f[65][161] = 9'b111111111;
assign f[65][164] = 9'b111111111;
assign f[65][165] = 9'b111111111;
assign f[65][166] = 9'b111111111;
assign f[65][167] = 9'b111111111;
assign f[65][168] = 9'b111111111;
assign f[65][176] = 9'b111111111;
assign f[65][177] = 9'b111111111;
assign f[65][178] = 9'b111111111;
assign f[65][179] = 9'b111111111;
assign f[65][180] = 9'b111111111;
assign f[65][181] = 9'b111111111;
assign f[65][182] = 9'b111111111;
assign f[65][183] = 9'b111111111;
assign f[65][184] = 9'b111111111;
//Total de Lineas = 3080
endmodule


